-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 23 2022 02:01:15

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    led : out std_logic_vector(7 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__34843\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \M_this_map_ram_read_data_4\ : std_logic;
signal \M_this_ppu_sprites_addr_9\ : std_logic;
signal \M_this_ppu_sprites_addr_8\ : std_logic;
signal \M_this_ppu_sprites_addr_7\ : std_logic;
signal \M_this_ppu_sprites_addr_6\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal port_nmib_0_i : std_logic;
signal port_clk_c : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal rgb_c_5 : std_logic;
signal port_data_rw_0_i : std_logic;
signal rgb_c_0 : std_logic;
signal rgb_c_1 : std_logic;
signal rgb_c_3 : std_logic;
signal rgb_c_4 : std_logic;
signal \this_vga_ramdac.N_2870_reto\ : std_logic;
signal rgb_c_2 : std_logic;
signal \this_vga_ramdac.i2_mux_0\ : std_logic;
signal \this_vga_ramdac.N_2875_reto\ : std_logic;
signal \this_vga_signals.un4_hsynclto7_0_cascade_\ : std_logic;
signal this_vga_signals_hsync_1_i : std_logic;
signal \this_vga_signals.un2_hsynclt7_cascade_\ : std_logic;
signal \this_vga_signals.hsync_1_0\ : std_logic;
signal this_vga_signals_hvisibility_i : std_logic;
signal \this_vga_signals.if_N_8_i_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_9_0_0_cascade_\ : std_logic;
signal \this_pixel_clk.M_counter_q_i_1\ : std_logic;
signal \this_pixel_clk.M_counter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_0_3_cascade_\ : std_logic;
signal \this_vga_signals.N_614_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_0\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_2\ : std_logic;
signal \this_vga_signals.N_931_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNI0JBR6Z0Z_9\ : std_logic;
signal \this_vga_signals.un4_hsynclto3_0\ : std_logic;
signal \this_vga_signals.un2_hsynclt6_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lt7_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lto7_1\ : std_logic;
signal this_vga_signals_vvisibility_i : std_logic;
signal \this_vga_signals.N_5_i_5\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0\ : std_logic;
signal \this_vga_signals.g0_4_cascade_\ : std_logic;
signal \this_vga_signals.g0_7_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \this_vga_ramdac.N_24_mux\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1\ : std_logic;
signal \this_vga_signals.g1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g2_0_0\ : std_logic;
signal \this_vga_signals.if_N_9_0_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_1\ : std_logic;
signal \this_vga_signals.N_236_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_3_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_\ : std_logic;
signal \this_vga_signals.N_3_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.SUM_3_i_0_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\ : std_logic;
signal \this_vga_signals.N_236\ : std_logic;
signal \this_vga_signals.SUM_3_i_0_0_3\ : std_logic;
signal \this_vga_signals.g0_1\ : std_logic;
signal \this_vga_signals.un6_vvisibilitylt8_cascade_\ : std_logic;
signal \this_vga_signals.vvisibility_1_cascade_\ : std_logic;
signal \this_vga_signals.vsync_1_3\ : std_logic;
signal \this_vga_signals.vsync_1_2_cascade_\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \this_vga_signals.if_m7_0_x4_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_9_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.d_N_12\ : std_logic;
signal \this_vga_signals.d_N_11\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNIUAKU9Z0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3\ : std_logic;
signal \this_vga_signals.N_2_7_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_3_d\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lt4\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.N_614_0\ : std_logic;
signal \this_vga_signals.N_931_1\ : std_logic;
signal \this_vga_signals.vaddress_0_5_cascade_\ : std_logic;
signal \this_vga_signals.g0_31_N_4L6\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_4_cascade_\ : std_logic;
signal \this_vga_signals.g0_31_N_3L3\ : std_logic;
signal \this_vga_signals.g3_3_0\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_2_cascade_\ : std_logic;
signal \this_vga_signals.g0_8_0_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_2_5_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_3_0_6_cascade_\ : std_logic;
signal \this_vga_signals.g2_3_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_2_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_6_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_1_0_0\ : std_logic;
signal \this_vga_signals.vaddress_3_0_6\ : std_logic;
signal \this_vga_signals.vaddress_3_5_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_3_6_cascade_\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_3\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_3\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_3\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \this_vga_ramdac.m19\ : std_logic;
signal \this_vga_ramdac.N_2874_reto\ : std_logic;
signal \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_3\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\ : std_logic;
signal \bfn_10_11_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.vaddress_c2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_1\ : std_logic;
signal \this_vga_signals.g0_31_N_5L8\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_0\ : std_logic;
signal \this_vga_signals.m9_1_cascade_\ : std_logic;
signal \this_vga_signals.g2_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_1_0\ : std_logic;
signal \this_vga_signals.g1_0_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g2_0_1_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_6_6\ : std_logic;
signal \this_vga_signals.N_4_1_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_0\ : std_logic;
signal \this_vga_signals.g1_4_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_1_0_0_1\ : std_logic;
signal \this_vga_signals.g0_2_0_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_3_2\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \this_sprites_ram.mem_WE_6\ : std_logic;
signal \this_vga_signals.N_3_2_1\ : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lto8_1\ : std_logic;
signal \this_vga_signals.M_lcounter_d_0_sqmuxa\ : std_logic;
signal \this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_\ : std_logic;
signal \N_2_0_cascade_\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_0\ : std_logic;
signal \M_counter_q_RNILQS8_1\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_1_cascade_\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_1\ : std_logic;
signal \N_3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_5_1\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_5_0\ : std_logic;
signal \this_vga_signals.M_hcounter_d7_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_0\ : std_logic;
signal \this_sprites_ram.mem_WE_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.N_1_4_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_0\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_2_3_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_8_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_0_3\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5Z0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJHZ0Z5\ : std_logic;
signal \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i_cascade_\ : std_logic;
signal \this_vga_signals.N_50\ : std_logic;
signal \this_vga_signals.vaddress_1_6_cascade_\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals.N_614_1_g\ : std_logic;
signal \this_vga_signals.N_931_g\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_1_cascade_\ : std_logic;
signal \this_vga_signals.if_N_5_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_5_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_0\ : std_logic;
signal \this_vga_signals.g0_1_2_0_1\ : std_logic;
signal \this_vga_signals.g0_1_2_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_1_0_0\ : std_logic;
signal \this_vga_signals.g2_0\ : std_logic;
signal \this_vga_signals.g1_1_1\ : std_logic;
signal \this_vga_signals.N_5_i_0\ : std_logic;
signal \this_vga_signals.g0_2_0_2_x1\ : std_logic;
signal \this_vga_signals.g0_2_0_2_x0_cascade_\ : std_logic;
signal \this_vga_signals.g0_2_0_2_cascade_\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_0\ : std_logic;
signal \this_sprites_ram.mem_WE_8\ : std_logic;
signal \this_vga_ramdac.m6\ : std_logic;
signal \this_vga_ramdac.N_2871_reto\ : std_logic;
signal \G_384_cascade_\ : std_logic;
signal \this_vga_ramdac.N_2872_reto\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \G_384\ : std_logic;
signal \this_vga_ramdac.N_2873_reto\ : std_logic;
signal \N_3_0\ : std_logic;
signal \N_2_0\ : std_logic;
signal \M_this_vga_signals_pixel_clk_0_0\ : std_logic;
signal \this_sprites_ram.mem_WE_2\ : std_logic;
signal \M_this_ppu_vram_addr_7\ : std_logic;
signal \M_this_ppu_sprites_addr_4\ : std_logic;
signal \this_vga_signals.vaddress_4_5\ : std_logic;
signal \this_vga_signals.vaddress_5\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.N_5_i_0_0\ : std_logic;
signal \this_vga_signals.i2_mux\ : std_logic;
signal \this_vga_signals.i2_mux_cascade_\ : std_logic;
signal \this_vga_signals.if_i2_mux_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_0_6\ : std_logic;
signal \this_vga_signals.g2_2\ : std_logic;
signal \m18x_N_3LZ0Z3\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNI5BS7NZ0Z_5\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_0_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_0_x1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0\ : std_logic;
signal \this_vga_signals.g0_2_0_2\ : std_logic;
signal \this_vga_signals.g1_0_0_0_1\ : std_logic;
signal \this_vga_signals.N_51\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0\ : std_logic;
signal \this_vga_signals.g2_1\ : std_logic;
signal \this_vga_signals.g1_0\ : std_logic;
signal \this_vga_signals.g1_N_4L5_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5EZ0Z1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2\ : std_logic;
signal \this_vga_signals.g0_1_1\ : std_logic;
signal \this_vga_signals.d_N_3_0_i\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_x0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.g0_7\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_0\ : std_logic;
signal this_vga_signals_un5_vaddress_g1_1_0 : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_0\ : std_logic;
signal \this_vga_signals.g1_2\ : std_logic;
signal \this_vga_signals.m21_0_1_1\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\ : std_logic;
signal \M_this_ppu_vram_data_0\ : std_logic;
signal \this_vga_ramdac.m16\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \this_vga_ramdac.i2_mux\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.line_clk_1\ : std_logic;
signal \M_this_vga_signals_line_clk_0_cascade_\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_cascade_\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_1\ : std_logic;
signal this_vga_signals_vvisibility : std_logic;
signal \this_vga_signals.vaddress_2_5\ : std_logic;
signal \this_vga_signals.g1_1_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_0_0\ : std_logic;
signal \this_vga_signals.g1_2_0_0\ : std_logic;
signal \this_vga_signals.if_i2_mux\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt3\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt9_1\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt9_1_cascade_\ : std_logic;
signal \this_vga_signals.un4_lvisibility_1\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_0\ : std_logic;
signal \this_vga_signals.g0_0\ : std_logic;
signal \this_vga_signals.vaddress_1_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_0_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_1_5\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \this_vga_signals.vaddress_2_6_cascade_\ : std_logic;
signal \this_vga_signals.g1_2_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNITP439_0Z0Z_2_cascade_\ : std_logic;
signal \this_vga_signals.m16_0_1\ : std_logic;
signal this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i : std_logic;
signal this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0 : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_12\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNITP439Z0Z_2\ : std_logic;
signal \this_vga_signals.g2_1_1\ : std_logic;
signal \this_vga_signals.g1_1_1_0\ : std_logic;
signal \this_vga_signals.if_N_5_1\ : std_logic;
signal \this_vga_signals.g0_5_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2_0\ : std_logic;
signal \this_vga_signals.g0_1_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3\ : std_logic;
signal \this_vga_signals.g0_1_2_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1\ : std_logic;
signal if_generate_plus_mult1_un68_sum_axb1_520 : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_i\ : std_logic;
signal \this_vga_signals.g2_0_0_0\ : std_logic;
signal \this_vga_signals.g1_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i\ : std_logic;
signal \this_vga_signals.g1_0_2\ : std_logic;
signal \this_vga_signals.g0_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_0_0_0\ : std_logic;
signal \this_vga_signals.m21_0_1\ : std_logic;
signal \this_vga_signals.i14_mux_i\ : std_logic;
signal \this_vga_signals.N_25_0_0_cascade_\ : std_logic;
signal \this_vga_signals.i13_mux_0_i\ : std_logic;
signal \this_vga_signals.if_i1_mux\ : std_logic;
signal \this_vga_signals.g1_0_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_N_4L5_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_N_4L5_cascade_\ : std_logic;
signal \this_vga_signals.N_5_i\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_2\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2\ : std_logic;
signal \this_ppu.M_last_q_RNIMRAD5_4\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4\ : std_logic;
signal \this_ppu.M_last_q_RNIMRAD5_5\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_6\ : std_logic;
signal \this_ppu.M_last_q_RNIMRAD5_1\ : std_logic;
signal \this_ppu.M_last_q_RNIMRAD5_0\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_4\ : std_logic;
signal \this_ppu.un1_M_count_q_1_axb_0_cascade_\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_6\ : std_logic;
signal \this_ppu.line_clk.M_last_qZ0\ : std_logic;
signal \M_this_vga_signals_line_clk_0\ : std_logic;
signal \this_ppu.N_82_i_cascade_\ : std_logic;
signal \this_ppu.M_last_q_RNIMRAD5_3\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_0\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z2\ : std_logic;
signal \this_vga_signals.if_N_5_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_4\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_5\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_2\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_1\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\ : std_logic;
signal \this_ppu.N_91_cascade_\ : std_logic;
signal \this_ppu.M_count_qZ1Z_1\ : std_logic;
signal \this_ppu.M_count_qZ1Z_2\ : std_logic;
signal \this_ppu.M_count_qZ1Z_0\ : std_logic;
signal \this_ppu.M_state_q_i_1_cascade_\ : std_logic;
signal \this_ppu.M_last_q_RNIMRAD5_2\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_3\ : std_logic;
signal \this_ppu.M_count_qZ1Z_3\ : std_logic;
signal \this_ppu.M_count_qZ1Z_4\ : std_logic;
signal \this_ppu.M_count_qZ0Z_6\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_5\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4_cascade_\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_1\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_1_cascade_\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_5\ : std_logic;
signal \this_ppu.M_count_qZ1Z_5\ : std_logic;
signal \this_ppu.M_state_q_i_1\ : std_logic;
signal \this_ppu.M_count_qZ0Z_7\ : std_logic;
signal \this_ppu.N_82_i\ : std_logic;
signal \this_ppu.un1_M_count_q_1_axb_7\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_1\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2\ : std_logic;
signal \M_this_ppu_vram_data_2\ : std_logic;
signal \this_ppu.M_state_qZ0Z_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_1\ : std_logic;
signal \this_sprites_ram.mem_WE_0\ : std_logic;
signal \M_this_ppu_map_addr_6\ : std_logic;
signal \M_this_ppu_map_addr_5\ : std_logic;
signal \M_this_ppu_sprites_addr_5\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c2\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \this_sprites_ram.mem_WE_14\ : std_logic;
signal \this_sprites_ram.mem_WE_12\ : std_logic;
signal \M_this_sprites_ram_write_en_0\ : std_logic;
signal \this_sprites_ram.mem_WE_10\ : std_logic;
signal \M_this_sprites_ram_write_data_0\ : std_logic;
signal \M_this_sprites_ram_write_data_1\ : std_logic;
signal \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux_cascade_\ : std_logic;
signal \M_this_sprites_ram_write_data_2\ : std_logic;
signal \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\ : std_logic;
signal \M_this_sprites_ram_write_data_3\ : std_logic;
signal \M_this_vga_ramdac_en_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \M_this_ppu_map_addr_7\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c5\ : std_logic;
signal \this_ppu.M_last_q_RNIQKTIG\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_7\ : std_logic;
signal \M_this_ppu_map_addr_9\ : std_logic;
signal \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_8\ : std_logic;
signal \this_vga_signals.un23_i_a2_x1Z0Z_0_cascade_\ : std_logic;
signal \dma_ac0Z0Z_5\ : std_logic;
signal this_vga_signals_un23_i_a2_1_3 : std_logic;
signal this_vga_signals_un23_i_a2_4_2 : std_logic;
signal \this_vga_signals_un23_i_a2_3_2_cascade_\ : std_logic;
signal dma_c3_0 : std_logic;
signal dma_axb0 : std_logic;
signal \M_this_state_q_RNI2S2SZ0Z_13\ : std_logic;
signal \M_this_state_q_RNITS9I4Z0Z_7_cascade_\ : std_logic;
signal dma_ac0_5_i : std_logic;
signal \dma_ac0_5_i_cascade_\ : std_logic;
signal dma_ac0_5_i_i : std_logic;
signal \this_vga_signals.un23_i_a2_4Z0Z_0\ : std_logic;
signal \M_this_state_q_RNI6Q0SZ0Z_7\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_3\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \M_this_ppu_vram_en_0\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_1\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_9\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2_cascade_\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_2\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_3\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_10\ : std_logic;
signal \M_this_state_q_RNIMJ231Z0Z_8\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_15\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7\ : std_logic;
signal \M_this_sprites_address_qZ0Z_8\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \M_this_sprites_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8\ : std_logic;
signal \M_this_sprites_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_13\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_13\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_o2_0_0_0\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_o2_0_1Z0Z_0_cascade_\ : std_logic;
signal \M_this_sprites_address_q_RNI1DGI7Z0Z_0\ : std_logic;
signal \M_this_map_ram_read_data_5\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_11\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_2_cascade_\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_8_mZ0Z_2\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_9\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_5_mZ0Z_9\ : std_logic;
signal \M_this_ppu_map_addr_1\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c2\ : std_logic;
signal \M_this_ppu_map_addr_0\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_6\ : std_logic;
signal \this_ppu_M_vaddress_q_i_6\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_6\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6_cascade_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_5\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_6\ : std_logic;
signal \this_vga_signals.N_294_cascade_\ : std_logic;
signal \this_vga_signals.un1_M_this_state_q_14Z0Z_1_cascade_\ : std_logic;
signal \un1_M_this_state_q_14_0\ : std_logic;
signal this_vga_signals_un23_i_a2_1_1 : std_logic;
signal un23_i_a2_1 : std_logic;
signal \this_vga_signals.N_486\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_5\ : std_logic;
signal \this_vga_signals.N_486_cascade_\ : std_logic;
signal \this_vga_signals.N_438_1\ : std_logic;
signal \this_vga_signals_M_this_state_q_ns_i_o2_0_12\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_11\ : std_logic;
signal \this_vga_signals.N_446_1\ : std_logic;
signal \M_this_sprites_address_qZ0Z_11\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_7\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_4\ : std_logic;
signal \this_vga_signals.un1_M_this_state_q_19_0\ : std_logic;
signal \this_vga_signals.M_this_state_d_1_sqmuxaZ0_cascade_\ : std_logic;
signal \this_vga_signals.N_399_0\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_5_mZ0Z_5\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_5_cascade_\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_0\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_6\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_5_mZ0Z_6_cascade_\ : std_logic;
signal \M_this_map_address_q_RNICF7V6Z0Z_0\ : std_logic;
signal \bfn_19_22_0_\ : std_logic;
signal \un1_M_this_map_address_q_cry_0\ : std_logic;
signal \M_this_map_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_map_address_q_cry_1_c_RNI8JSRZ0\ : std_logic;
signal \un1_M_this_map_address_q_cry_1\ : std_logic;
signal \un1_M_this_map_address_q_cry_2\ : std_logic;
signal \un1_M_this_map_address_q_cry_3\ : std_logic;
signal \M_this_map_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_map_address_q_cry_4_c_RNIESVRZ0\ : std_logic;
signal \un1_M_this_map_address_q_cry_4\ : std_logic;
signal \M_this_map_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_5_c_RNIGV0SZ0\ : std_logic;
signal \un1_M_this_map_address_q_cry_5\ : std_logic;
signal \un1_M_this_map_address_q_cry_6_c_RNII22SZ0\ : std_logic;
signal \un1_M_this_map_address_q_cry_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_7\ : std_logic;
signal \bfn_19_23_0_\ : std_logic;
signal \M_this_map_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_map_address_q_cry_8\ : std_logic;
signal \un1_M_this_map_address_q_cry_8_c_RNIM84SZ0\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_5_mZ0Z_7\ : std_logic;
signal \M_this_map_address_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_7\ : std_logic;
signal \M_this_ppu_map_addr_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c5\ : std_logic;
signal \this_ppu.M_last_q_RNI21NK5\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_6\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \M_this_sprites_address_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5\ : std_logic;
signal \M_this_sprites_address_qZ0Z_1\ : std_logic;
signal \N_389_0_cascade_\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1\ : std_logic;
signal \M_this_state_q_fastZ0Z_15\ : std_logic;
signal \N_297\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_9\ : std_logic;
signal \M_this_state_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_a3_sxZ0Z_9_cascade_\ : std_logic;
signal port_address_in_4 : std_logic;
signal port_rw_in : std_logic;
signal port_address_in_7 : std_logic;
signal \this_vga_signals.N_291\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1\ : std_logic;
signal port_address_in_5 : std_logic;
signal port_address_in_6 : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_4_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0\ : std_logic;
signal \this_vga_signals.N_444_1\ : std_logic;
signal \this_vga_signals_M_this_state_q_ns_i_o2_0_14\ : std_logic;
signal \M_this_state_q_fastZ0Z_14\ : std_logic;
signal \M_this_sprites_address_qZ0Z_12\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_12\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_5Z0Z_14\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_14\ : std_logic;
signal \M_this_sprites_address_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4\ : std_logic;
signal \M_this_map_address_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_8_mZ0Z_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_8_mZ0Z_1\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_1_cascade_\ : std_logic;
signal \un1_M_this_map_address_q_cry_0_c_RNI6GRRZ0\ : std_logic;
signal \M_this_map_address_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_8_mZ0Z_3_cascade_\ : std_logic;
signal \un1_M_this_map_address_q_cry_2_c_RNIAMTRZ0\ : std_logic;
signal \M_this_map_address_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_3\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_8_mZ0Z_4\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_4\ : std_logic;
signal \un1_M_this_map_address_q_cry_3_c_RNICPURZ0\ : std_logic;
signal \M_this_map_address_qZ0Z_4\ : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \un1_M_this_state_q_12_0\ : std_logic;
signal \this_vga_signals.M_this_map_address_d_5_mZ0Z_8\ : std_logic;
signal \this_vga_signals.un1_M_this_map_ram_write_en_0\ : std_logic;
signal \un1_M_this_map_address_q_cry_7_c_RNIK53SZ0\ : std_logic;
signal \N_989_g\ : std_logic;
signal \this_vga_signals.N_469\ : std_logic;
signal \M_this_state_qZ0Z_14\ : std_logic;
signal \this_start_data_delay_M_last_q\ : std_logic;
signal port_enb_c : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal port_address_in_2 : std_logic;
signal port_address_in_0 : std_logic;
signal port_address_in_3 : std_logic;
signal port_address_in_1 : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_10\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_5Z0Z_13_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_d_1_sqmuxaZ0\ : std_logic;
signal \this_vga_signals.M_this_state_d_0_sqmuxaZ0Z_1\ : std_logic;
signal \this_vga_signals.un1_M_this_state_q_21_0_cascade_\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_13\ : std_logic;
signal \M_this_state_qZ0Z_12\ : std_logic;
signal \this_vga_signals.N_293_1\ : std_logic;
signal \M_this_state_qZ0Z_15\ : std_logic;
signal \this_vga_signals.M_this_map_ram_write_data_1_sqmuxa\ : std_logic;
signal \this_vga_signals.N_293_cascade_\ : std_logic;
signal \M_this_map_ram_read_data_7\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_8_mZ0Z_5\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_5\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_6\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_8_mZ0Z_6_cascade_\ : std_logic;
signal \M_this_map_address_qZ0Z_8\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_this_map_address_q_mZ0Z_8\ : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_7\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_8\ : std_logic;
signal \M_this_sprites_address_qZ0Z_3\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3\ : std_logic;
signal \M_this_state_d88_1_cascade_\ : std_logic;
signal \this_vga_signals.N_390_0\ : std_logic;
signal \M_this_state_d88_12_cascade_\ : std_logic;
signal \N_507_cascade_\ : std_logic;
signal \N_508_cascade_\ : std_logic;
signal \M_this_state_d88_11\ : std_logic;
signal \M_this_state_d88_11_cascade_\ : std_logic;
signal \M_this_state_d88_12\ : std_logic;
signal \N_436\ : std_logic;
signal \N_465\ : std_logic;
signal \N_435\ : std_logic;
signal \M_this_state_qsr_0_cascade_\ : std_logic;
signal \N_466\ : std_logic;
signal led_c_1 : std_logic;
signal \M_this_state_d88\ : std_logic;
signal \un1_M_this_state_q_16_0\ : std_logic;
signal \bfn_22_20_0_\ : std_logic;
signal \un1_M_this_external_address_q_cry_0\ : std_logic;
signal \un1_M_this_external_address_q_cry_1\ : std_logic;
signal \un1_M_this_external_address_q_cry_2\ : std_logic;
signal \un1_M_this_external_address_q_cry_3\ : std_logic;
signal \M_this_external_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_external_address_q_cry_4_c_RNIOSKBZ0\ : std_logic;
signal \un1_M_this_external_address_q_cry_4\ : std_logic;
signal \M_this_external_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_5_c_RNIQVLBZ0\ : std_logic;
signal \un1_M_this_external_address_q_cry_5\ : std_logic;
signal \un1_M_this_external_address_q_cry_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_7\ : std_logic;
signal \bfn_22_21_0_\ : std_logic;
signal \un1_M_this_external_address_q_cry_8\ : std_logic;
signal \un1_M_this_external_address_q_cry_9\ : std_logic;
signal \un1_M_this_external_address_q_cry_10\ : std_logic;
signal \un1_M_this_external_address_q_cry_11\ : std_logic;
signal \M_this_external_address_qZ0Z_13\ : std_logic;
signal \un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0\ : std_logic;
signal \un1_M_this_external_address_q_cry_12\ : std_logic;
signal \M_this_external_address_qZ0Z_14\ : std_logic;
signal \un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0\ : std_logic;
signal \un1_M_this_external_address_q_cry_13\ : std_logic;
signal \un1_M_this_external_address_q_cry_14\ : std_logic;
signal \un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_8_cascade_\ : std_logic;
signal \M_this_external_address_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_5_mZ0Z_8\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_8_mZ0Z_0_cascade_\ : std_logic;
signal \M_this_external_address_q_RNIE44V9Z0Z_0\ : std_logic;
signal \M_this_external_address_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_0\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_5_mZ0Z_9\ : std_logic;
signal \un1_M_this_external_address_q_cry_8_c_RNI09PBZ0\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_5_mZ0Z_11_cascade_\ : std_logic;
signal \un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_11\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_11\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_3_cascade_\ : std_logic;
signal \un1_M_this_external_address_q_cry_2_c_RNIKMIBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_8_mZ0Z_3\ : std_logic;
signal \M_this_data_count_q_s_0\ : std_logic;
signal \M_this_state_qZ0Z_10\ : std_logic;
signal \this_vga_signals.N_292_cascade_\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_2_sqmuxaZ0\ : std_logic;
signal \M_this_state_d88_9\ : std_logic;
signal \N_506\ : std_logic;
signal \N_509\ : std_logic;
signal \N_510_cascade_\ : std_logic;
signal \N_511\ : std_logic;
signal \N_512\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \bfn_23_17_0_\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_data_count_q_s_1\ : std_logic;
signal \M_this_data_count_q_cry_0\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_q_s_2\ : std_logic;
signal \M_this_data_count_q_cry_1\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_q_s_3\ : std_logic;
signal \M_this_data_count_q_cry_2\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \M_this_data_count_q_s_4\ : std_logic;
signal \M_this_data_count_q_cry_3\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_q_s_5\ : std_logic;
signal \M_this_data_count_q_cry_4\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \M_this_data_count_q_s_6\ : std_logic;
signal \M_this_data_count_q_cry_5\ : std_logic;
signal \M_this_data_count_q_cry_6\ : std_logic;
signal \M_this_data_count_q_cry_7\ : std_logic;
signal \bfn_23_18_0_\ : std_logic;
signal \M_this_data_count_q_cry_8\ : std_logic;
signal \M_this_data_count_q_cry_9\ : std_logic;
signal \M_this_data_count_q_cry_10\ : std_logic;
signal \M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_data_count_q_cry_12\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \M_this_data_count_q_cry_13\ : std_logic;
signal \M_this_data_count_q_cry_14\ : std_logic;
signal \M_this_map_ram_read_data_6\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_12\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_1\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_8_mZ0Z_1_cascade_\ : std_logic;
signal \un1_M_this_external_address_q_cry_0_c_RNIGGGBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_2\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_8_mZ0Z_2_cascade_\ : std_logic;
signal \un1_M_this_external_address_q_cry_1_c_RNIIJHBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_8_mZ0Z_4\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_4\ : std_logic;
signal \un1_M_this_external_address_q_cry_3_c_RNIMPJBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_5_i_mZ0Z_15_cascade_\ : std_logic;
signal \un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_15\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_i_mZ0Z_15\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_7\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_8_mZ0Z_7_cascade_\ : std_logic;
signal \un1_M_this_external_address_q_cry_6_c_RNIS2NBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_5_mZ0Z_10_cascade_\ : std_logic;
signal \un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_10\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_10\ : std_logic;
signal \M_this_external_address_qZ0Z_9\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_9\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_5_mZ0Z_12\ : std_logic;
signal \this_vga_signals.un1_M_this_state_q_21_0\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_mZ0Z_12\ : std_logic;
signal \un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_12\ : std_logic;
signal \M_this_map_ram_write_data_3\ : std_logic;
signal \M_this_state_qZ0Z_13\ : std_logic;
signal \N_391_0\ : std_logic;
signal \this_vga_signals.un1_M_this_state_q_18Z0Z_1\ : std_logic;
signal \M_this_state_qZ0Z_11\ : std_logic;
signal \this_vga_signals.N_387_0\ : std_logic;
signal \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0\ : std_logic;
signal \N_513\ : std_logic;
signal \M_this_data_count_q_s_7\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \M_this_data_count_q_s_8\ : std_logic;
signal \N_514_cascade_\ : std_logic;
signal \M_this_data_count_q_s_9\ : std_logic;
signal \N_515_cascade_\ : std_logic;
signal \M_this_data_count_q_s_11\ : std_logic;
signal \M_this_data_count_q_s_12\ : std_logic;
signal \N_518_cascade_\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \M_this_data_count_q_s_14\ : std_logic;
signal \N_520_cascade_\ : std_logic;
signal \M_this_data_count_qZ0Z_14\ : std_logic;
signal \M_this_data_count_q_s_15\ : std_logic;
signal \N_521_cascade_\ : std_logic;
signal \M_this_data_count_qZ0Z_15\ : std_logic;
signal \N_517\ : std_logic;
signal \this_vga_signals.M_this_data_count_q_3_bmZ0Z_10\ : std_logic;
signal \M_this_data_count_q_cry_9_THRU_CO\ : std_logic;
signal \M_this_data_count_q_3_10_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_8\ : std_logic;
signal \N_389_0\ : std_logic;
signal \M_this_reset_cond_out_g_0\ : std_logic;
signal \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8_cascade_\ : std_logic;
signal \this_vga_signals.M_this_data_count_q_3_bmZ0Z_13\ : std_logic;
signal \this_vga_signals.M_this_data_count_q_3_amZ0Z_13_cascade_\ : std_logic;
signal \M_this_data_count_q_3_sn_N_2\ : std_logic;
signal \M_this_data_count_q_cry_12_THRU_CO\ : std_logic;
signal \M_this_data_count_q_3_13_cascade_\ : std_logic;
signal \N_570_0_i\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal clk_0_c_g : std_logic;
signal \M_this_data_count_qe_0_i\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \M_this_state_d88_10\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8\ : std_logic;
signal \this_vga_signals.M_this_data_count_q_3_amZ0Z_10\ : std_logic;
signal \M_this_map_ram_write_data_6\ : std_logic;
signal \M_this_map_ram_write_data_7\ : std_logic;
signal \this_ppu.M_haddress_qZ0Z_7\ : std_logic;
signal \M_this_ppu_map_addr_4\ : std_logic;
signal \M_this_ppu_vram_addr_6\ : std_logic;
signal \M_this_ppu_vram_addr_i_6\ : std_logic;
signal \M_this_map_ram_write_data_2\ : std_logic;
signal \M_this_map_ram_write_data_1\ : std_logic;
signal \M_this_map_ram_write_data_0\ : std_logic;
signal \M_this_map_ram_write_data_5\ : std_logic;
signal \M_this_map_ram_write_en_0\ : std_logic;
signal \M_this_map_ram_write_data_4\ : std_logic;
signal port_data_c_3 : std_logic;
signal port_data_c_2 : std_logic;
signal \this_vga_signals.M_this_external_address_d21Z0Z_2_cascade_\ : std_logic;
signal \this_vga_signals.M_this_external_address_dZ0Z21\ : std_logic;
signal port_data_c_1 : std_logic;
signal \this_vga_signals.M_this_external_address_d21Z0Z_2\ : std_logic;
signal port_data_c_0 : std_logic;
signal \this_vga_signals.M_this_external_address_dZ0Z22\ : std_logic;
signal port_data_c_5 : std_logic;
signal port_data_c_6 : std_logic;
signal port_data_c_7 : std_logic;
signal port_data_c_4 : std_logic;
signal \this_vga_signals.M_this_external_address_d21Z0Z_6\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_map_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    led <= led_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \M_this_ppu_sprites_addr_9\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_ppu_sprites_addr_8\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_ppu_sprites_addr_7\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_ppu_sprites_addr_6\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&\N__21433\&\N__23860\&\N__21574\&\N__20539\&\N__20506\&\N__33160\&\N__33094\&\N__25120\&\N__23595\&\N__23959\;
    \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&\N__25234\&\N__27676\&\N__25171\&\N__24697\&\N__24748\&\N__26518\&\N__26593\&\N__24808\&\N__26647\&\N__26119\;
    \this_map_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&\N__30400\&'0'&'0'&'0'&\N__33073\&'0'&'0'&'0'&\N__33067\&'0'&'0'&'0'&\N__33058\&'0';
    \M_this_map_ram_read_data_7\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_6\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_5\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_4\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&\N__21427\&\N__23854\&\N__21568\&\N__20533\&\N__20500\&\N__33154\&\N__33088\&\N__25113\&\N__23583\&\N__23949\;
    \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&\N__25228\&\N__27670\&\N__25165\&\N__24691\&\N__24742\&\N__26512\&\N__26587\&\N__24802\&\N__26641\&\N__26113\;
    \this_map_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&\N__33187\&'0'&'0'&'0'&\N__31471\&'0'&'0'&'0'&\N__33052\&'0'&'0'&'0'&\N__32947\&'0';
    \this_sprites_ram.mem_out_bus0_1\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_0\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__11326\&\N__11773\&\N__11665\&\N__11551\&\N__11437\&\N__20455\&\N__15613\&\N__15763\&\N__23545\&\N__22177\&\N__22372\;
    \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__22819\&\N__22966\&\N__23113\&\N__24340\&\N__23812\&\N__24973\&\N__26263\&\N__28366\&\N__22618\&\N__25618\&\N__26062\;
    \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21297\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21388\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus0_3\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_2\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__11320\&\N__11767\&\N__11659\&\N__11545\&\N__11431\&\N__20449\&\N__15607\&\N__15757\&\N__23539\&\N__22171\&\N__22366\;
    \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__22813\&\N__22960\&\N__23107\&\N__24334\&\N__23806\&\N__24967\&\N__26257\&\N__28360\&\N__22612\&\N__25612\&\N__26056\;
    \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21089\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21195\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_1\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_0\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__11314\&\N__11761\&\N__11653\&\N__11539\&\N__11425\&\N__20443\&\N__15601\&\N__15751\&\N__23533\&\N__22165\&\N__22360\;
    \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__22807\&\N__22954\&\N__23101\&\N__24328\&\N__23800\&\N__24961\&\N__26251\&\N__28354\&\N__22606\&\N__25606\&\N__26050\;
    \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21289\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21383\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_3\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_2\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__11308\&\N__11755\&\N__11647\&\N__11533\&\N__11419\&\N__20437\&\N__15595\&\N__15745\&\N__23527\&\N__22159\&\N__22354\;
    \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__22801\&\N__22948\&\N__23095\&\N__24322\&\N__23794\&\N__24955\&\N__26245\&\N__28348\&\N__22600\&\N__25600\&\N__26044\;
    \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21077\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21182\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_1\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_0\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__11302\&\N__11749\&\N__11641\&\N__11527\&\N__11413\&\N__20431\&\N__15589\&\N__15739\&\N__23521\&\N__22153\&\N__22348\;
    \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__22795\&\N__22942\&\N__23089\&\N__24316\&\N__23788\&\N__24949\&\N__26239\&\N__28342\&\N__22594\&\N__25594\&\N__26038\;
    \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21275\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21372\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_3\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_2\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__11296\&\N__11743\&\N__11635\&\N__11521\&\N__11407\&\N__20425\&\N__15583\&\N__15733\&\N__23515\&\N__22147\&\N__22342\;
    \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__22789\&\N__22936\&\N__23083\&\N__24310\&\N__23782\&\N__24943\&\N__26233\&\N__28336\&\N__22588\&\N__25588\&\N__26032\;
    \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21090\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21196\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_1\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_0\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__11290\&\N__11737\&\N__11629\&\N__11515\&\N__11401\&\N__20419\&\N__15577\&\N__15727\&\N__23509\&\N__22141\&\N__22336\;
    \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__22783\&\N__22930\&\N__23077\&\N__24304\&\N__23776\&\N__24937\&\N__26227\&\N__28330\&\N__22582\&\N__25582\&\N__26026\;
    \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21252\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21355\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_3\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_2\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__11284\&\N__11731\&\N__11623\&\N__11509\&\N__11395\&\N__20413\&\N__15571\&\N__15721\&\N__23503\&\N__22135\&\N__22330\;
    \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__22777\&\N__22924\&\N__23071\&\N__24298\&\N__23770\&\N__24931\&\N__26221\&\N__28324\&\N__22576\&\N__25576\&\N__26020\;
    \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21081\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21177\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_1\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_0\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__11278\&\N__11725\&\N__11617\&\N__11503\&\N__11389\&\N__20407\&\N__15565\&\N__15715\&\N__23497\&\N__22129\&\N__22324\;
    \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__22771\&\N__22918\&\N__23065\&\N__24292\&\N__23764\&\N__24925\&\N__26215\&\N__28318\&\N__22570\&\N__25570\&\N__26014\;
    \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21237\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21346\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_3\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_2\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__11272\&\N__11719\&\N__11611\&\N__11497\&\N__11383\&\N__20401\&\N__15559\&\N__15709\&\N__23491\&\N__22123\&\N__22318\;
    \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__22765\&\N__22912\&\N__23059\&\N__24286\&\N__23758\&\N__24919\&\N__26209\&\N__28312\&\N__22564\&\N__25564\&\N__26008\;
    \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21049\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21181\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_1\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_0\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__11266\&\N__11713\&\N__11605\&\N__11491\&\N__11377\&\N__20395\&\N__15553\&\N__15703\&\N__23485\&\N__22117\&\N__22312\;
    \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__22759\&\N__22906\&\N__23053\&\N__24280\&\N__23752\&\N__24913\&\N__26203\&\N__28306\&\N__22558\&\N__25558\&\N__26002\;
    \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21282\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21365\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_3\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_2\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__11260\&\N__11707\&\N__11599\&\N__11485\&\N__11371\&\N__20389\&\N__15547\&\N__15697\&\N__23479\&\N__22111\&\N__22306\;
    \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__22753\&\N__22900\&\N__23047\&\N__24274\&\N__23746\&\N__24907\&\N__26197\&\N__28300\&\N__22552\&\N__25552\&\N__25996\;
    \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21070\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21197\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_1\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_0\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__11254\&\N__11701\&\N__11593\&\N__11479\&\N__11365\&\N__20383\&\N__15541\&\N__15691\&\N__23473\&\N__22105\&\N__22300\;
    \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__22747\&\N__22894\&\N__23041\&\N__24268\&\N__23740\&\N__24901\&\N__26191\&\N__28294\&\N__22546\&\N__25546\&\N__25990\;
    \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21293\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21379\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_3\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_2\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__11248\&\N__11695\&\N__11587\&\N__11473\&\N__11359\&\N__20377\&\N__15535\&\N__15685\&\N__23467\&\N__22099\&\N__22294\;
    \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__22741\&\N__22888\&\N__23035\&\N__24262\&\N__23734\&\N__24895\&\N__26185\&\N__28288\&\N__22540\&\N__25540\&\N__25984\;
    \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21085\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21198\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_1\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_0\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__11242\&\N__11689\&\N__11581\&\N__11467\&\N__11353\&\N__20371\&\N__15529\&\N__15678\&\N__23461\&\N__22093\&\N__22288\;
    \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__22735\&\N__22882\&\N__23029\&\N__24256\&\N__23728\&\N__24889\&\N__26179\&\N__28282\&\N__22534\&\N__25534\&\N__25978\;
    \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21298\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21387\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_3\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_2\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__11236\&\N__11683\&\N__11575\&\N__11461\&\N__11347\&\N__20365\&\N__15523\&\N__15666\&\N__23455\&\N__22087\&\N__22281\;
    \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__22729\&\N__22876\&\N__23023\&\N__24250\&\N__23722\&\N__24883\&\N__26173\&\N__28276\&\N__22528\&\N__25528\&\N__25972\;
    \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21091\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21202\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__18607\&\N__14278\&\N__20893\&\N__13963\&\N__14353\&\N__13900\&\N__12184\&\N__12625\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__15681\&\N__33139\&\N__25116\&\N__23596\&\N__23958\&\N__23454\&\N__22086\&\N__22284\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__13720\&\N__20635\&\N__19912\&\N__16894\;

    \this_map_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32057\,
            RE => \N__30145\,
            WCLKE => \N__33044\,
            WCLK => \N__32058\,
            WE => \N__30156\
        );

    \this_map_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32061\,
            RE => \N__30160\,
            WCLKE => \N__33045\,
            WCLK => \N__32062\,
            WE => \N__30155\
        );

    \this_sprites_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__31937\,
            RE => \N__30039\,
            WCLKE => \N__20866\,
            WCLK => \N__31938\,
            WE => \N__30041\
        );

    \this_sprites_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__31939\,
            RE => \N__30038\,
            WCLKE => \N__20862\,
            WCLK => \N__31940\,
            WE => \N__30040\
        );

    \this_sprites_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__31942\,
            RE => \N__29948\,
            WCLKE => \N__20836\,
            WCLK => \N__31943\,
            WE => \N__30042\
        );

    \this_sprites_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__31947\,
            RE => \N__29947\,
            WCLKE => \N__20832\,
            WCLK => \N__31948\,
            WE => \N__29961\
        );

    \this_sprites_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__31960\,
            RE => \N__29848\,
            WCLKE => \N__20752\,
            WCLK => \N__31959\,
            WE => \N__29962\
        );

    \this_sprites_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__31970\,
            RE => \N__29836\,
            WCLKE => \N__20751\,
            WCLK => \N__31971\,
            WE => \N__29766\
        );

    \this_sprites_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__31985\,
            RE => \N__29869\,
            WCLKE => \N__15403\,
            WCLK => \N__31986\,
            WE => \N__29935\
        );

    \this_sprites_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__31999\,
            RE => \N__29876\,
            WCLKE => \N__15402\,
            WCLK => \N__32000\,
            WE => \N__30030\
        );

    \this_sprites_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32013\,
            RE => \N__29966\,
            WCLKE => \N__14334\,
            WCLK => \N__32014\,
            WE => \N__30031\
        );

    \this_sprites_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32030\,
            RE => \N__29967\,
            WCLKE => \N__14338\,
            WCLK => \N__32031\,
            WE => \N__30085\
        );

    \this_sprites_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32042\,
            RE => \N__30043\,
            WCLKE => \N__14445\,
            WCLK => \N__32043\,
            WE => \N__30054\
        );

    \this_sprites_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32049\,
            RE => \N__30044\,
            WCLKE => \N__14446\,
            WCLK => \N__32050\,
            WE => \N__30089\
        );

    \this_sprites_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32051\,
            RE => \N__30090\,
            WCLKE => \N__15792\,
            WCLK => \N__32052\,
            WE => \N__30092\
        );

    \this_sprites_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32053\,
            RE => \N__30091\,
            WCLKE => \N__15793\,
            WCLK => \N__32054\,
            WE => \N__30093\
        );

    \this_sprites_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32055\,
            RE => \N__30115\,
            WCLKE => \N__20556\,
            WCLK => \N__32056\,
            WE => \N__30117\
        );

    \this_sprites_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32059\,
            RE => \N__30116\,
            WCLKE => \N__20563\,
            WCLK => \N__32060\,
            WE => \N__30118\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32023\,
            RE => \N__30078\,
            WCLKE => \N__22225\,
            WCLK => \N__32024\,
            WE => \N__30106\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__34841\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34843\,
            DIN => \N__34842\,
            DOUT => \N__34841\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34843\,
            PADOUT => \N__34842\,
            PADIN => \N__34841\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34832\,
            DIN => \N__34831\,
            DOUT => \N__34830\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34832\,
            PADOUT => \N__34831\,
            PADIN => \N__34830\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34823\,
            DIN => \N__34822\,
            DOUT => \N__34821\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34823\,
            PADOUT => \N__34822\,
            PADIN => \N__34821\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34814\,
            DIN => \N__34813\,
            DOUT => \N__34812\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34814\,
            PADOUT => \N__34813\,
            PADIN => \N__34812\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12025\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34805\,
            DIN => \N__34804\,
            DOUT => \N__34803\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34805\,
            PADOUT => \N__34804\,
            PADIN => \N__34803\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11881\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34796\,
            DIN => \N__34795\,
            DOUT => \N__34794\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34796\,
            PADOUT => \N__34795\,
            PADIN => \N__34794\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29934\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34787\,
            DIN => \N__34786\,
            DOUT => \N__34785\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34787\,
            PADOUT => \N__34786\,
            PADIN => \N__34785\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__28585\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34778\,
            DIN => \N__34777\,
            DOUT => \N__34776\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34778\,
            PADOUT => \N__34777\,
            PADIN => \N__34776\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34769\,
            DIN => \N__34768\,
            DOUT => \N__34767\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34769\,
            PADOUT => \N__34768\,
            PADIN => \N__34767\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34760\,
            DIN => \N__34759\,
            DOUT => \N__34758\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34760\,
            PADOUT => \N__34759\,
            PADIN => \N__34758\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34751\,
            DIN => \N__34750\,
            DOUT => \N__34749\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34751\,
            PADOUT => \N__34750\,
            PADIN => \N__34749\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34742\,
            DIN => \N__34741\,
            DOUT => \N__34740\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34742\,
            PADOUT => \N__34741\,
            PADIN => \N__34740\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34733\,
            DIN => \N__34732\,
            DOUT => \N__34731\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34733\,
            PADOUT => \N__34732\,
            PADIN => \N__34731\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34724\,
            DIN => \N__34723\,
            DOUT => \N__34722\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34724\,
            PADOUT => \N__34723\,
            PADIN => \N__34722\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__28984\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21734\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34715\,
            DIN => \N__34714\,
            DOUT => \N__34713\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34715\,
            PADOUT => \N__34714\,
            PADIN => \N__34713\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__30376\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21867\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34706\,
            DIN => \N__34705\,
            DOUT => \N__34704\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34706\,
            PADOUT => \N__34705\,
            PADIN => \N__34704\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__30316\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21839\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34697\,
            DIN => \N__34696\,
            DOUT => \N__34695\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34697\,
            PADOUT => \N__34696\,
            PADIN => \N__34695\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__29251\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21866\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34688\,
            DIN => \N__34687\,
            DOUT => \N__34686\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34688\,
            PADOUT => \N__34687\,
            PADIN => \N__34686\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__30247\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21853\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34679\,
            DIN => \N__34678\,
            DOUT => \N__34677\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34679\,
            PADOUT => \N__34678\,
            PADIN => \N__34677\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__28753\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21826\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34670\,
            DIN => \N__34669\,
            DOUT => \N__34668\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34670\,
            PADOUT => \N__34669\,
            PADIN => \N__34668\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__28708\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21743\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34661\,
            DIN => \N__34660\,
            DOUT => \N__34659\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34661\,
            PADOUT => \N__34660\,
            PADIN => \N__34659\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__30994\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21775\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34652\,
            DIN => \N__34651\,
            DOUT => \N__34650\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34652\,
            PADOUT => \N__34651\,
            PADIN => \N__34650\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__30940\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21810\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34643\,
            DIN => \N__34642\,
            DOUT => \N__34641\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34643\,
            PADOUT => \N__34642\,
            PADIN => \N__34641\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29305\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21871\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34634\,
            DIN => \N__34633\,
            DOUT => \N__34632\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34634\,
            PADOUT => \N__34633\,
            PADIN => \N__34632\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__30436\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21854\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34625\,
            DIN => \N__34624\,
            DOUT => \N__34623\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34625\,
            PADOUT => \N__34624\,
            PADIN => \N__34623\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__28894\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21852\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34616\,
            DIN => \N__34615\,
            DOUT => \N__34614\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34616\,
            PADOUT => \N__34615\,
            PADIN => \N__34614\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__28849\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21822\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34607\,
            DIN => \N__34606\,
            DOUT => \N__34605\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34607\,
            PADOUT => \N__34606\,
            PADIN => \N__34605\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__30205\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21865\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34598\,
            DIN => \N__34597\,
            DOUT => \N__34596\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34598\,
            PADOUT => \N__34597\,
            PADIN => \N__34596\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29038\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21809\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34589\,
            DIN => \N__34588\,
            DOUT => \N__34587\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34589\,
            PADOUT => \N__34588\,
            PADIN => \N__34587\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__30901\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21858\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34580\,
            DIN => \N__34579\,
            DOUT => \N__34578\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34580\,
            PADOUT => \N__34579\,
            PADIN => \N__34578\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34571\,
            DIN => \N__34570\,
            DOUT => \N__34569\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34571\,
            PADOUT => \N__34570\,
            PADIN => \N__34569\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34562\,
            DIN => \N__34561\,
            DOUT => \N__34560\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34562\,
            PADOUT => \N__34561\,
            PADIN => \N__34560\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34553\,
            DIN => \N__34552\,
            DOUT => \N__34551\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34553\,
            PADOUT => \N__34552\,
            PADIN => \N__34551\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34544\,
            DIN => \N__34543\,
            DOUT => \N__34542\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34544\,
            PADOUT => \N__34543\,
            PADIN => \N__34542\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34535\,
            DIN => \N__34534\,
            DOUT => \N__34533\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34535\,
            PADOUT => \N__34534\,
            PADIN => \N__34533\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34526\,
            DIN => \N__34525\,
            DOUT => \N__34524\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34526\,
            PADOUT => \N__34525\,
            PADIN => \N__34524\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34517\,
            DIN => \N__34516\,
            DOUT => \N__34515\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34517\,
            PADOUT => \N__34516\,
            PADIN => \N__34515\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34508\,
            DIN => \N__34507\,
            DOUT => \N__34506\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34508\,
            PADOUT => \N__34507\,
            PADIN => \N__34506\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34499\,
            DIN => \N__34498\,
            DOUT => \N__34497\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34499\,
            PADOUT => \N__34498\,
            PADIN => \N__34497\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11812\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34490\,
            DIN => \N__34489\,
            DOUT => \N__34488\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34490\,
            PADOUT => \N__34489\,
            PADIN => \N__34488\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21898\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34481\,
            DIN => \N__34480\,
            DOUT => \N__34479\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34481\,
            PADOUT => \N__34480\,
            PADIN => \N__34479\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34472\,
            DIN => \N__34471\,
            DOUT => \N__34470\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34472\,
            PADOUT => \N__34471\,
            PADIN => \N__34470\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11863\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34463\,
            DIN => \N__34462\,
            DOUT => \N__34461\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__34463\,
            PADOUT => \N__34462\,
            PADIN => \N__34461\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__30144\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21848\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34454\,
            DIN => \N__34453\,
            DOUT => \N__34452\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34454\,
            PADOUT => \N__34453\,
            PADIN => \N__34452\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11797\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34445\,
            DIN => \N__34444\,
            DOUT => \N__34443\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34445\,
            PADOUT => \N__34444\,
            PADIN => \N__34443\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11782\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34436\,
            DIN => \N__34435\,
            DOUT => \N__34434\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34436\,
            PADOUT => \N__34435\,
            PADIN => \N__34434\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11917\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34427\,
            DIN => \N__34426\,
            DOUT => \N__34425\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34427\,
            PADOUT => \N__34426\,
            PADIN => \N__34425\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11965\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34418\,
            DIN => \N__34417\,
            DOUT => \N__34416\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34418\,
            PADOUT => \N__34417\,
            PADIN => \N__34416\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11950\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34409\,
            DIN => \N__34408\,
            DOUT => \N__34407\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34409\,
            PADOUT => \N__34408\,
            PADIN => \N__34407\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11830\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34400\,
            DIN => \N__34399\,
            DOUT => \N__34398\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__34400\,
            PADOUT => \N__34399\,
            PADIN => \N__34398\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34391\,
            DIN => \N__34390\,
            DOUT => \N__34389\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34391\,
            PADOUT => \N__34390\,
            PADIN => \N__34389\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12223\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34382\,
            DIN => \N__34381\,
            DOUT => \N__34380\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__34382\,
            PADOUT => \N__34381\,
            PADIN => \N__34380\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12469\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__8553\ : CascadeMux
    port map (
            O => \N__34363\,
            I => \N__34359\
        );

    \I__8552\ : CascadeMux
    port map (
            O => \N__34362\,
            I => \N__34354\
        );

    \I__8551\ : InMux
    port map (
            O => \N__34359\,
            I => \N__34351\
        );

    \I__8550\ : InMux
    port map (
            O => \N__34358\,
            I => \N__34348\
        );

    \I__8549\ : InMux
    port map (
            O => \N__34357\,
            I => \N__34344\
        );

    \I__8548\ : InMux
    port map (
            O => \N__34354\,
            I => \N__34340\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__34351\,
            I => \N__34337\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__34348\,
            I => \N__34334\
        );

    \I__8545\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34328\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__34344\,
            I => \N__34325\
        );

    \I__8543\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34322\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__34340\,
            I => \N__34319\
        );

    \I__8541\ : Span4Mux_v
    port map (
            O => \N__34337\,
            I => \N__34313\
        );

    \I__8540\ : Span4Mux_v
    port map (
            O => \N__34334\,
            I => \N__34313\
        );

    \I__8539\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34310\
        );

    \I__8538\ : CascadeMux
    port map (
            O => \N__34332\,
            I => \N__34307\
        );

    \I__8537\ : CascadeMux
    port map (
            O => \N__34331\,
            I => \N__34303\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__34328\,
            I => \N__34300\
        );

    \I__8535\ : Span4Mux_v
    port map (
            O => \N__34325\,
            I => \N__34297\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__34322\,
            I => \N__34294\
        );

    \I__8533\ : Span4Mux_v
    port map (
            O => \N__34319\,
            I => \N__34291\
        );

    \I__8532\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34288\
        );

    \I__8531\ : Sp12to4
    port map (
            O => \N__34313\,
            I => \N__34285\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__34310\,
            I => \N__34282\
        );

    \I__8529\ : InMux
    port map (
            O => \N__34307\,
            I => \N__34279\
        );

    \I__8528\ : InMux
    port map (
            O => \N__34306\,
            I => \N__34274\
        );

    \I__8527\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34274\
        );

    \I__8526\ : Sp12to4
    port map (
            O => \N__34300\,
            I => \N__34271\
        );

    \I__8525\ : Span4Mux_h
    port map (
            O => \N__34297\,
            I => \N__34266\
        );

    \I__8524\ : Span4Mux_h
    port map (
            O => \N__34294\,
            I => \N__34266\
        );

    \I__8523\ : Span4Mux_v
    port map (
            O => \N__34291\,
            I => \N__34261\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__34288\,
            I => \N__34261\
        );

    \I__8521\ : Span12Mux_h
    port map (
            O => \N__34285\,
            I => \N__34258\
        );

    \I__8520\ : Span12Mux_v
    port map (
            O => \N__34282\,
            I => \N__34251\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__34279\,
            I => \N__34251\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__34274\,
            I => \N__34251\
        );

    \I__8517\ : Span12Mux_h
    port map (
            O => \N__34271\,
            I => \N__34246\
        );

    \I__8516\ : Sp12to4
    port map (
            O => \N__34266\,
            I => \N__34246\
        );

    \I__8515\ : Span4Mux_h
    port map (
            O => \N__34261\,
            I => \N__34243\
        );

    \I__8514\ : Span12Mux_v
    port map (
            O => \N__34258\,
            I => \N__34240\
        );

    \I__8513\ : Span12Mux_h
    port map (
            O => \N__34251\,
            I => \N__34237\
        );

    \I__8512\ : Span12Mux_v
    port map (
            O => \N__34246\,
            I => \N__34234\
        );

    \I__8511\ : Span4Mux_h
    port map (
            O => \N__34243\,
            I => \N__34231\
        );

    \I__8510\ : Odrv12
    port map (
            O => \N__34240\,
            I => port_data_c_3
        );

    \I__8509\ : Odrv12
    port map (
            O => \N__34237\,
            I => port_data_c_3
        );

    \I__8508\ : Odrv12
    port map (
            O => \N__34234\,
            I => port_data_c_3
        );

    \I__8507\ : Odrv4
    port map (
            O => \N__34231\,
            I => port_data_c_3
        );

    \I__8506\ : CascadeMux
    port map (
            O => \N__34222\,
            I => \N__34217\
        );

    \I__8505\ : CascadeMux
    port map (
            O => \N__34221\,
            I => \N__34214\
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__34220\,
            I => \N__34209\
        );

    \I__8503\ : InMux
    port map (
            O => \N__34217\,
            I => \N__34206\
        );

    \I__8502\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34203\
        );

    \I__8501\ : CascadeMux
    port map (
            O => \N__34213\,
            I => \N__34199\
        );

    \I__8500\ : InMux
    port map (
            O => \N__34212\,
            I => \N__34196\
        );

    \I__8499\ : InMux
    port map (
            O => \N__34209\,
            I => \N__34193\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__34206\,
            I => \N__34189\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__34203\,
            I => \N__34186\
        );

    \I__8496\ : CascadeMux
    port map (
            O => \N__34202\,
            I => \N__34183\
        );

    \I__8495\ : InMux
    port map (
            O => \N__34199\,
            I => \N__34180\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__34196\,
            I => \N__34177\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__34193\,
            I => \N__34174\
        );

    \I__8492\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34171\
        );

    \I__8491\ : Span4Mux_v
    port map (
            O => \N__34189\,
            I => \N__34166\
        );

    \I__8490\ : Span4Mux_v
    port map (
            O => \N__34186\,
            I => \N__34166\
        );

    \I__8489\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34163\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__34180\,
            I => \N__34160\
        );

    \I__8487\ : Span4Mux_h
    port map (
            O => \N__34177\,
            I => \N__34155\
        );

    \I__8486\ : Span4Mux_v
    port map (
            O => \N__34174\,
            I => \N__34155\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__34171\,
            I => \N__34152\
        );

    \I__8484\ : Span4Mux_h
    port map (
            O => \N__34166\,
            I => \N__34145\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__34163\,
            I => \N__34145\
        );

    \I__8482\ : Span4Mux_v
    port map (
            O => \N__34160\,
            I => \N__34141\
        );

    \I__8481\ : Span4Mux_h
    port map (
            O => \N__34155\,
            I => \N__34136\
        );

    \I__8480\ : Span4Mux_v
    port map (
            O => \N__34152\,
            I => \N__34136\
        );

    \I__8479\ : InMux
    port map (
            O => \N__34151\,
            I => \N__34133\
        );

    \I__8478\ : CascadeMux
    port map (
            O => \N__34150\,
            I => \N__34130\
        );

    \I__8477\ : Span4Mux_h
    port map (
            O => \N__34145\,
            I => \N__34126\
        );

    \I__8476\ : InMux
    port map (
            O => \N__34144\,
            I => \N__34123\
        );

    \I__8475\ : Sp12to4
    port map (
            O => \N__34141\,
            I => \N__34120\
        );

    \I__8474\ : Span4Mux_h
    port map (
            O => \N__34136\,
            I => \N__34115\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__34133\,
            I => \N__34115\
        );

    \I__8472\ : InMux
    port map (
            O => \N__34130\,
            I => \N__34112\
        );

    \I__8471\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34109\
        );

    \I__8470\ : Span4Mux_v
    port map (
            O => \N__34126\,
            I => \N__34106\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__34123\,
            I => \N__34103\
        );

    \I__8468\ : Span12Mux_h
    port map (
            O => \N__34120\,
            I => \N__34100\
        );

    \I__8467\ : Sp12to4
    port map (
            O => \N__34115\,
            I => \N__34097\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__34112\,
            I => \N__34092\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__34109\,
            I => \N__34092\
        );

    \I__8464\ : Span4Mux_v
    port map (
            O => \N__34106\,
            I => \N__34087\
        );

    \I__8463\ : Span4Mux_h
    port map (
            O => \N__34103\,
            I => \N__34087\
        );

    \I__8462\ : Span12Mux_v
    port map (
            O => \N__34100\,
            I => \N__34084\
        );

    \I__8461\ : Span12Mux_v
    port map (
            O => \N__34097\,
            I => \N__34081\
        );

    \I__8460\ : Span12Mux_h
    port map (
            O => \N__34092\,
            I => \N__34078\
        );

    \I__8459\ : Span4Mux_v
    port map (
            O => \N__34087\,
            I => \N__34075\
        );

    \I__8458\ : Odrv12
    port map (
            O => \N__34084\,
            I => port_data_c_2
        );

    \I__8457\ : Odrv12
    port map (
            O => \N__34081\,
            I => port_data_c_2
        );

    \I__8456\ : Odrv12
    port map (
            O => \N__34078\,
            I => port_data_c_2
        );

    \I__8455\ : Odrv4
    port map (
            O => \N__34075\,
            I => port_data_c_2
        );

    \I__8454\ : CascadeMux
    port map (
            O => \N__34066\,
            I => \this_vga_signals.M_this_external_address_d21Z0Z_2_cascade_\
        );

    \I__8453\ : CascadeMux
    port map (
            O => \N__34063\,
            I => \N__34060\
        );

    \I__8452\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34054\
        );

    \I__8451\ : CascadeMux
    port map (
            O => \N__34059\,
            I => \N__34051\
        );

    \I__8450\ : InMux
    port map (
            O => \N__34058\,
            I => \N__34047\
        );

    \I__8449\ : InMux
    port map (
            O => \N__34057\,
            I => \N__34044\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__34054\,
            I => \N__34041\
        );

    \I__8447\ : InMux
    port map (
            O => \N__34051\,
            I => \N__34038\
        );

    \I__8446\ : CascadeMux
    port map (
            O => \N__34050\,
            I => \N__34035\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__34047\,
            I => \N__34032\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__34044\,
            I => \N__34029\
        );

    \I__8443\ : Span4Mux_h
    port map (
            O => \N__34041\,
            I => \N__34024\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__34038\,
            I => \N__34024\
        );

    \I__8441\ : InMux
    port map (
            O => \N__34035\,
            I => \N__34021\
        );

    \I__8440\ : Span12Mux_h
    port map (
            O => \N__34032\,
            I => \N__34018\
        );

    \I__8439\ : Span12Mux_h
    port map (
            O => \N__34029\,
            I => \N__34015\
        );

    \I__8438\ : Span4Mux_h
    port map (
            O => \N__34024\,
            I => \N__34012\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__34021\,
            I => \N__34009\
        );

    \I__8436\ : Odrv12
    port map (
            O => \N__34018\,
            I => \this_vga_signals.M_this_external_address_dZ0Z21\
        );

    \I__8435\ : Odrv12
    port map (
            O => \N__34015\,
            I => \this_vga_signals.M_this_external_address_dZ0Z21\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__34012\,
            I => \this_vga_signals.M_this_external_address_dZ0Z21\
        );

    \I__8433\ : Odrv12
    port map (
            O => \N__34009\,
            I => \this_vga_signals.M_this_external_address_dZ0Z21\
        );

    \I__8432\ : InMux
    port map (
            O => \N__34000\,
            I => \N__33996\
        );

    \I__8431\ : InMux
    port map (
            O => \N__33999\,
            I => \N__33993\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__33996\,
            I => \N__33986\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__33993\,
            I => \N__33983\
        );

    \I__8428\ : CascadeMux
    port map (
            O => \N__33992\,
            I => \N__33978\
        );

    \I__8427\ : CascadeMux
    port map (
            O => \N__33991\,
            I => \N__33975\
        );

    \I__8426\ : CascadeMux
    port map (
            O => \N__33990\,
            I => \N__33972\
        );

    \I__8425\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33967\
        );

    \I__8424\ : Span4Mux_h
    port map (
            O => \N__33986\,
            I => \N__33961\
        );

    \I__8423\ : Span4Mux_v
    port map (
            O => \N__33983\,
            I => \N__33961\
        );

    \I__8422\ : InMux
    port map (
            O => \N__33982\,
            I => \N__33958\
        );

    \I__8421\ : CascadeMux
    port map (
            O => \N__33981\,
            I => \N__33955\
        );

    \I__8420\ : InMux
    port map (
            O => \N__33978\,
            I => \N__33952\
        );

    \I__8419\ : InMux
    port map (
            O => \N__33975\,
            I => \N__33949\
        );

    \I__8418\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33946\
        );

    \I__8417\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33940\
        );

    \I__8416\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33940\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__33967\,
            I => \N__33937\
        );

    \I__8414\ : CascadeMux
    port map (
            O => \N__33966\,
            I => \N__33934\
        );

    \I__8413\ : Span4Mux_h
    port map (
            O => \N__33961\,
            I => \N__33929\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__33958\,
            I => \N__33929\
        );

    \I__8411\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33926\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__33952\,
            I => \N__33923\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__33949\,
            I => \N__33918\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__33946\,
            I => \N__33918\
        );

    \I__8407\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33915\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__33940\,
            I => \N__33912\
        );

    \I__8405\ : Span4Mux_v
    port map (
            O => \N__33937\,
            I => \N__33909\
        );

    \I__8404\ : InMux
    port map (
            O => \N__33934\,
            I => \N__33906\
        );

    \I__8403\ : Span4Mux_h
    port map (
            O => \N__33929\,
            I => \N__33901\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__33926\,
            I => \N__33901\
        );

    \I__8401\ : Span4Mux_v
    port map (
            O => \N__33923\,
            I => \N__33898\
        );

    \I__8400\ : Span4Mux_v
    port map (
            O => \N__33918\,
            I => \N__33895\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__33915\,
            I => \N__33892\
        );

    \I__8398\ : Span12Mux_s7_h
    port map (
            O => \N__33912\,
            I => \N__33885\
        );

    \I__8397\ : Sp12to4
    port map (
            O => \N__33909\,
            I => \N__33885\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__33906\,
            I => \N__33885\
        );

    \I__8395\ : Span4Mux_v
    port map (
            O => \N__33901\,
            I => \N__33882\
        );

    \I__8394\ : Span4Mux_v
    port map (
            O => \N__33898\,
            I => \N__33875\
        );

    \I__8393\ : Span4Mux_v
    port map (
            O => \N__33895\,
            I => \N__33875\
        );

    \I__8392\ : Span4Mux_v
    port map (
            O => \N__33892\,
            I => \N__33875\
        );

    \I__8391\ : Span12Mux_h
    port map (
            O => \N__33885\,
            I => \N__33872\
        );

    \I__8390\ : Span4Mux_h
    port map (
            O => \N__33882\,
            I => \N__33869\
        );

    \I__8389\ : Sp12to4
    port map (
            O => \N__33875\,
            I => \N__33866\
        );

    \I__8388\ : Span12Mux_v
    port map (
            O => \N__33872\,
            I => \N__33863\
        );

    \I__8387\ : Sp12to4
    port map (
            O => \N__33869\,
            I => \N__33860\
        );

    \I__8386\ : Span12Mux_h
    port map (
            O => \N__33866\,
            I => \N__33857\
        );

    \I__8385\ : Odrv12
    port map (
            O => \N__33863\,
            I => port_data_c_1
        );

    \I__8384\ : Odrv12
    port map (
            O => \N__33860\,
            I => port_data_c_1
        );

    \I__8383\ : Odrv12
    port map (
            O => \N__33857\,
            I => port_data_c_1
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__33850\,
            I => \N__33847\
        );

    \I__8381\ : InMux
    port map (
            O => \N__33847\,
            I => \N__33844\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__33844\,
            I => \this_vga_signals.M_this_external_address_d21Z0Z_2\
        );

    \I__8379\ : CascadeMux
    port map (
            O => \N__33841\,
            I => \N__33838\
        );

    \I__8378\ : InMux
    port map (
            O => \N__33838\,
            I => \N__33832\
        );

    \I__8377\ : CascadeMux
    port map (
            O => \N__33837\,
            I => \N__33829\
        );

    \I__8376\ : CascadeMux
    port map (
            O => \N__33836\,
            I => \N__33824\
        );

    \I__8375\ : InMux
    port map (
            O => \N__33835\,
            I => \N__33819\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__33832\,
            I => \N__33815\
        );

    \I__8373\ : InMux
    port map (
            O => \N__33829\,
            I => \N__33808\
        );

    \I__8372\ : InMux
    port map (
            O => \N__33828\,
            I => \N__33808\
        );

    \I__8371\ : InMux
    port map (
            O => \N__33827\,
            I => \N__33803\
        );

    \I__8370\ : InMux
    port map (
            O => \N__33824\,
            I => \N__33803\
        );

    \I__8369\ : InMux
    port map (
            O => \N__33823\,
            I => \N__33798\
        );

    \I__8368\ : InMux
    port map (
            O => \N__33822\,
            I => \N__33798\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__33819\,
            I => \N__33795\
        );

    \I__8366\ : InMux
    port map (
            O => \N__33818\,
            I => \N__33791\
        );

    \I__8365\ : Span4Mux_v
    port map (
            O => \N__33815\,
            I => \N__33788\
        );

    \I__8364\ : InMux
    port map (
            O => \N__33814\,
            I => \N__33785\
        );

    \I__8363\ : InMux
    port map (
            O => \N__33813\,
            I => \N__33782\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__33808\,
            I => \N__33779\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__33803\,
            I => \N__33776\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__33798\,
            I => \N__33773\
        );

    \I__8359\ : Span4Mux_v
    port map (
            O => \N__33795\,
            I => \N__33770\
        );

    \I__8358\ : InMux
    port map (
            O => \N__33794\,
            I => \N__33767\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__33791\,
            I => \N__33764\
        );

    \I__8356\ : Span4Mux_v
    port map (
            O => \N__33788\,
            I => \N__33761\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__33785\,
            I => \N__33758\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__33782\,
            I => \N__33755\
        );

    \I__8353\ : Span4Mux_v
    port map (
            O => \N__33779\,
            I => \N__33752\
        );

    \I__8352\ : Span4Mux_v
    port map (
            O => \N__33776\,
            I => \N__33749\
        );

    \I__8351\ : Sp12to4
    port map (
            O => \N__33773\,
            I => \N__33742\
        );

    \I__8350\ : Sp12to4
    port map (
            O => \N__33770\,
            I => \N__33742\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__33767\,
            I => \N__33742\
        );

    \I__8348\ : Span4Mux_h
    port map (
            O => \N__33764\,
            I => \N__33739\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__33761\,
            I => \N__33736\
        );

    \I__8346\ : Span4Mux_v
    port map (
            O => \N__33758\,
            I => \N__33733\
        );

    \I__8345\ : Span12Mux_h
    port map (
            O => \N__33755\,
            I => \N__33730\
        );

    \I__8344\ : Sp12to4
    port map (
            O => \N__33752\,
            I => \N__33725\
        );

    \I__8343\ : Sp12to4
    port map (
            O => \N__33749\,
            I => \N__33725\
        );

    \I__8342\ : Span12Mux_h
    port map (
            O => \N__33742\,
            I => \N__33720\
        );

    \I__8341\ : Sp12to4
    port map (
            O => \N__33739\,
            I => \N__33720\
        );

    \I__8340\ : Sp12to4
    port map (
            O => \N__33736\,
            I => \N__33715\
        );

    \I__8339\ : Sp12to4
    port map (
            O => \N__33733\,
            I => \N__33715\
        );

    \I__8338\ : Span12Mux_v
    port map (
            O => \N__33730\,
            I => \N__33712\
        );

    \I__8337\ : Span12Mux_h
    port map (
            O => \N__33725\,
            I => \N__33709\
        );

    \I__8336\ : Span12Mux_v
    port map (
            O => \N__33720\,
            I => \N__33704\
        );

    \I__8335\ : Span12Mux_h
    port map (
            O => \N__33715\,
            I => \N__33704\
        );

    \I__8334\ : Odrv12
    port map (
            O => \N__33712\,
            I => port_data_c_0
        );

    \I__8333\ : Odrv12
    port map (
            O => \N__33709\,
            I => port_data_c_0
        );

    \I__8332\ : Odrv12
    port map (
            O => \N__33704\,
            I => port_data_c_0
        );

    \I__8331\ : CascadeMux
    port map (
            O => \N__33697\,
            I => \N__33694\
        );

    \I__8330\ : InMux
    port map (
            O => \N__33694\,
            I => \N__33689\
        );

    \I__8329\ : InMux
    port map (
            O => \N__33693\,
            I => \N__33686\
        );

    \I__8328\ : InMux
    port map (
            O => \N__33692\,
            I => \N__33683\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__33689\,
            I => \N__33679\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__33686\,
            I => \N__33676\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__33683\,
            I => \N__33673\
        );

    \I__8324\ : InMux
    port map (
            O => \N__33682\,
            I => \N__33670\
        );

    \I__8323\ : Span4Mux_v
    port map (
            O => \N__33679\,
            I => \N__33665\
        );

    \I__8322\ : Span4Mux_v
    port map (
            O => \N__33676\,
            I => \N__33665\
        );

    \I__8321\ : Span4Mux_v
    port map (
            O => \N__33673\,
            I => \N__33662\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__33670\,
            I => \N__33659\
        );

    \I__8319\ : Span4Mux_h
    port map (
            O => \N__33665\,
            I => \N__33656\
        );

    \I__8318\ : Span4Mux_h
    port map (
            O => \N__33662\,
            I => \N__33651\
        );

    \I__8317\ : Span4Mux_v
    port map (
            O => \N__33659\,
            I => \N__33651\
        );

    \I__8316\ : Odrv4
    port map (
            O => \N__33656\,
            I => \this_vga_signals.M_this_external_address_dZ0Z22\
        );

    \I__8315\ : Odrv4
    port map (
            O => \N__33651\,
            I => \this_vga_signals.M_this_external_address_dZ0Z22\
        );

    \I__8314\ : CascadeMux
    port map (
            O => \N__33646\,
            I => \N__33643\
        );

    \I__8313\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33638\
        );

    \I__8312\ : CascadeMux
    port map (
            O => \N__33642\,
            I => \N__33634\
        );

    \I__8311\ : CascadeMux
    port map (
            O => \N__33641\,
            I => \N__33631\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__33638\,
            I => \N__33627\
        );

    \I__8309\ : InMux
    port map (
            O => \N__33637\,
            I => \N__33624\
        );

    \I__8308\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33621\
        );

    \I__8307\ : InMux
    port map (
            O => \N__33631\,
            I => \N__33618\
        );

    \I__8306\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33615\
        );

    \I__8305\ : Span4Mux_h
    port map (
            O => \N__33627\,
            I => \N__33608\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__33624\,
            I => \N__33608\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__33621\,
            I => \N__33605\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__33618\,
            I => \N__33602\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__33615\,
            I => \N__33599\
        );

    \I__8300\ : InMux
    port map (
            O => \N__33614\,
            I => \N__33596\
        );

    \I__8299\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33592\
        );

    \I__8298\ : Span4Mux_h
    port map (
            O => \N__33608\,
            I => \N__33589\
        );

    \I__8297\ : Span4Mux_v
    port map (
            O => \N__33605\,
            I => \N__33582\
        );

    \I__8296\ : Span4Mux_v
    port map (
            O => \N__33602\,
            I => \N__33582\
        );

    \I__8295\ : Span4Mux_v
    port map (
            O => \N__33599\,
            I => \N__33582\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__33596\,
            I => \N__33579\
        );

    \I__8293\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33575\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__33592\,
            I => \N__33572\
        );

    \I__8291\ : Span4Mux_v
    port map (
            O => \N__33589\,
            I => \N__33565\
        );

    \I__8290\ : Span4Mux_h
    port map (
            O => \N__33582\,
            I => \N__33565\
        );

    \I__8289\ : Span4Mux_v
    port map (
            O => \N__33579\,
            I => \N__33565\
        );

    \I__8288\ : InMux
    port map (
            O => \N__33578\,
            I => \N__33562\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__33575\,
            I => \N__33559\
        );

    \I__8286\ : Span12Mux_h
    port map (
            O => \N__33572\,
            I => \N__33556\
        );

    \I__8285\ : Sp12to4
    port map (
            O => \N__33565\,
            I => \N__33551\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__33562\,
            I => \N__33551\
        );

    \I__8283\ : Span12Mux_v
    port map (
            O => \N__33559\,
            I => \N__33548\
        );

    \I__8282\ : Span12Mux_v
    port map (
            O => \N__33556\,
            I => \N__33543\
        );

    \I__8281\ : Span12Mux_h
    port map (
            O => \N__33551\,
            I => \N__33543\
        );

    \I__8280\ : Odrv12
    port map (
            O => \N__33548\,
            I => port_data_c_5
        );

    \I__8279\ : Odrv12
    port map (
            O => \N__33543\,
            I => port_data_c_5
        );

    \I__8278\ : CascadeMux
    port map (
            O => \N__33538\,
            I => \N__33533\
        );

    \I__8277\ : InMux
    port map (
            O => \N__33537\,
            I => \N__33529\
        );

    \I__8276\ : CascadeMux
    port map (
            O => \N__33536\,
            I => \N__33526\
        );

    \I__8275\ : InMux
    port map (
            O => \N__33533\,
            I => \N__33523\
        );

    \I__8274\ : CascadeMux
    port map (
            O => \N__33532\,
            I => \N__33520\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__33529\,
            I => \N__33516\
        );

    \I__8272\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33513\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33509\
        );

    \I__8270\ : InMux
    port map (
            O => \N__33520\,
            I => \N__33505\
        );

    \I__8269\ : InMux
    port map (
            O => \N__33519\,
            I => \N__33502\
        );

    \I__8268\ : Span4Mux_v
    port map (
            O => \N__33516\,
            I => \N__33497\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__33513\,
            I => \N__33497\
        );

    \I__8266\ : InMux
    port map (
            O => \N__33512\,
            I => \N__33493\
        );

    \I__8265\ : Span4Mux_v
    port map (
            O => \N__33509\,
            I => \N__33490\
        );

    \I__8264\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33487\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__33505\,
            I => \N__33484\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__33502\,
            I => \N__33481\
        );

    \I__8261\ : Span4Mux_v
    port map (
            O => \N__33497\,
            I => \N__33477\
        );

    \I__8260\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33474\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__33493\,
            I => \N__33471\
        );

    \I__8258\ : Span4Mux_v
    port map (
            O => \N__33490\,
            I => \N__33468\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__33487\,
            I => \N__33465\
        );

    \I__8256\ : Span4Mux_h
    port map (
            O => \N__33484\,
            I => \N__33460\
        );

    \I__8255\ : Span4Mux_h
    port map (
            O => \N__33481\,
            I => \N__33460\
        );

    \I__8254\ : InMux
    port map (
            O => \N__33480\,
            I => \N__33457\
        );

    \I__8253\ : Span4Mux_h
    port map (
            O => \N__33477\,
            I => \N__33452\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__33474\,
            I => \N__33452\
        );

    \I__8251\ : Span12Mux_v
    port map (
            O => \N__33471\,
            I => \N__33447\
        );

    \I__8250\ : Sp12to4
    port map (
            O => \N__33468\,
            I => \N__33447\
        );

    \I__8249\ : Span12Mux_s9_v
    port map (
            O => \N__33465\,
            I => \N__33438\
        );

    \I__8248\ : Sp12to4
    port map (
            O => \N__33460\,
            I => \N__33438\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__33457\,
            I => \N__33438\
        );

    \I__8246\ : Sp12to4
    port map (
            O => \N__33452\,
            I => \N__33438\
        );

    \I__8245\ : Span12Mux_h
    port map (
            O => \N__33447\,
            I => \N__33435\
        );

    \I__8244\ : Span12Mux_v
    port map (
            O => \N__33438\,
            I => \N__33432\
        );

    \I__8243\ : Odrv12
    port map (
            O => \N__33435\,
            I => port_data_c_6
        );

    \I__8242\ : Odrv12
    port map (
            O => \N__33432\,
            I => port_data_c_6
        );

    \I__8241\ : CascadeMux
    port map (
            O => \N__33427\,
            I => \N__33423\
        );

    \I__8240\ : CascadeMux
    port map (
            O => \N__33426\,
            I => \N__33418\
        );

    \I__8239\ : InMux
    port map (
            O => \N__33423\,
            I => \N__33415\
        );

    \I__8238\ : InMux
    port map (
            O => \N__33422\,
            I => \N__33412\
        );

    \I__8237\ : InMux
    port map (
            O => \N__33421\,
            I => \N__33407\
        );

    \I__8236\ : InMux
    port map (
            O => \N__33418\,
            I => \N__33407\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__33415\,
            I => \N__33403\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__33412\,
            I => \N__33400\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__33407\,
            I => \N__33397\
        );

    \I__8232\ : InMux
    port map (
            O => \N__33406\,
            I => \N__33394\
        );

    \I__8231\ : Span4Mux_v
    port map (
            O => \N__33403\,
            I => \N__33391\
        );

    \I__8230\ : Span4Mux_v
    port map (
            O => \N__33400\,
            I => \N__33382\
        );

    \I__8229\ : Span4Mux_h
    port map (
            O => \N__33397\,
            I => \N__33382\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__33394\,
            I => \N__33382\
        );

    \I__8227\ : Span4Mux_h
    port map (
            O => \N__33391\,
            I => \N__33379\
        );

    \I__8226\ : InMux
    port map (
            O => \N__33390\,
            I => \N__33376\
        );

    \I__8225\ : CascadeMux
    port map (
            O => \N__33389\,
            I => \N__33373\
        );

    \I__8224\ : Span4Mux_v
    port map (
            O => \N__33382\,
            I => \N__33370\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__33379\,
            I => \N__33365\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__33376\,
            I => \N__33365\
        );

    \I__8221\ : InMux
    port map (
            O => \N__33373\,
            I => \N__33362\
        );

    \I__8220\ : Span4Mux_v
    port map (
            O => \N__33370\,
            I => \N__33357\
        );

    \I__8219\ : Span4Mux_v
    port map (
            O => \N__33365\,
            I => \N__33357\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__33362\,
            I => \N__33354\
        );

    \I__8217\ : Span4Mux_h
    port map (
            O => \N__33357\,
            I => \N__33351\
        );

    \I__8216\ : Span12Mux_v
    port map (
            O => \N__33354\,
            I => \N__33348\
        );

    \I__8215\ : IoSpan4Mux
    port map (
            O => \N__33351\,
            I => \N__33345\
        );

    \I__8214\ : Odrv12
    port map (
            O => \N__33348\,
            I => port_data_c_7
        );

    \I__8213\ : Odrv4
    port map (
            O => \N__33345\,
            I => port_data_c_7
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__33340\,
            I => \N__33337\
        );

    \I__8211\ : InMux
    port map (
            O => \N__33337\,
            I => \N__33333\
        );

    \I__8210\ : CascadeMux
    port map (
            O => \N__33336\,
            I => \N__33330\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33323\
        );

    \I__8208\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33320\
        );

    \I__8207\ : CascadeMux
    port map (
            O => \N__33329\,
            I => \N__33316\
        );

    \I__8206\ : CascadeMux
    port map (
            O => \N__33328\,
            I => \N__33313\
        );

    \I__8205\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33308\
        );

    \I__8204\ : CascadeMux
    port map (
            O => \N__33326\,
            I => \N__33305\
        );

    \I__8203\ : Span4Mux_v
    port map (
            O => \N__33323\,
            I => \N__33300\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__33320\,
            I => \N__33300\
        );

    \I__8201\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33297\
        );

    \I__8200\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33294\
        );

    \I__8199\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33291\
        );

    \I__8198\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33288\
        );

    \I__8197\ : CascadeMux
    port map (
            O => \N__33311\,
            I => \N__33285\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__33308\,
            I => \N__33282\
        );

    \I__8195\ : InMux
    port map (
            O => \N__33305\,
            I => \N__33279\
        );

    \I__8194\ : Span4Mux_h
    port map (
            O => \N__33300\,
            I => \N__33270\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__33297\,
            I => \N__33270\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__33294\,
            I => \N__33270\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__33291\,
            I => \N__33270\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__33288\,
            I => \N__33267\
        );

    \I__8189\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33263\
        );

    \I__8188\ : Span4Mux_v
    port map (
            O => \N__33282\,
            I => \N__33258\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__33279\,
            I => \N__33258\
        );

    \I__8186\ : Span4Mux_v
    port map (
            O => \N__33270\,
            I => \N__33255\
        );

    \I__8185\ : Span4Mux_v
    port map (
            O => \N__33267\,
            I => \N__33252\
        );

    \I__8184\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33249\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__33263\,
            I => \N__33245\
        );

    \I__8182\ : Span4Mux_v
    port map (
            O => \N__33258\,
            I => \N__33242\
        );

    \I__8181\ : Span4Mux_h
    port map (
            O => \N__33255\,
            I => \N__33237\
        );

    \I__8180\ : Span4Mux_v
    port map (
            O => \N__33252\,
            I => \N__33237\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__33249\,
            I => \N__33234\
        );

    \I__8178\ : InMux
    port map (
            O => \N__33248\,
            I => \N__33231\
        );

    \I__8177\ : Span12Mux_v
    port map (
            O => \N__33245\,
            I => \N__33228\
        );

    \I__8176\ : Span4Mux_v
    port map (
            O => \N__33242\,
            I => \N__33225\
        );

    \I__8175\ : Span4Mux_v
    port map (
            O => \N__33237\,
            I => \N__33220\
        );

    \I__8174\ : Span4Mux_v
    port map (
            O => \N__33234\,
            I => \N__33220\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__33231\,
            I => \N__33217\
        );

    \I__8172\ : Span12Mux_h
    port map (
            O => \N__33228\,
            I => \N__33214\
        );

    \I__8171\ : Sp12to4
    port map (
            O => \N__33225\,
            I => \N__33211\
        );

    \I__8170\ : Sp12to4
    port map (
            O => \N__33220\,
            I => \N__33206\
        );

    \I__8169\ : Span12Mux_v
    port map (
            O => \N__33217\,
            I => \N__33206\
        );

    \I__8168\ : Odrv12
    port map (
            O => \N__33214\,
            I => port_data_c_4
        );

    \I__8167\ : Odrv12
    port map (
            O => \N__33211\,
            I => port_data_c_4
        );

    \I__8166\ : Odrv12
    port map (
            O => \N__33206\,
            I => port_data_c_4
        );

    \I__8165\ : InMux
    port map (
            O => \N__33199\,
            I => \N__33193\
        );

    \I__8164\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33193\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__33193\,
            I => \N__33190\
        );

    \I__8162\ : Odrv4
    port map (
            O => \N__33190\,
            I => \this_vga_signals.M_this_external_address_d21Z0Z_6\
        );

    \I__8161\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33184\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__33184\,
            I => \N__33181\
        );

    \I__8159\ : Span4Mux_v
    port map (
            O => \N__33181\,
            I => \N__33178\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__33178\,
            I => \M_this_map_ram_write_data_7\
        );

    \I__8157\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33171\
        );

    \I__8156\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33168\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__33171\,
            I => \N__33165\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__33168\,
            I => \this_ppu.M_haddress_qZ0Z_7\
        );

    \I__8153\ : Odrv12
    port map (
            O => \N__33165\,
            I => \this_ppu.M_haddress_qZ0Z_7\
        );

    \I__8152\ : CascadeMux
    port map (
            O => \N__33160\,
            I => \N__33157\
        );

    \I__8151\ : CascadeBuf
    port map (
            O => \N__33157\,
            I => \N__33154\
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__33154\,
            I => \N__33151\
        );

    \I__8149\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33148\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__33148\,
            I => \N__33145\
        );

    \I__8147\ : Span4Mux_v
    port map (
            O => \N__33145\,
            I => \N__33142\
        );

    \I__8146\ : Odrv4
    port map (
            O => \N__33142\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__8145\ : CascadeMux
    port map (
            O => \N__33139\,
            I => \N__33136\
        );

    \I__8144\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33133\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__33133\,
            I => \N__33130\
        );

    \I__8142\ : Span4Mux_h
    port map (
            O => \N__33130\,
            I => \N__33127\
        );

    \I__8141\ : Span4Mux_v
    port map (
            O => \N__33127\,
            I => \N__33122\
        );

    \I__8140\ : InMux
    port map (
            O => \N__33126\,
            I => \N__33117\
        );

    \I__8139\ : InMux
    port map (
            O => \N__33125\,
            I => \N__33117\
        );

    \I__8138\ : Span4Mux_v
    port map (
            O => \N__33122\,
            I => \N__33110\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33110\
        );

    \I__8136\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33107\
        );

    \I__8135\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33104\
        );

    \I__8134\ : Span4Mux_h
    port map (
            O => \N__33110\,
            I => \N__33101\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__33107\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__33104\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__8131\ : Odrv4
    port map (
            O => \N__33101\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__8130\ : CascadeMux
    port map (
            O => \N__33094\,
            I => \N__33091\
        );

    \I__8129\ : CascadeBuf
    port map (
            O => \N__33091\,
            I => \N__33088\
        );

    \I__8128\ : CascadeMux
    port map (
            O => \N__33088\,
            I => \N__33085\
        );

    \I__8127\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33082\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__33082\,
            I => \N__33079\
        );

    \I__8125\ : Span4Mux_s3_v
    port map (
            O => \N__33079\,
            I => \N__33076\
        );

    \I__8124\ : Odrv4
    port map (
            O => \N__33076\,
            I => \M_this_ppu_vram_addr_i_6\
        );

    \I__8123\ : InMux
    port map (
            O => \N__33073\,
            I => \N__33070\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__33070\,
            I => \M_this_map_ram_write_data_2\
        );

    \I__8121\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33064\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__33064\,
            I => \N__33061\
        );

    \I__8119\ : Odrv4
    port map (
            O => \N__33061\,
            I => \M_this_map_ram_write_data_1\
        );

    \I__8118\ : InMux
    port map (
            O => \N__33058\,
            I => \N__33055\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__33055\,
            I => \M_this_map_ram_write_data_0\
        );

    \I__8116\ : InMux
    port map (
            O => \N__33052\,
            I => \N__33049\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__33049\,
            I => \M_this_map_ram_write_data_5\
        );

    \I__8114\ : CascadeMux
    port map (
            O => \N__33046\,
            I => \N__33040\
        );

    \I__8113\ : CEMux
    port map (
            O => \N__33045\,
            I => \N__33036\
        );

    \I__8112\ : CEMux
    port map (
            O => \N__33044\,
            I => \N__33033\
        );

    \I__8111\ : InMux
    port map (
            O => \N__33043\,
            I => \N__33030\
        );

    \I__8110\ : InMux
    port map (
            O => \N__33040\,
            I => \N__33025\
        );

    \I__8109\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33025\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__33036\,
            I => \N__33019\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__33033\,
            I => \N__33012\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__33030\,
            I => \N__33012\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__33025\,
            I => \N__33012\
        );

    \I__8104\ : InMux
    port map (
            O => \N__33024\,
            I => \N__33007\
        );

    \I__8103\ : InMux
    port map (
            O => \N__33023\,
            I => \N__33007\
        );

    \I__8102\ : InMux
    port map (
            O => \N__33022\,
            I => \N__33002\
        );

    \I__8101\ : Span4Mux_v
    port map (
            O => \N__33019\,
            I => \N__32994\
        );

    \I__8100\ : Span4Mux_v
    port map (
            O => \N__33012\,
            I => \N__32994\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__33007\,
            I => \N__32994\
        );

    \I__8098\ : InMux
    port map (
            O => \N__33006\,
            I => \N__32989\
        );

    \I__8097\ : InMux
    port map (
            O => \N__33005\,
            I => \N__32989\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__33002\,
            I => \N__32986\
        );

    \I__8095\ : InMux
    port map (
            O => \N__33001\,
            I => \N__32981\
        );

    \I__8094\ : Span4Mux_h
    port map (
            O => \N__32994\,
            I => \N__32978\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__32989\,
            I => \N__32975\
        );

    \I__8092\ : Span12Mux_h
    port map (
            O => \N__32986\,
            I => \N__32972\
        );

    \I__8091\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32967\
        );

    \I__8090\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32967\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__32981\,
            I => \N__32960\
        );

    \I__8088\ : Span4Mux_v
    port map (
            O => \N__32978\,
            I => \N__32960\
        );

    \I__8087\ : Span4Mux_h
    port map (
            O => \N__32975\,
            I => \N__32960\
        );

    \I__8086\ : Span12Mux_v
    port map (
            O => \N__32972\,
            I => \N__32957\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__32967\,
            I => \N__32952\
        );

    \I__8084\ : Span4Mux_v
    port map (
            O => \N__32960\,
            I => \N__32952\
        );

    \I__8083\ : Odrv12
    port map (
            O => \N__32957\,
            I => \M_this_map_ram_write_en_0\
        );

    \I__8082\ : Odrv4
    port map (
            O => \N__32952\,
            I => \M_this_map_ram_write_en_0\
        );

    \I__8081\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32944\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__32944\,
            I => \M_this_map_ram_write_data_4\
        );

    \I__8079\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32938\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__32938\,
            I => \M_this_data_count_q_cry_9_THRU_CO\
        );

    \I__8077\ : CascadeMux
    port map (
            O => \N__32935\,
            I => \M_this_data_count_q_3_10_cascade_\
        );

    \I__8076\ : CascadeMux
    port map (
            O => \N__32932\,
            I => \N__32926\
        );

    \I__8075\ : InMux
    port map (
            O => \N__32931\,
            I => \N__32920\
        );

    \I__8074\ : InMux
    port map (
            O => \N__32930\,
            I => \N__32917\
        );

    \I__8073\ : InMux
    port map (
            O => \N__32929\,
            I => \N__32913\
        );

    \I__8072\ : InMux
    port map (
            O => \N__32926\,
            I => \N__32910\
        );

    \I__8071\ : InMux
    port map (
            O => \N__32925\,
            I => \N__32907\
        );

    \I__8070\ : InMux
    port map (
            O => \N__32924\,
            I => \N__32904\
        );

    \I__8069\ : InMux
    port map (
            O => \N__32923\,
            I => \N__32901\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__32920\,
            I => \N__32898\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__32917\,
            I => \N__32895\
        );

    \I__8066\ : InMux
    port map (
            O => \N__32916\,
            I => \N__32892\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__32913\,
            I => \N__32889\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__32910\,
            I => \N__32886\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__32907\,
            I => \N__32883\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__32904\,
            I => \N__32880\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__32901\,
            I => \N__32877\
        );

    \I__8060\ : Span4Mux_h
    port map (
            O => \N__32898\,
            I => \N__32872\
        );

    \I__8059\ : Span4Mux_h
    port map (
            O => \N__32895\,
            I => \N__32872\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__32892\,
            I => \N__32861\
        );

    \I__8057\ : Span4Mux_v
    port map (
            O => \N__32889\,
            I => \N__32861\
        );

    \I__8056\ : Span4Mux_v
    port map (
            O => \N__32886\,
            I => \N__32861\
        );

    \I__8055\ : Span4Mux_v
    port map (
            O => \N__32883\,
            I => \N__32861\
        );

    \I__8054\ : Span4Mux_h
    port map (
            O => \N__32880\,
            I => \N__32861\
        );

    \I__8053\ : Odrv12
    port map (
            O => \N__32877\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__8052\ : Odrv4
    port map (
            O => \N__32872\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__8051\ : Odrv4
    port map (
            O => \N__32861\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__8050\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32840\
        );

    \I__8049\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32835\
        );

    \I__8048\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32835\
        );

    \I__8047\ : CascadeMux
    port map (
            O => \N__32851\,
            I => \N__32831\
        );

    \I__8046\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32818\
        );

    \I__8045\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32815\
        );

    \I__8044\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32812\
        );

    \I__8043\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32805\
        );

    \I__8042\ : InMux
    port map (
            O => \N__32846\,
            I => \N__32805\
        );

    \I__8041\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32805\
        );

    \I__8040\ : InMux
    port map (
            O => \N__32844\,
            I => \N__32800\
        );

    \I__8039\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32800\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__32840\,
            I => \N__32795\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__32835\,
            I => \N__32795\
        );

    \I__8036\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32792\
        );

    \I__8035\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32781\
        );

    \I__8034\ : InMux
    port map (
            O => \N__32830\,
            I => \N__32778\
        );

    \I__8033\ : InMux
    port map (
            O => \N__32829\,
            I => \N__32765\
        );

    \I__8032\ : InMux
    port map (
            O => \N__32828\,
            I => \N__32765\
        );

    \I__8031\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32762\
        );

    \I__8030\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32747\
        );

    \I__8029\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32743\
        );

    \I__8028\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32740\
        );

    \I__8027\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32735\
        );

    \I__8026\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32735\
        );

    \I__8025\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32732\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__32818\,
            I => \N__32727\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__32815\,
            I => \N__32727\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__32812\,
            I => \N__32724\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__32805\,
            I => \N__32716\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__32800\,
            I => \N__32716\
        );

    \I__8019\ : Span4Mux_h
    port map (
            O => \N__32795\,
            I => \N__32716\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__32792\,
            I => \N__32713\
        );

    \I__8017\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32710\
        );

    \I__8016\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32707\
        );

    \I__8015\ : InMux
    port map (
            O => \N__32789\,
            I => \N__32704\
        );

    \I__8014\ : InMux
    port map (
            O => \N__32788\,
            I => \N__32699\
        );

    \I__8013\ : InMux
    port map (
            O => \N__32787\,
            I => \N__32699\
        );

    \I__8012\ : InMux
    port map (
            O => \N__32786\,
            I => \N__32696\
        );

    \I__8011\ : InMux
    port map (
            O => \N__32785\,
            I => \N__32691\
        );

    \I__8010\ : InMux
    port map (
            O => \N__32784\,
            I => \N__32691\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__32781\,
            I => \N__32688\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__32778\,
            I => \N__32685\
        );

    \I__8007\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32682\
        );

    \I__8006\ : InMux
    port map (
            O => \N__32776\,
            I => \N__32675\
        );

    \I__8005\ : InMux
    port map (
            O => \N__32775\,
            I => \N__32675\
        );

    \I__8004\ : InMux
    port map (
            O => \N__32774\,
            I => \N__32675\
        );

    \I__8003\ : InMux
    port map (
            O => \N__32773\,
            I => \N__32672\
        );

    \I__8002\ : InMux
    port map (
            O => \N__32772\,
            I => \N__32669\
        );

    \I__8001\ : InMux
    port map (
            O => \N__32771\,
            I => \N__32664\
        );

    \I__8000\ : InMux
    port map (
            O => \N__32770\,
            I => \N__32664\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__32765\,
            I => \N__32659\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__32762\,
            I => \N__32659\
        );

    \I__7997\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32650\
        );

    \I__7996\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32650\
        );

    \I__7995\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32650\
        );

    \I__7994\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32650\
        );

    \I__7993\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32645\
        );

    \I__7992\ : InMux
    port map (
            O => \N__32756\,
            I => \N__32645\
        );

    \I__7991\ : InMux
    port map (
            O => \N__32755\,
            I => \N__32640\
        );

    \I__7990\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32640\
        );

    \I__7989\ : InMux
    port map (
            O => \N__32753\,
            I => \N__32634\
        );

    \I__7988\ : InMux
    port map (
            O => \N__32752\,
            I => \N__32629\
        );

    \I__7987\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32629\
        );

    \I__7986\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32626\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__32747\,
            I => \N__32617\
        );

    \I__7984\ : InMux
    port map (
            O => \N__32746\,
            I => \N__32613\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__32743\,
            I => \N__32600\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__32740\,
            I => \N__32600\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__32735\,
            I => \N__32600\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__32732\,
            I => \N__32600\
        );

    \I__7979\ : Sp12to4
    port map (
            O => \N__32727\,
            I => \N__32600\
        );

    \I__7978\ : Sp12to4
    port map (
            O => \N__32724\,
            I => \N__32600\
        );

    \I__7977\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32597\
        );

    \I__7976\ : Span4Mux_v
    port map (
            O => \N__32716\,
            I => \N__32590\
        );

    \I__7975\ : Span4Mux_h
    port map (
            O => \N__32713\,
            I => \N__32590\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__32710\,
            I => \N__32590\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__32707\,
            I => \N__32585\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__32704\,
            I => \N__32582\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__32699\,
            I => \N__32577\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__32696\,
            I => \N__32577\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__32691\,
            I => \N__32574\
        );

    \I__7968\ : Span4Mux_v
    port map (
            O => \N__32688\,
            I => \N__32567\
        );

    \I__7967\ : Span4Mux_v
    port map (
            O => \N__32685\,
            I => \N__32567\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__32682\,
            I => \N__32567\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__32675\,
            I => \N__32564\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__32672\,
            I => \N__32561\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__32669\,
            I => \N__32548\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__32664\,
            I => \N__32548\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__32659\,
            I => \N__32548\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__32650\,
            I => \N__32548\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__32645\,
            I => \N__32548\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__32640\,
            I => \N__32548\
        );

    \I__7957\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32545\
        );

    \I__7956\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32542\
        );

    \I__7955\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32539\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__32634\,
            I => \N__32532\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__32629\,
            I => \N__32532\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32532\
        );

    \I__7951\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32529\
        );

    \I__7950\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32526\
        );

    \I__7949\ : InMux
    port map (
            O => \N__32623\,
            I => \N__32523\
        );

    \I__7948\ : InMux
    port map (
            O => \N__32622\,
            I => \N__32518\
        );

    \I__7947\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32518\
        );

    \I__7946\ : InMux
    port map (
            O => \N__32620\,
            I => \N__32515\
        );

    \I__7945\ : Span12Mux_h
    port map (
            O => \N__32617\,
            I => \N__32512\
        );

    \I__7944\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32509\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32502\
        );

    \I__7942\ : Span12Mux_v
    port map (
            O => \N__32600\,
            I => \N__32502\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__32597\,
            I => \N__32502\
        );

    \I__7940\ : Span4Mux_v
    port map (
            O => \N__32590\,
            I => \N__32499\
        );

    \I__7939\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32494\
        );

    \I__7938\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32494\
        );

    \I__7937\ : Span4Mux_h
    port map (
            O => \N__32585\,
            I => \N__32487\
        );

    \I__7936\ : Span4Mux_h
    port map (
            O => \N__32582\,
            I => \N__32487\
        );

    \I__7935\ : Span4Mux_h
    port map (
            O => \N__32577\,
            I => \N__32487\
        );

    \I__7934\ : Span4Mux_h
    port map (
            O => \N__32574\,
            I => \N__32476\
        );

    \I__7933\ : Span4Mux_h
    port map (
            O => \N__32567\,
            I => \N__32476\
        );

    \I__7932\ : Span4Mux_h
    port map (
            O => \N__32564\,
            I => \N__32476\
        );

    \I__7931\ : Span4Mux_h
    port map (
            O => \N__32561\,
            I => \N__32476\
        );

    \I__7930\ : Span4Mux_v
    port map (
            O => \N__32548\,
            I => \N__32476\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__32545\,
            I => \N__32471\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__32542\,
            I => \N__32471\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__32539\,
            I => \N__32464\
        );

    \I__7926\ : Span4Mux_v
    port map (
            O => \N__32532\,
            I => \N__32464\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__32529\,
            I => \N__32464\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__32526\,
            I => \N_389_0\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__32523\,
            I => \N_389_0\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__32518\,
            I => \N_389_0\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__32515\,
            I => \N_389_0\
        );

    \I__7920\ : Odrv12
    port map (
            O => \N__32512\,
            I => \N_389_0\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__32509\,
            I => \N_389_0\
        );

    \I__7918\ : Odrv12
    port map (
            O => \N__32502\,
            I => \N_389_0\
        );

    \I__7917\ : Odrv4
    port map (
            O => \N__32499\,
            I => \N_389_0\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__32494\,
            I => \N_389_0\
        );

    \I__7915\ : Odrv4
    port map (
            O => \N__32487\,
            I => \N_389_0\
        );

    \I__7914\ : Odrv4
    port map (
            O => \N__32476\,
            I => \N_389_0\
        );

    \I__7913\ : Odrv12
    port map (
            O => \N__32471\,
            I => \N_389_0\
        );

    \I__7912\ : Odrv4
    port map (
            O => \N__32464\,
            I => \N_389_0\
        );

    \I__7911\ : InMux
    port map (
            O => \N__32437\,
            I => \N__32424\
        );

    \I__7910\ : InMux
    port map (
            O => \N__32436\,
            I => \N__32421\
        );

    \I__7909\ : InMux
    port map (
            O => \N__32435\,
            I => \N__32418\
        );

    \I__7908\ : InMux
    port map (
            O => \N__32434\,
            I => \N__32415\
        );

    \I__7907\ : InMux
    port map (
            O => \N__32433\,
            I => \N__32412\
        );

    \I__7906\ : InMux
    port map (
            O => \N__32432\,
            I => \N__32409\
        );

    \I__7905\ : InMux
    port map (
            O => \N__32431\,
            I => \N__32406\
        );

    \I__7904\ : InMux
    port map (
            O => \N__32430\,
            I => \N__32403\
        );

    \I__7903\ : InMux
    port map (
            O => \N__32429\,
            I => \N__32400\
        );

    \I__7902\ : InMux
    port map (
            O => \N__32428\,
            I => \N__32397\
        );

    \I__7901\ : InMux
    port map (
            O => \N__32427\,
            I => \N__32394\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__32424\,
            I => \N__32370\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__32421\,
            I => \N__32367\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32364\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__32415\,
            I => \N__32361\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__32412\,
            I => \N__32358\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__32409\,
            I => \N__32355\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__32406\,
            I => \N__32352\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__32403\,
            I => \N__32349\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__32400\,
            I => \N__32346\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__32397\,
            I => \N__32343\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__32394\,
            I => \N__32340\
        );

    \I__7889\ : SRMux
    port map (
            O => \N__32393\,
            I => \N__32275\
        );

    \I__7888\ : SRMux
    port map (
            O => \N__32392\,
            I => \N__32275\
        );

    \I__7887\ : SRMux
    port map (
            O => \N__32391\,
            I => \N__32275\
        );

    \I__7886\ : SRMux
    port map (
            O => \N__32390\,
            I => \N__32275\
        );

    \I__7885\ : SRMux
    port map (
            O => \N__32389\,
            I => \N__32275\
        );

    \I__7884\ : SRMux
    port map (
            O => \N__32388\,
            I => \N__32275\
        );

    \I__7883\ : SRMux
    port map (
            O => \N__32387\,
            I => \N__32275\
        );

    \I__7882\ : SRMux
    port map (
            O => \N__32386\,
            I => \N__32275\
        );

    \I__7881\ : SRMux
    port map (
            O => \N__32385\,
            I => \N__32275\
        );

    \I__7880\ : SRMux
    port map (
            O => \N__32384\,
            I => \N__32275\
        );

    \I__7879\ : SRMux
    port map (
            O => \N__32383\,
            I => \N__32275\
        );

    \I__7878\ : SRMux
    port map (
            O => \N__32382\,
            I => \N__32275\
        );

    \I__7877\ : SRMux
    port map (
            O => \N__32381\,
            I => \N__32275\
        );

    \I__7876\ : SRMux
    port map (
            O => \N__32380\,
            I => \N__32275\
        );

    \I__7875\ : SRMux
    port map (
            O => \N__32379\,
            I => \N__32275\
        );

    \I__7874\ : SRMux
    port map (
            O => \N__32378\,
            I => \N__32275\
        );

    \I__7873\ : SRMux
    port map (
            O => \N__32377\,
            I => \N__32275\
        );

    \I__7872\ : SRMux
    port map (
            O => \N__32376\,
            I => \N__32275\
        );

    \I__7871\ : SRMux
    port map (
            O => \N__32375\,
            I => \N__32275\
        );

    \I__7870\ : SRMux
    port map (
            O => \N__32374\,
            I => \N__32275\
        );

    \I__7869\ : SRMux
    port map (
            O => \N__32373\,
            I => \N__32275\
        );

    \I__7868\ : Glb2LocalMux
    port map (
            O => \N__32370\,
            I => \N__32275\
        );

    \I__7867\ : Glb2LocalMux
    port map (
            O => \N__32367\,
            I => \N__32275\
        );

    \I__7866\ : Glb2LocalMux
    port map (
            O => \N__32364\,
            I => \N__32275\
        );

    \I__7865\ : Glb2LocalMux
    port map (
            O => \N__32361\,
            I => \N__32275\
        );

    \I__7864\ : Glb2LocalMux
    port map (
            O => \N__32358\,
            I => \N__32275\
        );

    \I__7863\ : Glb2LocalMux
    port map (
            O => \N__32355\,
            I => \N__32275\
        );

    \I__7862\ : Glb2LocalMux
    port map (
            O => \N__32352\,
            I => \N__32275\
        );

    \I__7861\ : Glb2LocalMux
    port map (
            O => \N__32349\,
            I => \N__32275\
        );

    \I__7860\ : Glb2LocalMux
    port map (
            O => \N__32346\,
            I => \N__32275\
        );

    \I__7859\ : Glb2LocalMux
    port map (
            O => \N__32343\,
            I => \N__32275\
        );

    \I__7858\ : Glb2LocalMux
    port map (
            O => \N__32340\,
            I => \N__32275\
        );

    \I__7857\ : GlobalMux
    port map (
            O => \N__32275\,
            I => \N__32272\
        );

    \I__7856\ : gio2CtrlBuf
    port map (
            O => \N__32272\,
            I => \M_this_reset_cond_out_g_0\
        );

    \I__7855\ : CascadeMux
    port map (
            O => \N__32269\,
            I => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8_cascade_\
        );

    \I__7854\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32263\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__32263\,
            I => \N__32260\
        );

    \I__7852\ : Odrv4
    port map (
            O => \N__32260\,
            I => \this_vga_signals.M_this_data_count_q_3_bmZ0Z_13\
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__32257\,
            I => \this_vga_signals.M_this_data_count_q_3_amZ0Z_13_cascade_\
        );

    \I__7850\ : InMux
    port map (
            O => \N__32254\,
            I => \N__32242\
        );

    \I__7849\ : InMux
    port map (
            O => \N__32253\,
            I => \N__32242\
        );

    \I__7848\ : InMux
    port map (
            O => \N__32252\,
            I => \N__32242\
        );

    \I__7847\ : InMux
    port map (
            O => \N__32251\,
            I => \N__32227\
        );

    \I__7846\ : InMux
    port map (
            O => \N__32250\,
            I => \N__32227\
        );

    \I__7845\ : InMux
    port map (
            O => \N__32249\,
            I => \N__32227\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32224\
        );

    \I__7843\ : InMux
    port map (
            O => \N__32241\,
            I => \N__32219\
        );

    \I__7842\ : InMux
    port map (
            O => \N__32240\,
            I => \N__32219\
        );

    \I__7841\ : InMux
    port map (
            O => \N__32239\,
            I => \N__32214\
        );

    \I__7840\ : InMux
    port map (
            O => \N__32238\,
            I => \N__32214\
        );

    \I__7839\ : InMux
    port map (
            O => \N__32237\,
            I => \N__32205\
        );

    \I__7838\ : InMux
    port map (
            O => \N__32236\,
            I => \N__32205\
        );

    \I__7837\ : InMux
    port map (
            O => \N__32235\,
            I => \N__32205\
        );

    \I__7836\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32205\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__32227\,
            I => \N__32200\
        );

    \I__7834\ : Sp12to4
    port map (
            O => \N__32224\,
            I => \N__32193\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__32219\,
            I => \N__32193\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__32214\,
            I => \N__32193\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32190\
        );

    \I__7830\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32185\
        );

    \I__7829\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32185\
        );

    \I__7828\ : Odrv4
    port map (
            O => \N__32200\,
            I => \M_this_data_count_q_3_sn_N_2\
        );

    \I__7827\ : Odrv12
    port map (
            O => \N__32193\,
            I => \M_this_data_count_q_3_sn_N_2\
        );

    \I__7826\ : Odrv4
    port map (
            O => \N__32190\,
            I => \M_this_data_count_q_3_sn_N_2\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__32185\,
            I => \M_this_data_count_q_3_sn_N_2\
        );

    \I__7824\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32173\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__32173\,
            I => \M_this_data_count_q_cry_12_THRU_CO\
        );

    \I__7822\ : CascadeMux
    port map (
            O => \N__32170\,
            I => \M_this_data_count_q_3_13_cascade_\
        );

    \I__7821\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32147\
        );

    \I__7820\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32147\
        );

    \I__7819\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32147\
        );

    \I__7818\ : InMux
    port map (
            O => \N__32164\,
            I => \N__32138\
        );

    \I__7817\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32138\
        );

    \I__7816\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32138\
        );

    \I__7815\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32138\
        );

    \I__7814\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32127\
        );

    \I__7813\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32127\
        );

    \I__7812\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32127\
        );

    \I__7811\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32127\
        );

    \I__7810\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32120\
        );

    \I__7809\ : InMux
    port map (
            O => \N__32155\,
            I => \N__32120\
        );

    \I__7808\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32120\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__32147\,
            I => \N__32115\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__32138\,
            I => \N__32115\
        );

    \I__7805\ : InMux
    port map (
            O => \N__32137\,
            I => \N__32110\
        );

    \I__7804\ : InMux
    port map (
            O => \N__32136\,
            I => \N__32110\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__32127\,
            I => \N__32107\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__32120\,
            I => \N__32104\
        );

    \I__7801\ : Span4Mux_v
    port map (
            O => \N__32115\,
            I => \N__32099\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__32110\,
            I => \N__32099\
        );

    \I__7799\ : Odrv4
    port map (
            O => \N__32107\,
            I => \N_570_0_i\
        );

    \I__7798\ : Odrv4
    port map (
            O => \N__32104\,
            I => \N_570_0_i\
        );

    \I__7797\ : Odrv4
    port map (
            O => \N__32099\,
            I => \N_570_0_i\
        );

    \I__7796\ : InMux
    port map (
            O => \N__32092\,
            I => \N__32089\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__32089\,
            I => \N__32083\
        );

    \I__7794\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32080\
        );

    \I__7793\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32077\
        );

    \I__7792\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32074\
        );

    \I__7791\ : Span4Mux_h
    port map (
            O => \N__32083\,
            I => \N__32071\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__32080\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__32077\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__32074\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__7787\ : Odrv4
    port map (
            O => \N__32071\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__7786\ : ClkMux
    port map (
            O => \N__32062\,
            I => \N__31684\
        );

    \I__7785\ : ClkMux
    port map (
            O => \N__32061\,
            I => \N__31684\
        );

    \I__7784\ : ClkMux
    port map (
            O => \N__32060\,
            I => \N__31684\
        );

    \I__7783\ : ClkMux
    port map (
            O => \N__32059\,
            I => \N__31684\
        );

    \I__7782\ : ClkMux
    port map (
            O => \N__32058\,
            I => \N__31684\
        );

    \I__7781\ : ClkMux
    port map (
            O => \N__32057\,
            I => \N__31684\
        );

    \I__7780\ : ClkMux
    port map (
            O => \N__32056\,
            I => \N__31684\
        );

    \I__7779\ : ClkMux
    port map (
            O => \N__32055\,
            I => \N__31684\
        );

    \I__7778\ : ClkMux
    port map (
            O => \N__32054\,
            I => \N__31684\
        );

    \I__7777\ : ClkMux
    port map (
            O => \N__32053\,
            I => \N__31684\
        );

    \I__7776\ : ClkMux
    port map (
            O => \N__32052\,
            I => \N__31684\
        );

    \I__7775\ : ClkMux
    port map (
            O => \N__32051\,
            I => \N__31684\
        );

    \I__7774\ : ClkMux
    port map (
            O => \N__32050\,
            I => \N__31684\
        );

    \I__7773\ : ClkMux
    port map (
            O => \N__32049\,
            I => \N__31684\
        );

    \I__7772\ : ClkMux
    port map (
            O => \N__32048\,
            I => \N__31684\
        );

    \I__7771\ : ClkMux
    port map (
            O => \N__32047\,
            I => \N__31684\
        );

    \I__7770\ : ClkMux
    port map (
            O => \N__32046\,
            I => \N__31684\
        );

    \I__7769\ : ClkMux
    port map (
            O => \N__32045\,
            I => \N__31684\
        );

    \I__7768\ : ClkMux
    port map (
            O => \N__32044\,
            I => \N__31684\
        );

    \I__7767\ : ClkMux
    port map (
            O => \N__32043\,
            I => \N__31684\
        );

    \I__7766\ : ClkMux
    port map (
            O => \N__32042\,
            I => \N__31684\
        );

    \I__7765\ : ClkMux
    port map (
            O => \N__32041\,
            I => \N__31684\
        );

    \I__7764\ : ClkMux
    port map (
            O => \N__32040\,
            I => \N__31684\
        );

    \I__7763\ : ClkMux
    port map (
            O => \N__32039\,
            I => \N__31684\
        );

    \I__7762\ : ClkMux
    port map (
            O => \N__32038\,
            I => \N__31684\
        );

    \I__7761\ : ClkMux
    port map (
            O => \N__32037\,
            I => \N__31684\
        );

    \I__7760\ : ClkMux
    port map (
            O => \N__32036\,
            I => \N__31684\
        );

    \I__7759\ : ClkMux
    port map (
            O => \N__32035\,
            I => \N__31684\
        );

    \I__7758\ : ClkMux
    port map (
            O => \N__32034\,
            I => \N__31684\
        );

    \I__7757\ : ClkMux
    port map (
            O => \N__32033\,
            I => \N__31684\
        );

    \I__7756\ : ClkMux
    port map (
            O => \N__32032\,
            I => \N__31684\
        );

    \I__7755\ : ClkMux
    port map (
            O => \N__32031\,
            I => \N__31684\
        );

    \I__7754\ : ClkMux
    port map (
            O => \N__32030\,
            I => \N__31684\
        );

    \I__7753\ : ClkMux
    port map (
            O => \N__32029\,
            I => \N__31684\
        );

    \I__7752\ : ClkMux
    port map (
            O => \N__32028\,
            I => \N__31684\
        );

    \I__7751\ : ClkMux
    port map (
            O => \N__32027\,
            I => \N__31684\
        );

    \I__7750\ : ClkMux
    port map (
            O => \N__32026\,
            I => \N__31684\
        );

    \I__7749\ : ClkMux
    port map (
            O => \N__32025\,
            I => \N__31684\
        );

    \I__7748\ : ClkMux
    port map (
            O => \N__32024\,
            I => \N__31684\
        );

    \I__7747\ : ClkMux
    port map (
            O => \N__32023\,
            I => \N__31684\
        );

    \I__7746\ : ClkMux
    port map (
            O => \N__32022\,
            I => \N__31684\
        );

    \I__7745\ : ClkMux
    port map (
            O => \N__32021\,
            I => \N__31684\
        );

    \I__7744\ : ClkMux
    port map (
            O => \N__32020\,
            I => \N__31684\
        );

    \I__7743\ : ClkMux
    port map (
            O => \N__32019\,
            I => \N__31684\
        );

    \I__7742\ : ClkMux
    port map (
            O => \N__32018\,
            I => \N__31684\
        );

    \I__7741\ : ClkMux
    port map (
            O => \N__32017\,
            I => \N__31684\
        );

    \I__7740\ : ClkMux
    port map (
            O => \N__32016\,
            I => \N__31684\
        );

    \I__7739\ : ClkMux
    port map (
            O => \N__32015\,
            I => \N__31684\
        );

    \I__7738\ : ClkMux
    port map (
            O => \N__32014\,
            I => \N__31684\
        );

    \I__7737\ : ClkMux
    port map (
            O => \N__32013\,
            I => \N__31684\
        );

    \I__7736\ : ClkMux
    port map (
            O => \N__32012\,
            I => \N__31684\
        );

    \I__7735\ : ClkMux
    port map (
            O => \N__32011\,
            I => \N__31684\
        );

    \I__7734\ : ClkMux
    port map (
            O => \N__32010\,
            I => \N__31684\
        );

    \I__7733\ : ClkMux
    port map (
            O => \N__32009\,
            I => \N__31684\
        );

    \I__7732\ : ClkMux
    port map (
            O => \N__32008\,
            I => \N__31684\
        );

    \I__7731\ : ClkMux
    port map (
            O => \N__32007\,
            I => \N__31684\
        );

    \I__7730\ : ClkMux
    port map (
            O => \N__32006\,
            I => \N__31684\
        );

    \I__7729\ : ClkMux
    port map (
            O => \N__32005\,
            I => \N__31684\
        );

    \I__7728\ : ClkMux
    port map (
            O => \N__32004\,
            I => \N__31684\
        );

    \I__7727\ : ClkMux
    port map (
            O => \N__32003\,
            I => \N__31684\
        );

    \I__7726\ : ClkMux
    port map (
            O => \N__32002\,
            I => \N__31684\
        );

    \I__7725\ : ClkMux
    port map (
            O => \N__32001\,
            I => \N__31684\
        );

    \I__7724\ : ClkMux
    port map (
            O => \N__32000\,
            I => \N__31684\
        );

    \I__7723\ : ClkMux
    port map (
            O => \N__31999\,
            I => \N__31684\
        );

    \I__7722\ : ClkMux
    port map (
            O => \N__31998\,
            I => \N__31684\
        );

    \I__7721\ : ClkMux
    port map (
            O => \N__31997\,
            I => \N__31684\
        );

    \I__7720\ : ClkMux
    port map (
            O => \N__31996\,
            I => \N__31684\
        );

    \I__7719\ : ClkMux
    port map (
            O => \N__31995\,
            I => \N__31684\
        );

    \I__7718\ : ClkMux
    port map (
            O => \N__31994\,
            I => \N__31684\
        );

    \I__7717\ : ClkMux
    port map (
            O => \N__31993\,
            I => \N__31684\
        );

    \I__7716\ : ClkMux
    port map (
            O => \N__31992\,
            I => \N__31684\
        );

    \I__7715\ : ClkMux
    port map (
            O => \N__31991\,
            I => \N__31684\
        );

    \I__7714\ : ClkMux
    port map (
            O => \N__31990\,
            I => \N__31684\
        );

    \I__7713\ : ClkMux
    port map (
            O => \N__31989\,
            I => \N__31684\
        );

    \I__7712\ : ClkMux
    port map (
            O => \N__31988\,
            I => \N__31684\
        );

    \I__7711\ : ClkMux
    port map (
            O => \N__31987\,
            I => \N__31684\
        );

    \I__7710\ : ClkMux
    port map (
            O => \N__31986\,
            I => \N__31684\
        );

    \I__7709\ : ClkMux
    port map (
            O => \N__31985\,
            I => \N__31684\
        );

    \I__7708\ : ClkMux
    port map (
            O => \N__31984\,
            I => \N__31684\
        );

    \I__7707\ : ClkMux
    port map (
            O => \N__31983\,
            I => \N__31684\
        );

    \I__7706\ : ClkMux
    port map (
            O => \N__31982\,
            I => \N__31684\
        );

    \I__7705\ : ClkMux
    port map (
            O => \N__31981\,
            I => \N__31684\
        );

    \I__7704\ : ClkMux
    port map (
            O => \N__31980\,
            I => \N__31684\
        );

    \I__7703\ : ClkMux
    port map (
            O => \N__31979\,
            I => \N__31684\
        );

    \I__7702\ : ClkMux
    port map (
            O => \N__31978\,
            I => \N__31684\
        );

    \I__7701\ : ClkMux
    port map (
            O => \N__31977\,
            I => \N__31684\
        );

    \I__7700\ : ClkMux
    port map (
            O => \N__31976\,
            I => \N__31684\
        );

    \I__7699\ : ClkMux
    port map (
            O => \N__31975\,
            I => \N__31684\
        );

    \I__7698\ : ClkMux
    port map (
            O => \N__31974\,
            I => \N__31684\
        );

    \I__7697\ : ClkMux
    port map (
            O => \N__31973\,
            I => \N__31684\
        );

    \I__7696\ : ClkMux
    port map (
            O => \N__31972\,
            I => \N__31684\
        );

    \I__7695\ : ClkMux
    port map (
            O => \N__31971\,
            I => \N__31684\
        );

    \I__7694\ : ClkMux
    port map (
            O => \N__31970\,
            I => \N__31684\
        );

    \I__7693\ : ClkMux
    port map (
            O => \N__31969\,
            I => \N__31684\
        );

    \I__7692\ : ClkMux
    port map (
            O => \N__31968\,
            I => \N__31684\
        );

    \I__7691\ : ClkMux
    port map (
            O => \N__31967\,
            I => \N__31684\
        );

    \I__7690\ : ClkMux
    port map (
            O => \N__31966\,
            I => \N__31684\
        );

    \I__7689\ : ClkMux
    port map (
            O => \N__31965\,
            I => \N__31684\
        );

    \I__7688\ : ClkMux
    port map (
            O => \N__31964\,
            I => \N__31684\
        );

    \I__7687\ : ClkMux
    port map (
            O => \N__31963\,
            I => \N__31684\
        );

    \I__7686\ : ClkMux
    port map (
            O => \N__31962\,
            I => \N__31684\
        );

    \I__7685\ : ClkMux
    port map (
            O => \N__31961\,
            I => \N__31684\
        );

    \I__7684\ : ClkMux
    port map (
            O => \N__31960\,
            I => \N__31684\
        );

    \I__7683\ : ClkMux
    port map (
            O => \N__31959\,
            I => \N__31684\
        );

    \I__7682\ : ClkMux
    port map (
            O => \N__31958\,
            I => \N__31684\
        );

    \I__7681\ : ClkMux
    port map (
            O => \N__31957\,
            I => \N__31684\
        );

    \I__7680\ : ClkMux
    port map (
            O => \N__31956\,
            I => \N__31684\
        );

    \I__7679\ : ClkMux
    port map (
            O => \N__31955\,
            I => \N__31684\
        );

    \I__7678\ : ClkMux
    port map (
            O => \N__31954\,
            I => \N__31684\
        );

    \I__7677\ : ClkMux
    port map (
            O => \N__31953\,
            I => \N__31684\
        );

    \I__7676\ : ClkMux
    port map (
            O => \N__31952\,
            I => \N__31684\
        );

    \I__7675\ : ClkMux
    port map (
            O => \N__31951\,
            I => \N__31684\
        );

    \I__7674\ : ClkMux
    port map (
            O => \N__31950\,
            I => \N__31684\
        );

    \I__7673\ : ClkMux
    port map (
            O => \N__31949\,
            I => \N__31684\
        );

    \I__7672\ : ClkMux
    port map (
            O => \N__31948\,
            I => \N__31684\
        );

    \I__7671\ : ClkMux
    port map (
            O => \N__31947\,
            I => \N__31684\
        );

    \I__7670\ : ClkMux
    port map (
            O => \N__31946\,
            I => \N__31684\
        );

    \I__7669\ : ClkMux
    port map (
            O => \N__31945\,
            I => \N__31684\
        );

    \I__7668\ : ClkMux
    port map (
            O => \N__31944\,
            I => \N__31684\
        );

    \I__7667\ : ClkMux
    port map (
            O => \N__31943\,
            I => \N__31684\
        );

    \I__7666\ : ClkMux
    port map (
            O => \N__31942\,
            I => \N__31684\
        );

    \I__7665\ : ClkMux
    port map (
            O => \N__31941\,
            I => \N__31684\
        );

    \I__7664\ : ClkMux
    port map (
            O => \N__31940\,
            I => \N__31684\
        );

    \I__7663\ : ClkMux
    port map (
            O => \N__31939\,
            I => \N__31684\
        );

    \I__7662\ : ClkMux
    port map (
            O => \N__31938\,
            I => \N__31684\
        );

    \I__7661\ : ClkMux
    port map (
            O => \N__31937\,
            I => \N__31684\
        );

    \I__7660\ : GlobalMux
    port map (
            O => \N__31684\,
            I => \N__31681\
        );

    \I__7659\ : gio2CtrlBuf
    port map (
            O => \N__31681\,
            I => clk_0_c_g
        );

    \I__7658\ : CEMux
    port map (
            O => \N__31678\,
            I => \N__31673\
        );

    \I__7657\ : CEMux
    port map (
            O => \N__31677\,
            I => \N__31670\
        );

    \I__7656\ : CEMux
    port map (
            O => \N__31676\,
            I => \N__31665\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__31673\,
            I => \N__31660\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__31670\,
            I => \N__31660\
        );

    \I__7653\ : CEMux
    port map (
            O => \N__31669\,
            I => \N__31657\
        );

    \I__7652\ : CEMux
    port map (
            O => \N__31668\,
            I => \N__31654\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__31665\,
            I => \N__31651\
        );

    \I__7650\ : Span4Mux_v
    port map (
            O => \N__31660\,
            I => \N__31648\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__31657\,
            I => \N__31643\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__31654\,
            I => \N__31643\
        );

    \I__7647\ : Odrv4
    port map (
            O => \N__31651\,
            I => \M_this_data_count_qe_0_i\
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__31648\,
            I => \M_this_data_count_qe_0_i\
        );

    \I__7645\ : Odrv4
    port map (
            O => \N__31643\,
            I => \M_this_data_count_qe_0_i\
        );

    \I__7644\ : InMux
    port map (
            O => \N__31636\,
            I => \N__31631\
        );

    \I__7643\ : InMux
    port map (
            O => \N__31635\,
            I => \N__31628\
        );

    \I__7642\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31625\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__31631\,
            I => \N__31622\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__31628\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__31625\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__7638\ : Odrv4
    port map (
            O => \N__31622\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__7637\ : CascadeMux
    port map (
            O => \N__31615\,
            I => \N__31612\
        );

    \I__7636\ : InMux
    port map (
            O => \N__31612\,
            I => \N__31607\
        );

    \I__7635\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31604\
        );

    \I__7634\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31601\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__31607\,
            I => \N__31598\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__31604\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__31601\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__7630\ : Odrv4
    port map (
            O => \N__31598\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__7629\ : CascadeMux
    port map (
            O => \N__31591\,
            I => \N__31586\
        );

    \I__7628\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31583\
        );

    \I__7627\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31580\
        );

    \I__7626\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31577\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__31583\,
            I => \N__31574\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__31580\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__31577\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__7622\ : Odrv4
    port map (
            O => \N__31574\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__7621\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31563\
        );

    \I__7620\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31560\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__31563\,
            I => \N__31557\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__31560\,
            I => \N__31552\
        );

    \I__7617\ : Span4Mux_v
    port map (
            O => \N__31557\,
            I => \N__31552\
        );

    \I__7616\ : Span4Mux_v
    port map (
            O => \N__31552\,
            I => \N__31549\
        );

    \I__7615\ : Odrv4
    port map (
            O => \N__31549\,
            I => \M_this_state_d88_10\
        );

    \I__7614\ : CascadeMux
    port map (
            O => \N__31546\,
            I => \N__31541\
        );

    \I__7613\ : InMux
    port map (
            O => \N__31545\,
            I => \N__31538\
        );

    \I__7612\ : InMux
    port map (
            O => \N__31544\,
            I => \N__31534\
        );

    \I__7611\ : InMux
    port map (
            O => \N__31541\,
            I => \N__31531\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__31538\,
            I => \N__31528\
        );

    \I__7609\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31525\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__31534\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__31531\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__7606\ : Odrv4
    port map (
            O => \N__31528\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__31525\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__7604\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31509\
        );

    \I__7603\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31509\
        );

    \I__7602\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31502\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__31509\,
            I => \N__31499\
        );

    \I__7600\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31490\
        );

    \I__7599\ : InMux
    port map (
            O => \N__31507\,
            I => \N__31490\
        );

    \I__7598\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31490\
        );

    \I__7597\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31490\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__31502\,
            I => \N__31487\
        );

    \I__7595\ : Odrv4
    port map (
            O => \N__31499\,
            I => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__31490\,
            I => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8\
        );

    \I__7593\ : Odrv4
    port map (
            O => \N__31487\,
            I => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8\
        );

    \I__7592\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31477\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__31477\,
            I => \N__31474\
        );

    \I__7590\ : Odrv4
    port map (
            O => \N__31474\,
            I => \this_vga_signals.M_this_data_count_q_3_amZ0Z_10\
        );

    \I__7589\ : InMux
    port map (
            O => \N__31471\,
            I => \N__31468\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__31468\,
            I => \N__31465\
        );

    \I__7587\ : Span4Mux_s2_v
    port map (
            O => \N__31465\,
            I => \N__31462\
        );

    \I__7586\ : Span4Mux_v
    port map (
            O => \N__31462\,
            I => \N__31459\
        );

    \I__7585\ : Odrv4
    port map (
            O => \N__31459\,
            I => \M_this_map_ram_write_data_6\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__31456\,
            I => \N__31453\
        );

    \I__7583\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31450\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__31450\,
            I => \M_this_data_count_q_s_11\
        );

    \I__7581\ : InMux
    port map (
            O => \N__31447\,
            I => \N__31444\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__31444\,
            I => \M_this_data_count_q_s_12\
        );

    \I__7579\ : CascadeMux
    port map (
            O => \N__31441\,
            I => \N_518_cascade_\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__31438\,
            I => \N__31433\
        );

    \I__7577\ : InMux
    port map (
            O => \N__31437\,
            I => \N__31430\
        );

    \I__7576\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31427\
        );

    \I__7575\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31424\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__31430\,
            I => \N__31421\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__31427\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__31424\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__7571\ : Odrv4
    port map (
            O => \N__31421\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__7570\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31411\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__31411\,
            I => \M_this_data_count_q_s_14\
        );

    \I__7568\ : CascadeMux
    port map (
            O => \N__31408\,
            I => \N_520_cascade_\
        );

    \I__7567\ : CascadeMux
    port map (
            O => \N__31405\,
            I => \N__31400\
        );

    \I__7566\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31397\
        );

    \I__7565\ : InMux
    port map (
            O => \N__31403\,
            I => \N__31394\
        );

    \I__7564\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31391\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31388\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__31394\,
            I => \M_this_data_count_qZ0Z_14\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__31391\,
            I => \M_this_data_count_qZ0Z_14\
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__31388\,
            I => \M_this_data_count_qZ0Z_14\
        );

    \I__7559\ : InMux
    port map (
            O => \N__31381\,
            I => \N__31378\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__31378\,
            I => \M_this_data_count_q_s_15\
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__31375\,
            I => \N_521_cascade_\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__31372\,
            I => \N__31369\
        );

    \I__7555\ : InMux
    port map (
            O => \N__31369\,
            I => \N__31364\
        );

    \I__7554\ : InMux
    port map (
            O => \N__31368\,
            I => \N__31361\
        );

    \I__7553\ : InMux
    port map (
            O => \N__31367\,
            I => \N__31358\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__31364\,
            I => \N__31355\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__31361\,
            I => \M_this_data_count_qZ0Z_15\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__31358\,
            I => \M_this_data_count_qZ0Z_15\
        );

    \I__7549\ : Odrv4
    port map (
            O => \N__31355\,
            I => \M_this_data_count_qZ0Z_15\
        );

    \I__7548\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31345\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__31345\,
            I => \N_517\
        );

    \I__7546\ : InMux
    port map (
            O => \N__31342\,
            I => \N__31339\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__31339\,
            I => \N__31336\
        );

    \I__7544\ : Span4Mux_v
    port map (
            O => \N__31336\,
            I => \N__31333\
        );

    \I__7543\ : Span4Mux_h
    port map (
            O => \N__31333\,
            I => \N__31330\
        );

    \I__7542\ : Odrv4
    port map (
            O => \N__31330\,
            I => \this_vga_signals.M_this_data_count_q_3_bmZ0Z_10\
        );

    \I__7541\ : CascadeMux
    port map (
            O => \N__31327\,
            I => \N__31324\
        );

    \I__7540\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31320\
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__31323\,
            I => \N__31313\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__31320\,
            I => \N__31310\
        );

    \I__7537\ : InMux
    port map (
            O => \N__31319\,
            I => \N__31307\
        );

    \I__7536\ : InMux
    port map (
            O => \N__31318\,
            I => \N__31304\
        );

    \I__7535\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31301\
        );

    \I__7534\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31296\
        );

    \I__7533\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31296\
        );

    \I__7532\ : Span4Mux_v
    port map (
            O => \N__31310\,
            I => \N__31290\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__31307\,
            I => \N__31290\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__31304\,
            I => \N__31287\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__31301\,
            I => \N__31284\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__31296\,
            I => \N__31281\
        );

    \I__7527\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31278\
        );

    \I__7526\ : Span4Mux_h
    port map (
            O => \N__31290\,
            I => \N__31275\
        );

    \I__7525\ : Span4Mux_h
    port map (
            O => \N__31287\,
            I => \N__31272\
        );

    \I__7524\ : Span4Mux_h
    port map (
            O => \N__31284\,
            I => \N__31267\
        );

    \I__7523\ : Span4Mux_h
    port map (
            O => \N__31281\,
            I => \N__31267\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__31278\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__7521\ : Odrv4
    port map (
            O => \N__31275\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__7520\ : Odrv4
    port map (
            O => \N__31272\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__31267\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__7518\ : CascadeMux
    port map (
            O => \N__31258\,
            I => \N__31255\
        );

    \I__7517\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31249\
        );

    \I__7516\ : InMux
    port map (
            O => \N__31254\,
            I => \N__31246\
        );

    \I__7515\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31243\
        );

    \I__7514\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31240\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__31249\,
            I => \N__31237\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__31246\,
            I => \N__31232\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__31243\,
            I => \N__31232\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__31240\,
            I => \N__31228\
        );

    \I__7509\ : Span4Mux_h
    port map (
            O => \N__31237\,
            I => \N__31223\
        );

    \I__7508\ : Span4Mux_v
    port map (
            O => \N__31232\,
            I => \N__31223\
        );

    \I__7507\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31220\
        );

    \I__7506\ : Span12Mux_h
    port map (
            O => \N__31228\,
            I => \N__31217\
        );

    \I__7505\ : Odrv4
    port map (
            O => \N__31223\,
            I => \N_391_0\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__31220\,
            I => \N_391_0\
        );

    \I__7503\ : Odrv12
    port map (
            O => \N__31217\,
            I => \N_391_0\
        );

    \I__7502\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31207\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__31207\,
            I => \this_vga_signals.un1_M_this_state_q_18Z0Z_1\
        );

    \I__7500\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31194\
        );

    \I__7499\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31194\
        );

    \I__7498\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31191\
        );

    \I__7497\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31188\
        );

    \I__7496\ : InMux
    port map (
            O => \N__31200\,
            I => \N__31185\
        );

    \I__7495\ : CascadeMux
    port map (
            O => \N__31199\,
            I => \N__31182\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31179\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__31191\,
            I => \N__31176\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__31188\,
            I => \N__31171\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__31185\,
            I => \N__31171\
        );

    \I__7490\ : InMux
    port map (
            O => \N__31182\,
            I => \N__31168\
        );

    \I__7489\ : Span4Mux_v
    port map (
            O => \N__31179\,
            I => \N__31165\
        );

    \I__7488\ : Span4Mux_v
    port map (
            O => \N__31176\,
            I => \N__31162\
        );

    \I__7487\ : Span4Mux_v
    port map (
            O => \N__31171\,
            I => \N__31159\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__31168\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__7485\ : Odrv4
    port map (
            O => \N__31165\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__31162\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__7483\ : Odrv4
    port map (
            O => \N__31159\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__7482\ : InMux
    port map (
            O => \N__31150\,
            I => \N__31143\
        );

    \I__7481\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31143\
        );

    \I__7480\ : CascadeMux
    port map (
            O => \N__31148\,
            I => \N__31140\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__31143\,
            I => \N__31137\
        );

    \I__7478\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31134\
        );

    \I__7477\ : Span4Mux_v
    port map (
            O => \N__31137\,
            I => \N__31129\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31129\
        );

    \I__7475\ : Span4Mux_h
    port map (
            O => \N__31129\,
            I => \N__31125\
        );

    \I__7474\ : InMux
    port map (
            O => \N__31128\,
            I => \N__31122\
        );

    \I__7473\ : Odrv4
    port map (
            O => \N__31125\,
            I => \this_vga_signals.N_387_0\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__31122\,
            I => \this_vga_signals.N_387_0\
        );

    \I__7471\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31108\
        );

    \I__7470\ : InMux
    port map (
            O => \N__31116\,
            I => \N__31108\
        );

    \I__7469\ : InMux
    port map (
            O => \N__31115\,
            I => \N__31108\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__31108\,
            I => \N__31104\
        );

    \I__7467\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31097\
        );

    \I__7466\ : Span4Mux_h
    port map (
            O => \N__31104\,
            I => \N__31094\
        );

    \I__7465\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31091\
        );

    \I__7464\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31088\
        );

    \I__7463\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31083\
        );

    \I__7462\ : InMux
    port map (
            O => \N__31100\,
            I => \N__31083\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__31097\,
            I => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0\
        );

    \I__7460\ : Odrv4
    port map (
            O => \N__31094\,
            I => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__31091\,
            I => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__31088\,
            I => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__31083\,
            I => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0\
        );

    \I__7456\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31069\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__31069\,
            I => \N_513\
        );

    \I__7454\ : CascadeMux
    port map (
            O => \N__31066\,
            I => \N__31063\
        );

    \I__7453\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31060\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__31060\,
            I => \M_this_data_count_q_s_7\
        );

    \I__7451\ : CascadeMux
    port map (
            O => \N__31057\,
            I => \N__31054\
        );

    \I__7450\ : InMux
    port map (
            O => \N__31054\,
            I => \N__31049\
        );

    \I__7449\ : InMux
    port map (
            O => \N__31053\,
            I => \N__31046\
        );

    \I__7448\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31043\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__31049\,
            I => \N__31040\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__31046\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__31043\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__7444\ : Odrv4
    port map (
            O => \N__31040\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__7443\ : InMux
    port map (
            O => \N__31033\,
            I => \N__31030\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__31030\,
            I => \M_this_data_count_q_s_8\
        );

    \I__7441\ : CascadeMux
    port map (
            O => \N__31027\,
            I => \N_514_cascade_\
        );

    \I__7440\ : InMux
    port map (
            O => \N__31024\,
            I => \N__31021\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__31021\,
            I => \M_this_data_count_q_s_9\
        );

    \I__7438\ : CascadeMux
    port map (
            O => \N__31018\,
            I => \N_515_cascade_\
        );

    \I__7437\ : InMux
    port map (
            O => \N__31015\,
            I => \N__31012\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__31012\,
            I => \N__31009\
        );

    \I__7435\ : Span4Mux_v
    port map (
            O => \N__31009\,
            I => \N__31006\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__31006\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_7\
        );

    \I__7433\ : CascadeMux
    port map (
            O => \N__31003\,
            I => \this_vga_signals.M_this_external_address_d_8_mZ0Z_7_cascade_\
        );

    \I__7432\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30997\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__30997\,
            I => \un1_M_this_external_address_q_cry_6_c_RNIS2NBZ0\
        );

    \I__7430\ : IoInMux
    port map (
            O => \N__30994\,
            I => \N__30991\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__30991\,
            I => \N__30988\
        );

    \I__7428\ : Span4Mux_s1_h
    port map (
            O => \N__30988\,
            I => \N__30985\
        );

    \I__7427\ : Span4Mux_v
    port map (
            O => \N__30985\,
            I => \N__30982\
        );

    \I__7426\ : Span4Mux_v
    port map (
            O => \N__30982\,
            I => \N__30979\
        );

    \I__7425\ : Span4Mux_h
    port map (
            O => \N__30979\,
            I => \N__30975\
        );

    \I__7424\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30972\
        );

    \I__7423\ : Span4Mux_h
    port map (
            O => \N__30975\,
            I => \N__30966\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__30972\,
            I => \N__30966\
        );

    \I__7421\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30962\
        );

    \I__7420\ : Span4Mux_v
    port map (
            O => \N__30966\,
            I => \N__30959\
        );

    \I__7419\ : InMux
    port map (
            O => \N__30965\,
            I => \N__30956\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__30962\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__7417\ : Odrv4
    port map (
            O => \N__30959\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__30956\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__7415\ : CascadeMux
    port map (
            O => \N__30949\,
            I => \this_vga_signals.M_this_external_address_d_5_mZ0Z_10_cascade_\
        );

    \I__7414\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30943\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__30943\,
            I => \un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0\
        );

    \I__7412\ : IoInMux
    port map (
            O => \N__30940\,
            I => \N__30937\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__30937\,
            I => \N__30933\
        );

    \I__7410\ : InMux
    port map (
            O => \N__30936\,
            I => \N__30929\
        );

    \I__7409\ : Span12Mux_s11_v
    port map (
            O => \N__30933\,
            I => \N__30925\
        );

    \I__7408\ : InMux
    port map (
            O => \N__30932\,
            I => \N__30922\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__30929\,
            I => \N__30919\
        );

    \I__7406\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30916\
        );

    \I__7405\ : Odrv12
    port map (
            O => \N__30925\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__30922\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__7403\ : Odrv4
    port map (
            O => \N__30919\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__30916\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__7401\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30904\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__30904\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_10\
        );

    \I__7399\ : IoInMux
    port map (
            O => \N__30901\,
            I => \N__30898\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__30898\,
            I => \N__30895\
        );

    \I__7397\ : Span4Mux_s2_v
    port map (
            O => \N__30895\,
            I => \N__30892\
        );

    \I__7396\ : Span4Mux_v
    port map (
            O => \N__30892\,
            I => \N__30888\
        );

    \I__7395\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30884\
        );

    \I__7394\ : Span4Mux_v
    port map (
            O => \N__30888\,
            I => \N__30880\
        );

    \I__7393\ : InMux
    port map (
            O => \N__30887\,
            I => \N__30877\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__30884\,
            I => \N__30874\
        );

    \I__7391\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30871\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__30880\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__30877\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__7388\ : Odrv12
    port map (
            O => \N__30874\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__30871\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__7386\ : CascadeMux
    port map (
            O => \N__30862\,
            I => \N__30853\
        );

    \I__7385\ : CascadeMux
    port map (
            O => \N__30861\,
            I => \N__30849\
        );

    \I__7384\ : InMux
    port map (
            O => \N__30860\,
            I => \N__30844\
        );

    \I__7383\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30835\
        );

    \I__7382\ : InMux
    port map (
            O => \N__30858\,
            I => \N__30828\
        );

    \I__7381\ : InMux
    port map (
            O => \N__30857\,
            I => \N__30828\
        );

    \I__7380\ : InMux
    port map (
            O => \N__30856\,
            I => \N__30828\
        );

    \I__7379\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30823\
        );

    \I__7378\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30823\
        );

    \I__7377\ : InMux
    port map (
            O => \N__30849\,
            I => \N__30818\
        );

    \I__7376\ : InMux
    port map (
            O => \N__30848\,
            I => \N__30818\
        );

    \I__7375\ : InMux
    port map (
            O => \N__30847\,
            I => \N__30815\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__30844\,
            I => \N__30812\
        );

    \I__7373\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30809\
        );

    \I__7372\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30806\
        );

    \I__7371\ : InMux
    port map (
            O => \N__30841\,
            I => \N__30801\
        );

    \I__7370\ : InMux
    port map (
            O => \N__30840\,
            I => \N__30801\
        );

    \I__7369\ : InMux
    port map (
            O => \N__30839\,
            I => \N__30797\
        );

    \I__7368\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30794\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__30835\,
            I => \N__30785\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__30828\,
            I => \N__30785\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__30823\,
            I => \N__30785\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__30818\,
            I => \N__30785\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__30815\,
            I => \N__30781\
        );

    \I__7362\ : Span4Mux_h
    port map (
            O => \N__30812\,
            I => \N__30778\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__30809\,
            I => \N__30771\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__30806\,
            I => \N__30771\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__30801\,
            I => \N__30771\
        );

    \I__7358\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30768\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__30797\,
            I => \N__30765\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30760\
        );

    \I__7355\ : Span4Mux_v
    port map (
            O => \N__30785\,
            I => \N__30760\
        );

    \I__7354\ : InMux
    port map (
            O => \N__30784\,
            I => \N__30757\
        );

    \I__7353\ : Span4Mux_h
    port map (
            O => \N__30781\,
            I => \N__30745\
        );

    \I__7352\ : Span4Mux_v
    port map (
            O => \N__30778\,
            I => \N__30745\
        );

    \I__7351\ : Span4Mux_v
    port map (
            O => \N__30771\,
            I => \N__30745\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__30768\,
            I => \N__30745\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__30765\,
            I => \N__30740\
        );

    \I__7348\ : Span4Mux_v
    port map (
            O => \N__30760\,
            I => \N__30740\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__30757\,
            I => \N__30737\
        );

    \I__7346\ : InMux
    port map (
            O => \N__30756\,
            I => \N__30734\
        );

    \I__7345\ : InMux
    port map (
            O => \N__30755\,
            I => \N__30731\
        );

    \I__7344\ : InMux
    port map (
            O => \N__30754\,
            I => \N__30728\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__30745\,
            I => \N__30725\
        );

    \I__7342\ : Span4Mux_h
    port map (
            O => \N__30740\,
            I => \N__30720\
        );

    \I__7341\ : Span4Mux_h
    port map (
            O => \N__30737\,
            I => \N__30720\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__30734\,
            I => \N__30715\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__30731\,
            I => \N__30715\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__30728\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__7337\ : Odrv4
    port map (
            O => \N__30725\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__7336\ : Odrv4
    port map (
            O => \N__30720\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__7335\ : Odrv12
    port map (
            O => \N__30715\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__7334\ : InMux
    port map (
            O => \N__30706\,
            I => \N__30703\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__30703\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_9\
        );

    \I__7332\ : InMux
    port map (
            O => \N__30700\,
            I => \N__30692\
        );

    \I__7331\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30689\
        );

    \I__7330\ : CascadeMux
    port map (
            O => \N__30698\,
            I => \N__30686\
        );

    \I__7329\ : InMux
    port map (
            O => \N__30697\,
            I => \N__30677\
        );

    \I__7328\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30677\
        );

    \I__7327\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30672\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__30692\,
            I => \N__30664\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__30689\,
            I => \N__30664\
        );

    \I__7324\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30661\
        );

    \I__7323\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30658\
        );

    \I__7322\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30655\
        );

    \I__7321\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30652\
        );

    \I__7320\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30649\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__30677\,
            I => \N__30645\
        );

    \I__7318\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30640\
        );

    \I__7317\ : InMux
    port map (
            O => \N__30675\,
            I => \N__30640\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__30672\,
            I => \N__30637\
        );

    \I__7315\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30633\
        );

    \I__7314\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30630\
        );

    \I__7313\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30627\
        );

    \I__7312\ : Span4Mux_v
    port map (
            O => \N__30664\,
            I => \N__30618\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__30661\,
            I => \N__30618\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__30658\,
            I => \N__30618\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30618\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__30652\,
            I => \N__30613\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30613\
        );

    \I__7306\ : CascadeMux
    port map (
            O => \N__30648\,
            I => \N__30610\
        );

    \I__7305\ : Span4Mux_v
    port map (
            O => \N__30645\,
            I => \N__30602\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__30640\,
            I => \N__30602\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__30637\,
            I => \N__30602\
        );

    \I__7302\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30599\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__30633\,
            I => \N__30592\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__30630\,
            I => \N__30592\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__30627\,
            I => \N__30585\
        );

    \I__7298\ : Span4Mux_v
    port map (
            O => \N__30618\,
            I => \N__30585\
        );

    \I__7297\ : Span4Mux_v
    port map (
            O => \N__30613\,
            I => \N__30585\
        );

    \I__7296\ : InMux
    port map (
            O => \N__30610\,
            I => \N__30582\
        );

    \I__7295\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30579\
        );

    \I__7294\ : Span4Mux_h
    port map (
            O => \N__30602\,
            I => \N__30573\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__30599\,
            I => \N__30573\
        );

    \I__7292\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30570\
        );

    \I__7291\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30567\
        );

    \I__7290\ : Span12Mux_h
    port map (
            O => \N__30592\,
            I => \N__30564\
        );

    \I__7289\ : Span4Mux_h
    port map (
            O => \N__30585\,
            I => \N__30561\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__30582\,
            I => \N__30556\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__30579\,
            I => \N__30556\
        );

    \I__7286\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30553\
        );

    \I__7285\ : Span4Mux_h
    port map (
            O => \N__30573\,
            I => \N__30550\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__30570\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__30567\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__7282\ : Odrv12
    port map (
            O => \N__30564\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__7281\ : Odrv4
    port map (
            O => \N__30561\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__7280\ : Odrv4
    port map (
            O => \N__30556\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__30553\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__7278\ : Odrv4
    port map (
            O => \N__30550\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__7277\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30532\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__30532\,
            I => \this_vga_signals.M_this_external_address_d_5_mZ0Z_12\
        );

    \I__7275\ : InMux
    port map (
            O => \N__30529\,
            I => \N__30515\
        );

    \I__7274\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30510\
        );

    \I__7273\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30510\
        );

    \I__7272\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30503\
        );

    \I__7271\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30503\
        );

    \I__7270\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30503\
        );

    \I__7269\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30496\
        );

    \I__7268\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30496\
        );

    \I__7267\ : InMux
    port map (
            O => \N__30521\,
            I => \N__30496\
        );

    \I__7266\ : InMux
    port map (
            O => \N__30520\,
            I => \N__30489\
        );

    \I__7265\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30489\
        );

    \I__7264\ : InMux
    port map (
            O => \N__30518\,
            I => \N__30489\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__30515\,
            I => \N__30476\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__30510\,
            I => \N__30476\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__30503\,
            I => \N__30476\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__30496\,
            I => \N__30476\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__30489\,
            I => \N__30476\
        );

    \I__7258\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30471\
        );

    \I__7257\ : InMux
    port map (
            O => \N__30487\,
            I => \N__30471\
        );

    \I__7256\ : Span4Mux_v
    port map (
            O => \N__30476\,
            I => \N__30467\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__30471\,
            I => \N__30464\
        );

    \I__7254\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30461\
        );

    \I__7253\ : Odrv4
    port map (
            O => \N__30467\,
            I => \this_vga_signals.un1_M_this_state_q_21_0\
        );

    \I__7252\ : Odrv4
    port map (
            O => \N__30464\,
            I => \this_vga_signals.un1_M_this_state_q_21_0\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__30461\,
            I => \this_vga_signals.un1_M_this_state_q_21_0\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__30454\,
            I => \N__30451\
        );

    \I__7249\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30448\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__30448\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_12\
        );

    \I__7247\ : InMux
    port map (
            O => \N__30445\,
            I => \N__30442\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__30442\,
            I => \N__30439\
        );

    \I__7245\ : Odrv4
    port map (
            O => \N__30439\,
            I => \un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0\
        );

    \I__7244\ : IoInMux
    port map (
            O => \N__30436\,
            I => \N__30433\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__30433\,
            I => \N__30430\
        );

    \I__7242\ : IoSpan4Mux
    port map (
            O => \N__30430\,
            I => \N__30427\
        );

    \I__7241\ : Span4Mux_s2_h
    port map (
            O => \N__30427\,
            I => \N__30423\
        );

    \I__7240\ : InMux
    port map (
            O => \N__30426\,
            I => \N__30418\
        );

    \I__7239\ : Span4Mux_h
    port map (
            O => \N__30423\,
            I => \N__30415\
        );

    \I__7238\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30410\
        );

    \I__7237\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30410\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__30418\,
            I => \N__30407\
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__30415\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__30410\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__30407\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__7232\ : InMux
    port map (
            O => \N__30400\,
            I => \N__30397\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30394\
        );

    \I__7230\ : Odrv4
    port map (
            O => \N__30394\,
            I => \M_this_map_ram_write_data_3\
        );

    \I__7229\ : InMux
    port map (
            O => \N__30391\,
            I => \N__30388\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__30388\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_1\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__30385\,
            I => \this_vga_signals.M_this_external_address_d_8_mZ0Z_1_cascade_\
        );

    \I__7226\ : InMux
    port map (
            O => \N__30382\,
            I => \N__30379\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__30379\,
            I => \un1_M_this_external_address_q_cry_0_c_RNIGGGBZ0\
        );

    \I__7224\ : IoInMux
    port map (
            O => \N__30376\,
            I => \N__30373\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__30373\,
            I => \N__30370\
        );

    \I__7222\ : IoSpan4Mux
    port map (
            O => \N__30370\,
            I => \N__30367\
        );

    \I__7221\ : Sp12to4
    port map (
            O => \N__30367\,
            I => \N__30364\
        );

    \I__7220\ : Span12Mux_v
    port map (
            O => \N__30364\,
            I => \N__30358\
        );

    \I__7219\ : InMux
    port map (
            O => \N__30363\,
            I => \N__30355\
        );

    \I__7218\ : InMux
    port map (
            O => \N__30362\,
            I => \N__30352\
        );

    \I__7217\ : InMux
    port map (
            O => \N__30361\,
            I => \N__30349\
        );

    \I__7216\ : Odrv12
    port map (
            O => \N__30358\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__30355\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__30352\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__30349\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__7212\ : InMux
    port map (
            O => \N__30340\,
            I => \N__30337\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__30337\,
            I => \N__30334\
        );

    \I__7210\ : Span4Mux_v
    port map (
            O => \N__30334\,
            I => \N__30331\
        );

    \I__7209\ : Span4Mux_h
    port map (
            O => \N__30331\,
            I => \N__30328\
        );

    \I__7208\ : Odrv4
    port map (
            O => \N__30328\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_2\
        );

    \I__7207\ : CascadeMux
    port map (
            O => \N__30325\,
            I => \this_vga_signals.M_this_external_address_d_8_mZ0Z_2_cascade_\
        );

    \I__7206\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30319\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__30319\,
            I => \un1_M_this_external_address_q_cry_1_c_RNIIJHBZ0\
        );

    \I__7204\ : IoInMux
    port map (
            O => \N__30316\,
            I => \N__30313\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__30313\,
            I => \N__30310\
        );

    \I__7202\ : Span4Mux_s0_v
    port map (
            O => \N__30310\,
            I => \N__30307\
        );

    \I__7201\ : Sp12to4
    port map (
            O => \N__30307\,
            I => \N__30303\
        );

    \I__7200\ : InMux
    port map (
            O => \N__30306\,
            I => \N__30300\
        );

    \I__7199\ : Span12Mux_h
    port map (
            O => \N__30303\,
            I => \N__30296\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__30300\,
            I => \N__30293\
        );

    \I__7197\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30289\
        );

    \I__7196\ : Span12Mux_v
    port map (
            O => \N__30296\,
            I => \N__30284\
        );

    \I__7195\ : Span12Mux_v
    port map (
            O => \N__30293\,
            I => \N__30284\
        );

    \I__7194\ : InMux
    port map (
            O => \N__30292\,
            I => \N__30281\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__30289\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__7192\ : Odrv12
    port map (
            O => \N__30284\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__30281\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__7190\ : InMux
    port map (
            O => \N__30274\,
            I => \N__30271\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__30271\,
            I => \N__30268\
        );

    \I__7188\ : Odrv4
    port map (
            O => \N__30268\,
            I => \this_vga_signals.M_this_external_address_d_8_mZ0Z_4\
        );

    \I__7187\ : CascadeMux
    port map (
            O => \N__30265\,
            I => \N__30262\
        );

    \I__7186\ : InMux
    port map (
            O => \N__30262\,
            I => \N__30259\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__30259\,
            I => \N__30256\
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__30256\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_4\
        );

    \I__7183\ : InMux
    port map (
            O => \N__30253\,
            I => \N__30250\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__30250\,
            I => \un1_M_this_external_address_q_cry_3_c_RNIMPJBZ0\
        );

    \I__7181\ : IoInMux
    port map (
            O => \N__30247\,
            I => \N__30244\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__30244\,
            I => \N__30241\
        );

    \I__7179\ : IoSpan4Mux
    port map (
            O => \N__30241\,
            I => \N__30238\
        );

    \I__7178\ : Span4Mux_s3_h
    port map (
            O => \N__30238\,
            I => \N__30233\
        );

    \I__7177\ : InMux
    port map (
            O => \N__30237\,
            I => \N__30228\
        );

    \I__7176\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30228\
        );

    \I__7175\ : Span4Mux_h
    port map (
            O => \N__30233\,
            I => \N__30222\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__30228\,
            I => \N__30222\
        );

    \I__7173\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30219\
        );

    \I__7172\ : Odrv4
    port map (
            O => \N__30222\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__30219\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__7170\ : CascadeMux
    port map (
            O => \N__30214\,
            I => \this_vga_signals.M_this_external_address_d_5_i_mZ0Z_15_cascade_\
        );

    \I__7169\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30208\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__30208\,
            I => \un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0\
        );

    \I__7167\ : IoInMux
    port map (
            O => \N__30205\,
            I => \N__30202\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__30202\,
            I => \N__30199\
        );

    \I__7165\ : Span12Mux_s9_h
    port map (
            O => \N__30199\,
            I => \N__30196\
        );

    \I__7164\ : Span12Mux_v
    port map (
            O => \N__30196\,
            I => \N__30190\
        );

    \I__7163\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30187\
        );

    \I__7162\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30182\
        );

    \I__7161\ : InMux
    port map (
            O => \N__30193\,
            I => \N__30182\
        );

    \I__7160\ : Odrv12
    port map (
            O => \N__30190\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__30187\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__30182\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__7157\ : InMux
    port map (
            O => \N__30175\,
            I => \N__30172\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__30172\,
            I => \this_vga_signals.M_this_external_address_q_i_mZ0Z_15\
        );

    \I__7155\ : InMux
    port map (
            O => \N__30169\,
            I => \M_this_data_count_q_cry_10\
        );

    \I__7154\ : InMux
    port map (
            O => \N__30166\,
            I => \M_this_data_count_q_cry_11\
        );

    \I__7153\ : InMux
    port map (
            O => \N__30163\,
            I => \M_this_data_count_q_cry_12\
        );

    \I__7152\ : SRMux
    port map (
            O => \N__30160\,
            I => \N__30157\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__30157\,
            I => \N__30152\
        );

    \I__7150\ : SRMux
    port map (
            O => \N__30156\,
            I => \N__30149\
        );

    \I__7149\ : SRMux
    port map (
            O => \N__30155\,
            I => \N__30146\
        );

    \I__7148\ : Span4Mux_s2_v
    port map (
            O => \N__30152\,
            I => \N__30141\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__30149\,
            I => \N__30138\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__30146\,
            I => \N__30135\
        );

    \I__7145\ : SRMux
    port map (
            O => \N__30145\,
            I => \N__30132\
        );

    \I__7144\ : IoInMux
    port map (
            O => \N__30144\,
            I => \N__30129\
        );

    \I__7143\ : Span4Mux_h
    port map (
            O => \N__30141\,
            I => \N__30124\
        );

    \I__7142\ : Span4Mux_h
    port map (
            O => \N__30138\,
            I => \N__30124\
        );

    \I__7141\ : Span4Mux_s2_v
    port map (
            O => \N__30135\,
            I => \N__30119\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__30132\,
            I => \N__30119\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__30129\,
            I => \N__30112\
        );

    \I__7138\ : Span4Mux_v
    port map (
            O => \N__30124\,
            I => \N__30107\
        );

    \I__7137\ : Span4Mux_v
    port map (
            O => \N__30119\,
            I => \N__30107\
        );

    \I__7136\ : SRMux
    port map (
            O => \N__30118\,
            I => \N__30103\
        );

    \I__7135\ : SRMux
    port map (
            O => \N__30117\,
            I => \N__30100\
        );

    \I__7134\ : SRMux
    port map (
            O => \N__30116\,
            I => \N__30097\
        );

    \I__7133\ : SRMux
    port map (
            O => \N__30115\,
            I => \N__30094\
        );

    \I__7132\ : IoSpan4Mux
    port map (
            O => \N__30112\,
            I => \N__30086\
        );

    \I__7131\ : Span4Mux_v
    port map (
            O => \N__30107\,
            I => \N__30082\
        );

    \I__7130\ : SRMux
    port map (
            O => \N__30106\,
            I => \N__30079\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__30103\,
            I => \N__30066\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__30100\,
            I => \N__30066\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__30097\,
            I => \N__30061\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__30094\,
            I => \N__30061\
        );

    \I__7125\ : SRMux
    port map (
            O => \N__30093\,
            I => \N__30058\
        );

    \I__7124\ : SRMux
    port map (
            O => \N__30092\,
            I => \N__30055\
        );

    \I__7123\ : SRMux
    port map (
            O => \N__30091\,
            I => \N__30051\
        );

    \I__7122\ : SRMux
    port map (
            O => \N__30090\,
            I => \N__30048\
        );

    \I__7121\ : SRMux
    port map (
            O => \N__30089\,
            I => \N__30045\
        );

    \I__7120\ : Span4Mux_s0_h
    port map (
            O => \N__30086\,
            I => \N__30035\
        );

    \I__7119\ : SRMux
    port map (
            O => \N__30085\,
            I => \N__30032\
        );

    \I__7118\ : Span4Mux_v
    port map (
            O => \N__30082\,
            I => \N__30025\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__30079\,
            I => \N__30025\
        );

    \I__7116\ : SRMux
    port map (
            O => \N__30078\,
            I => \N__30022\
        );

    \I__7115\ : CascadeMux
    port map (
            O => \N__30077\,
            I => \N__30018\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__30076\,
            I => \N__30015\
        );

    \I__7113\ : CascadeMux
    port map (
            O => \N__30075\,
            I => \N__30009\
        );

    \I__7112\ : CascadeMux
    port map (
            O => \N__30074\,
            I => \N__30006\
        );

    \I__7111\ : CascadeMux
    port map (
            O => \N__30073\,
            I => \N__30002\
        );

    \I__7110\ : CascadeMux
    port map (
            O => \N__30072\,
            I => \N__29998\
        );

    \I__7109\ : CascadeMux
    port map (
            O => \N__30071\,
            I => \N__29994\
        );

    \I__7108\ : Span4Mux_v
    port map (
            O => \N__30066\,
            I => \N__29985\
        );

    \I__7107\ : Span4Mux_v
    port map (
            O => \N__30061\,
            I => \N__29985\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__30058\,
            I => \N__29985\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__30055\,
            I => \N__29985\
        );

    \I__7104\ : SRMux
    port map (
            O => \N__30054\,
            I => \N__29982\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__30051\,
            I => \N__29977\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__30048\,
            I => \N__29977\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__30045\,
            I => \N__29974\
        );

    \I__7100\ : SRMux
    port map (
            O => \N__30044\,
            I => \N__29971\
        );

    \I__7099\ : SRMux
    port map (
            O => \N__30043\,
            I => \N__29968\
        );

    \I__7098\ : SRMux
    port map (
            O => \N__30042\,
            I => \N__29963\
        );

    \I__7097\ : SRMux
    port map (
            O => \N__30041\,
            I => \N__29958\
        );

    \I__7096\ : SRMux
    port map (
            O => \N__30040\,
            I => \N__29955\
        );

    \I__7095\ : SRMux
    port map (
            O => \N__30039\,
            I => \N__29952\
        );

    \I__7094\ : SRMux
    port map (
            O => \N__30038\,
            I => \N__29949\
        );

    \I__7093\ : Span4Mux_h
    port map (
            O => \N__30035\,
            I => \N__29942\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__30032\,
            I => \N__29942\
        );

    \I__7091\ : SRMux
    port map (
            O => \N__30031\,
            I => \N__29939\
        );

    \I__7090\ : SRMux
    port map (
            O => \N__30030\,
            I => \N__29936\
        );

    \I__7089\ : Span4Mux_v
    port map (
            O => \N__30025\,
            I => \N__29931\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__30022\,
            I => \N__29928\
        );

    \I__7087\ : InMux
    port map (
            O => \N__30021\,
            I => \N__29913\
        );

    \I__7086\ : InMux
    port map (
            O => \N__30018\,
            I => \N__29913\
        );

    \I__7085\ : InMux
    port map (
            O => \N__30015\,
            I => \N__29913\
        );

    \I__7084\ : InMux
    port map (
            O => \N__30014\,
            I => \N__29913\
        );

    \I__7083\ : InMux
    port map (
            O => \N__30013\,
            I => \N__29913\
        );

    \I__7082\ : InMux
    port map (
            O => \N__30012\,
            I => \N__29913\
        );

    \I__7081\ : InMux
    port map (
            O => \N__30009\,
            I => \N__29913\
        );

    \I__7080\ : InMux
    port map (
            O => \N__30006\,
            I => \N__29898\
        );

    \I__7079\ : InMux
    port map (
            O => \N__30005\,
            I => \N__29898\
        );

    \I__7078\ : InMux
    port map (
            O => \N__30002\,
            I => \N__29898\
        );

    \I__7077\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29898\
        );

    \I__7076\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29898\
        );

    \I__7075\ : InMux
    port map (
            O => \N__29997\,
            I => \N__29898\
        );

    \I__7074\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29898\
        );

    \I__7073\ : Span4Mux_v
    port map (
            O => \N__29985\,
            I => \N__29895\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__29982\,
            I => \N__29892\
        );

    \I__7071\ : Span4Mux_v
    port map (
            O => \N__29977\,
            I => \N__29883\
        );

    \I__7070\ : Span4Mux_h
    port map (
            O => \N__29974\,
            I => \N__29883\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__29971\,
            I => \N__29883\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__29968\,
            I => \N__29883\
        );

    \I__7067\ : SRMux
    port map (
            O => \N__29967\,
            I => \N__29880\
        );

    \I__7066\ : SRMux
    port map (
            O => \N__29966\,
            I => \N__29877\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__29963\,
            I => \N__29873\
        );

    \I__7064\ : SRMux
    port map (
            O => \N__29962\,
            I => \N__29870\
        );

    \I__7063\ : SRMux
    port map (
            O => \N__29961\,
            I => \N__29866\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__29958\,
            I => \N__29863\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__29955\,
            I => \N__29860\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__29952\,
            I => \N__29855\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__29949\,
            I => \N__29855\
        );

    \I__7058\ : SRMux
    port map (
            O => \N__29948\,
            I => \N__29852\
        );

    \I__7057\ : SRMux
    port map (
            O => \N__29947\,
            I => \N__29849\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__29942\,
            I => \N__29843\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__29939\,
            I => \N__29843\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__29936\,
            I => \N__29840\
        );

    \I__7053\ : SRMux
    port map (
            O => \N__29935\,
            I => \N__29837\
        );

    \I__7052\ : IoInMux
    port map (
            O => \N__29934\,
            I => \N__29833\
        );

    \I__7051\ : Span4Mux_v
    port map (
            O => \N__29931\,
            I => \N__29828\
        );

    \I__7050\ : Span4Mux_v
    port map (
            O => \N__29928\,
            I => \N__29828\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__29913\,
            I => \N__29822\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__29898\,
            I => \N__29822\
        );

    \I__7047\ : Span4Mux_v
    port map (
            O => \N__29895\,
            I => \N__29811\
        );

    \I__7046\ : Span4Mux_v
    port map (
            O => \N__29892\,
            I => \N__29811\
        );

    \I__7045\ : Span4Mux_v
    port map (
            O => \N__29883\,
            I => \N__29811\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__29880\,
            I => \N__29811\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__29877\,
            I => \N__29811\
        );

    \I__7042\ : SRMux
    port map (
            O => \N__29876\,
            I => \N__29808\
        );

    \I__7041\ : Span4Mux_v
    port map (
            O => \N__29873\,
            I => \N__29803\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__29870\,
            I => \N__29803\
        );

    \I__7039\ : SRMux
    port map (
            O => \N__29869\,
            I => \N__29800\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29797\
        );

    \I__7037\ : Span4Mux_s3_v
    port map (
            O => \N__29863\,
            I => \N__29786\
        );

    \I__7036\ : Span4Mux_h
    port map (
            O => \N__29860\,
            I => \N__29786\
        );

    \I__7035\ : Span4Mux_s3_v
    port map (
            O => \N__29855\,
            I => \N__29786\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__29852\,
            I => \N__29786\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__29849\,
            I => \N__29786\
        );

    \I__7032\ : SRMux
    port map (
            O => \N__29848\,
            I => \N__29783\
        );

    \I__7031\ : Span4Mux_v
    port map (
            O => \N__29843\,
            I => \N__29776\
        );

    \I__7030\ : Span4Mux_h
    port map (
            O => \N__29840\,
            I => \N__29776\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__29837\,
            I => \N__29776\
        );

    \I__7028\ : SRMux
    port map (
            O => \N__29836\,
            I => \N__29773\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__29833\,
            I => \N__29770\
        );

    \I__7026\ : Span4Mux_h
    port map (
            O => \N__29828\,
            I => \N__29767\
        );

    \I__7025\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29763\
        );

    \I__7024\ : Span4Mux_v
    port map (
            O => \N__29822\,
            I => \N__29760\
        );

    \I__7023\ : Span4Mux_v
    port map (
            O => \N__29811\,
            I => \N__29751\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__29808\,
            I => \N__29751\
        );

    \I__7021\ : Span4Mux_v
    port map (
            O => \N__29803\,
            I => \N__29751\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__29800\,
            I => \N__29751\
        );

    \I__7019\ : Span4Mux_h
    port map (
            O => \N__29797\,
            I => \N__29740\
        );

    \I__7018\ : Span4Mux_v
    port map (
            O => \N__29786\,
            I => \N__29740\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__29783\,
            I => \N__29740\
        );

    \I__7016\ : Span4Mux_v
    port map (
            O => \N__29776\,
            I => \N__29740\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__29773\,
            I => \N__29740\
        );

    \I__7014\ : Span12Mux_s8_h
    port map (
            O => \N__29770\,
            I => \N__29737\
        );

    \I__7013\ : Span4Mux_h
    port map (
            O => \N__29767\,
            I => \N__29734\
        );

    \I__7012\ : SRMux
    port map (
            O => \N__29766\,
            I => \N__29731\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__29763\,
            I => \N__29728\
        );

    \I__7010\ : Span4Mux_v
    port map (
            O => \N__29760\,
            I => \N__29725\
        );

    \I__7009\ : Span4Mux_v
    port map (
            O => \N__29751\,
            I => \N__29720\
        );

    \I__7008\ : Span4Mux_v
    port map (
            O => \N__29740\,
            I => \N__29720\
        );

    \I__7007\ : Span12Mux_h
    port map (
            O => \N__29737\,
            I => \N__29717\
        );

    \I__7006\ : Span4Mux_h
    port map (
            O => \N__29734\,
            I => \N__29714\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__29731\,
            I => \N__29711\
        );

    \I__7004\ : Span12Mux_v
    port map (
            O => \N__29728\,
            I => \N__29704\
        );

    \I__7003\ : Sp12to4
    port map (
            O => \N__29725\,
            I => \N__29704\
        );

    \I__7002\ : Sp12to4
    port map (
            O => \N__29720\,
            I => \N__29704\
        );

    \I__7001\ : Odrv12
    port map (
            O => \N__29717\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__29714\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6999\ : Odrv12
    port map (
            O => \N__29711\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6998\ : Odrv12
    port map (
            O => \N__29704\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6997\ : InMux
    port map (
            O => \N__29695\,
            I => \M_this_data_count_q_cry_13\
        );

    \I__6996\ : InMux
    port map (
            O => \N__29692\,
            I => \M_this_data_count_q_cry_14\
        );

    \I__6995\ : InMux
    port map (
            O => \N__29689\,
            I => \N__29686\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__29686\,
            I => \N__29683\
        );

    \I__6993\ : Span12Mux_v
    port map (
            O => \N__29683\,
            I => \N__29680\
        );

    \I__6992\ : Span12Mux_v
    port map (
            O => \N__29680\,
            I => \N__29677\
        );

    \I__6991\ : Odrv12
    port map (
            O => \N__29677\,
            I => \M_this_map_ram_read_data_6\
        );

    \I__6990\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29669\
        );

    \I__6989\ : CascadeMux
    port map (
            O => \N__29673\,
            I => \N__29666\
        );

    \I__6988\ : CascadeMux
    port map (
            O => \N__29672\,
            I => \N__29663\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__29669\,
            I => \N__29660\
        );

    \I__6986\ : InMux
    port map (
            O => \N__29666\,
            I => \N__29657\
        );

    \I__6985\ : InMux
    port map (
            O => \N__29663\,
            I => \N__29654\
        );

    \I__6984\ : Span4Mux_h
    port map (
            O => \N__29660\,
            I => \N__29651\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__29657\,
            I => \N__29646\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__29654\,
            I => \N__29646\
        );

    \I__6981\ : Span4Mux_h
    port map (
            O => \N__29651\,
            I => \N__29640\
        );

    \I__6980\ : Span4Mux_v
    port map (
            O => \N__29646\,
            I => \N__29640\
        );

    \I__6979\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29637\
        );

    \I__6978\ : Span4Mux_h
    port map (
            O => \N__29640\,
            I => \N__29634\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__29637\,
            I => \N__29631\
        );

    \I__6976\ : Span4Mux_h
    port map (
            O => \N__29634\,
            I => \N__29628\
        );

    \I__6975\ : Span12Mux_h
    port map (
            O => \N__29631\,
            I => \N__29625\
        );

    \I__6974\ : Odrv4
    port map (
            O => \N__29628\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__6973\ : Odrv12
    port map (
            O => \N__29625\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__6972\ : InMux
    port map (
            O => \N__29620\,
            I => \N__29613\
        );

    \I__6971\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29610\
        );

    \I__6970\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29607\
        );

    \I__6969\ : InMux
    port map (
            O => \N__29617\,
            I => \N__29603\
        );

    \I__6968\ : InMux
    port map (
            O => \N__29616\,
            I => \N__29600\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__29613\,
            I => \N__29597\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__29610\,
            I => \N__29592\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__29607\,
            I => \N__29589\
        );

    \I__6964\ : CascadeMux
    port map (
            O => \N__29606\,
            I => \N__29586\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__29603\,
            I => \N__29581\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__29600\,
            I => \N__29581\
        );

    \I__6961\ : Span4Mux_v
    port map (
            O => \N__29597\,
            I => \N__29578\
        );

    \I__6960\ : InMux
    port map (
            O => \N__29596\,
            I => \N__29575\
        );

    \I__6959\ : InMux
    port map (
            O => \N__29595\,
            I => \N__29572\
        );

    \I__6958\ : Span4Mux_h
    port map (
            O => \N__29592\,
            I => \N__29567\
        );

    \I__6957\ : Span4Mux_h
    port map (
            O => \N__29589\,
            I => \N__29567\
        );

    \I__6956\ : InMux
    port map (
            O => \N__29586\,
            I => \N__29564\
        );

    \I__6955\ : Span4Mux_h
    port map (
            O => \N__29581\,
            I => \N__29561\
        );

    \I__6954\ : Odrv4
    port map (
            O => \N__29578\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__29575\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__29572\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6951\ : Odrv4
    port map (
            O => \N__29567\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__29564\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6949\ : Odrv4
    port map (
            O => \N__29561\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6948\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29545\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__29545\,
            I => \M_this_data_count_q_s_2\
        );

    \I__6946\ : InMux
    port map (
            O => \N__29542\,
            I => \M_this_data_count_q_cry_1\
        );

    \I__6945\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29534\
        );

    \I__6944\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29531\
        );

    \I__6943\ : InMux
    port map (
            O => \N__29537\,
            I => \N__29528\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__29534\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__29531\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__29528\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__6939\ : CascadeMux
    port map (
            O => \N__29521\,
            I => \N__29518\
        );

    \I__6938\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29515\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__29515\,
            I => \M_this_data_count_q_s_3\
        );

    \I__6936\ : InMux
    port map (
            O => \N__29512\,
            I => \M_this_data_count_q_cry_2\
        );

    \I__6935\ : CascadeMux
    port map (
            O => \N__29509\,
            I => \N__29505\
        );

    \I__6934\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29501\
        );

    \I__6933\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29498\
        );

    \I__6932\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29495\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__29501\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__29498\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__29495\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__6928\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29485\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__29485\,
            I => \M_this_data_count_q_s_4\
        );

    \I__6926\ : InMux
    port map (
            O => \N__29482\,
            I => \M_this_data_count_q_cry_3\
        );

    \I__6925\ : InMux
    port map (
            O => \N__29479\,
            I => \N__29474\
        );

    \I__6924\ : InMux
    port map (
            O => \N__29478\,
            I => \N__29469\
        );

    \I__6923\ : InMux
    port map (
            O => \N__29477\,
            I => \N__29469\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__29474\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__29469\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__29464\,
            I => \N__29461\
        );

    \I__6919\ : InMux
    port map (
            O => \N__29461\,
            I => \N__29458\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__29458\,
            I => \M_this_data_count_q_s_5\
        );

    \I__6917\ : InMux
    port map (
            O => \N__29455\,
            I => \M_this_data_count_q_cry_4\
        );

    \I__6916\ : CascadeMux
    port map (
            O => \N__29452\,
            I => \N__29449\
        );

    \I__6915\ : InMux
    port map (
            O => \N__29449\,
            I => \N__29444\
        );

    \I__6914\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29439\
        );

    \I__6913\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29439\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__29444\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__29439\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__6910\ : CascadeMux
    port map (
            O => \N__29434\,
            I => \N__29431\
        );

    \I__6909\ : InMux
    port map (
            O => \N__29431\,
            I => \N__29428\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__29428\,
            I => \M_this_data_count_q_s_6\
        );

    \I__6907\ : InMux
    port map (
            O => \N__29425\,
            I => \M_this_data_count_q_cry_5\
        );

    \I__6906\ : InMux
    port map (
            O => \N__29422\,
            I => \M_this_data_count_q_cry_6\
        );

    \I__6905\ : InMux
    port map (
            O => \N__29419\,
            I => \bfn_23_18_0_\
        );

    \I__6904\ : InMux
    port map (
            O => \N__29416\,
            I => \M_this_data_count_q_cry_8\
        );

    \I__6903\ : InMux
    port map (
            O => \N__29413\,
            I => \M_this_data_count_q_cry_9\
        );

    \I__6902\ : InMux
    port map (
            O => \N__29410\,
            I => \N__29407\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__29407\,
            I => \N_509\
        );

    \I__6900\ : CascadeMux
    port map (
            O => \N__29404\,
            I => \N_510_cascade_\
        );

    \I__6899\ : InMux
    port map (
            O => \N__29401\,
            I => \N__29398\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__29398\,
            I => \N_511\
        );

    \I__6897\ : InMux
    port map (
            O => \N__29395\,
            I => \N__29392\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__29392\,
            I => \N_512\
        );

    \I__6895\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29386\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__29386\,
            I => \N__29383\
        );

    \I__6893\ : Span4Mux_v
    port map (
            O => \N__29383\,
            I => \N__29379\
        );

    \I__6892\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29374\
        );

    \I__6891\ : Span4Mux_v
    port map (
            O => \N__29379\,
            I => \N__29371\
        );

    \I__6890\ : InMux
    port map (
            O => \N__29378\,
            I => \N__29368\
        );

    \I__6889\ : InMux
    port map (
            O => \N__29377\,
            I => \N__29365\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__29374\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6887\ : Odrv4
    port map (
            O => \N__29371\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__29368\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__29365\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6884\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29351\
        );

    \I__6883\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29348\
        );

    \I__6882\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29345\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__29351\,
            I => \N__29342\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__29348\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__29345\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__6878\ : Odrv4
    port map (
            O => \N__29342\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__6877\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29332\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__29332\,
            I => \M_this_data_count_q_s_1\
        );

    \I__6875\ : InMux
    port map (
            O => \N__29329\,
            I => \M_this_data_count_q_cry_0\
        );

    \I__6874\ : CascadeMux
    port map (
            O => \N__29326\,
            I => \N__29322\
        );

    \I__6873\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29318\
        );

    \I__6872\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29315\
        );

    \I__6871\ : InMux
    port map (
            O => \N__29321\,
            I => \N__29312\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__29318\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__29315\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__29312\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__6867\ : IoInMux
    port map (
            O => \N__29305\,
            I => \N__29302\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__29302\,
            I => \N__29299\
        );

    \I__6865\ : Span4Mux_s0_v
    port map (
            O => \N__29299\,
            I => \N__29296\
        );

    \I__6864\ : Sp12to4
    port map (
            O => \N__29296\,
            I => \N__29292\
        );

    \I__6863\ : InMux
    port map (
            O => \N__29295\,
            I => \N__29287\
        );

    \I__6862\ : Span12Mux_s10_h
    port map (
            O => \N__29292\,
            I => \N__29284\
        );

    \I__6861\ : InMux
    port map (
            O => \N__29291\,
            I => \N__29279\
        );

    \I__6860\ : InMux
    port map (
            O => \N__29290\,
            I => \N__29279\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__29287\,
            I => \N__29276\
        );

    \I__6858\ : Odrv12
    port map (
            O => \N__29284\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__29279\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__6856\ : Odrv4
    port map (
            O => \N__29276\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__6855\ : InMux
    port map (
            O => \N__29269\,
            I => \N__29266\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__29266\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_11\
        );

    \I__6853\ : CascadeMux
    port map (
            O => \N__29263\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_3_cascade_\
        );

    \I__6852\ : InMux
    port map (
            O => \N__29260\,
            I => \N__29257\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__29257\,
            I => \N__29254\
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__29254\,
            I => \un1_M_this_external_address_q_cry_2_c_RNIKMIBZ0\
        );

    \I__6849\ : IoInMux
    port map (
            O => \N__29251\,
            I => \N__29248\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__29248\,
            I => \N__29245\
        );

    \I__6847\ : IoSpan4Mux
    port map (
            O => \N__29245\,
            I => \N__29242\
        );

    \I__6846\ : Span4Mux_s1_h
    port map (
            O => \N__29242\,
            I => \N__29239\
        );

    \I__6845\ : Span4Mux_v
    port map (
            O => \N__29239\,
            I => \N__29234\
        );

    \I__6844\ : CascadeMux
    port map (
            O => \N__29238\,
            I => \N__29231\
        );

    \I__6843\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29227\
        );

    \I__6842\ : Sp12to4
    port map (
            O => \N__29234\,
            I => \N__29224\
        );

    \I__6841\ : InMux
    port map (
            O => \N__29231\,
            I => \N__29219\
        );

    \I__6840\ : InMux
    port map (
            O => \N__29230\,
            I => \N__29219\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__29227\,
            I => \N__29216\
        );

    \I__6838\ : Odrv12
    port map (
            O => \N__29224\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__29219\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__6836\ : Odrv4
    port map (
            O => \N__29216\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__6835\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29206\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__29206\,
            I => \this_vga_signals.M_this_external_address_d_8_mZ0Z_3\
        );

    \I__6833\ : InMux
    port map (
            O => \N__29203\,
            I => \N__29200\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__29200\,
            I => \N__29197\
        );

    \I__6831\ : Span12Mux_v
    port map (
            O => \N__29197\,
            I => \N__29194\
        );

    \I__6830\ : Odrv12
    port map (
            O => \N__29194\,
            I => \M_this_data_count_q_s_0\
        );

    \I__6829\ : InMux
    port map (
            O => \N__29191\,
            I => \N__29182\
        );

    \I__6828\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29182\
        );

    \I__6827\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29177\
        );

    \I__6826\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29174\
        );

    \I__6825\ : InMux
    port map (
            O => \N__29187\,
            I => \N__29171\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__29182\,
            I => \N__29168\
        );

    \I__6823\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29165\
        );

    \I__6822\ : InMux
    port map (
            O => \N__29180\,
            I => \N__29156\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__29177\,
            I => \N__29153\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__29174\,
            I => \N__29146\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__29171\,
            I => \N__29146\
        );

    \I__6818\ : Span4Mux_h
    port map (
            O => \N__29168\,
            I => \N__29146\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__29165\,
            I => \N__29143\
        );

    \I__6816\ : InMux
    port map (
            O => \N__29164\,
            I => \N__29140\
        );

    \I__6815\ : InMux
    port map (
            O => \N__29163\,
            I => \N__29137\
        );

    \I__6814\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29134\
        );

    \I__6813\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29131\
        );

    \I__6812\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29128\
        );

    \I__6811\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29125\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__29156\,
            I => \N__29122\
        );

    \I__6809\ : Span4Mux_h
    port map (
            O => \N__29153\,
            I => \N__29119\
        );

    \I__6808\ : Span4Mux_v
    port map (
            O => \N__29146\,
            I => \N__29114\
        );

    \I__6807\ : Span4Mux_h
    port map (
            O => \N__29143\,
            I => \N__29114\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__29140\,
            I => \N__29111\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__29137\,
            I => \N__29102\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__29134\,
            I => \N__29102\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__29131\,
            I => \N__29102\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__29128\,
            I => \N__29102\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__29125\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6800\ : Odrv4
    port map (
            O => \N__29122\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6799\ : Odrv4
    port map (
            O => \N__29119\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__29114\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6797\ : Odrv12
    port map (
            O => \N__29111\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__29102\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6795\ : CascadeMux
    port map (
            O => \N__29089\,
            I => \this_vga_signals.N_292_cascade_\
        );

    \I__6794\ : InMux
    port map (
            O => \N__29086\,
            I => \N__29083\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__29083\,
            I => \N__29079\
        );

    \I__6792\ : InMux
    port map (
            O => \N__29082\,
            I => \N__29076\
        );

    \I__6791\ : Span4Mux_h
    port map (
            O => \N__29079\,
            I => \N__29073\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__29076\,
            I => \N__29070\
        );

    \I__6789\ : Odrv4
    port map (
            O => \N__29073\,
            I => \this_vga_signals.M_this_external_address_d_2_sqmuxaZ0\
        );

    \I__6788\ : Odrv4
    port map (
            O => \N__29070\,
            I => \this_vga_signals.M_this_external_address_d_2_sqmuxaZ0\
        );

    \I__6787\ : InMux
    port map (
            O => \N__29065\,
            I => \N__29062\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__29062\,
            I => \M_this_state_d88_9\
        );

    \I__6785\ : CascadeMux
    port map (
            O => \N__29059\,
            I => \N__29056\
        );

    \I__6784\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29053\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__29053\,
            I => \N__29050\
        );

    \I__6782\ : Odrv4
    port map (
            O => \N__29050\,
            I => \N_506\
        );

    \I__6781\ : InMux
    port map (
            O => \N__29047\,
            I => \N__29044\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__29044\,
            I => \un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0\
        );

    \I__6779\ : CascadeMux
    port map (
            O => \N__29041\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_8_cascade_\
        );

    \I__6778\ : IoInMux
    port map (
            O => \N__29038\,
            I => \N__29035\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__29035\,
            I => \N__29032\
        );

    \I__6776\ : Span4Mux_s1_v
    port map (
            O => \N__29032\,
            I => \N__29029\
        );

    \I__6775\ : Sp12to4
    port map (
            O => \N__29029\,
            I => \N__29025\
        );

    \I__6774\ : CascadeMux
    port map (
            O => \N__29028\,
            I => \N__29022\
        );

    \I__6773\ : Span12Mux_h
    port map (
            O => \N__29025\,
            I => \N__29017\
        );

    \I__6772\ : InMux
    port map (
            O => \N__29022\,
            I => \N__29012\
        );

    \I__6771\ : InMux
    port map (
            O => \N__29021\,
            I => \N__29012\
        );

    \I__6770\ : InMux
    port map (
            O => \N__29020\,
            I => \N__29009\
        );

    \I__6769\ : Odrv12
    port map (
            O => \N__29017\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__29012\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__29009\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__6766\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__28999\,
            I => \this_vga_signals.M_this_external_address_d_5_mZ0Z_8\
        );

    \I__6764\ : CascadeMux
    port map (
            O => \N__28996\,
            I => \this_vga_signals.M_this_external_address_d_8_mZ0Z_0_cascade_\
        );

    \I__6763\ : InMux
    port map (
            O => \N__28993\,
            I => \N__28990\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__28990\,
            I => \N__28987\
        );

    \I__6761\ : Odrv12
    port map (
            O => \N__28987\,
            I => \M_this_external_address_q_RNIE44V9Z0Z_0\
        );

    \I__6760\ : IoInMux
    port map (
            O => \N__28984\,
            I => \N__28981\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__28981\,
            I => \N__28978\
        );

    \I__6758\ : IoSpan4Mux
    port map (
            O => \N__28978\,
            I => \N__28975\
        );

    \I__6757\ : Span4Mux_s2_v
    port map (
            O => \N__28975\,
            I => \N__28972\
        );

    \I__6756\ : Span4Mux_v
    port map (
            O => \N__28972\,
            I => \N__28968\
        );

    \I__6755\ : InMux
    port map (
            O => \N__28971\,
            I => \N__28963\
        );

    \I__6754\ : Span4Mux_v
    port map (
            O => \N__28968\,
            I => \N__28960\
        );

    \I__6753\ : InMux
    port map (
            O => \N__28967\,
            I => \N__28955\
        );

    \I__6752\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28955\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__28963\,
            I => \N__28952\
        );

    \I__6750\ : Odrv4
    port map (
            O => \N__28960\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__28955\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__6748\ : Odrv4
    port map (
            O => \N__28952\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__6747\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28942\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__28942\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_0\
        );

    \I__6745\ : CascadeMux
    port map (
            O => \N__28939\,
            I => \N__28936\
        );

    \I__6744\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28933\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__28933\,
            I => \N__28930\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__28930\,
            I => \this_vga_signals.M_this_external_address_d_5_mZ0Z_9\
        );

    \I__6741\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28924\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__28924\,
            I => \un1_M_this_external_address_q_cry_8_c_RNI09PBZ0\
        );

    \I__6739\ : CascadeMux
    port map (
            O => \N__28921\,
            I => \this_vga_signals.M_this_external_address_d_5_mZ0Z_11_cascade_\
        );

    \I__6738\ : InMux
    port map (
            O => \N__28918\,
            I => \N__28915\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__28915\,
            I => \N__28912\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__28912\,
            I => \un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0\
        );

    \I__6735\ : InMux
    port map (
            O => \N__28909\,
            I => \bfn_22_21_0_\
        );

    \I__6734\ : InMux
    port map (
            O => \N__28906\,
            I => \un1_M_this_external_address_q_cry_8\
        );

    \I__6733\ : InMux
    port map (
            O => \N__28903\,
            I => \un1_M_this_external_address_q_cry_9\
        );

    \I__6732\ : InMux
    port map (
            O => \N__28900\,
            I => \un1_M_this_external_address_q_cry_10\
        );

    \I__6731\ : InMux
    port map (
            O => \N__28897\,
            I => \un1_M_this_external_address_q_cry_11\
        );

    \I__6730\ : IoInMux
    port map (
            O => \N__28894\,
            I => \N__28891\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__28891\,
            I => \N__28888\
        );

    \I__6728\ : Span4Mux_s2_h
    port map (
            O => \N__28888\,
            I => \N__28885\
        );

    \I__6727\ : Span4Mux_h
    port map (
            O => \N__28885\,
            I => \N__28881\
        );

    \I__6726\ : InMux
    port map (
            O => \N__28884\,
            I => \N__28878\
        );

    \I__6725\ : Span4Mux_h
    port map (
            O => \N__28881\,
            I => \N__28871\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__28878\,
            I => \N__28871\
        );

    \I__6723\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28866\
        );

    \I__6722\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28866\
        );

    \I__6721\ : Odrv4
    port map (
            O => \N__28871\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__28866\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__6719\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28858\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28855\
        );

    \I__6717\ : Odrv4
    port map (
            O => \N__28855\,
            I => \un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0\
        );

    \I__6716\ : InMux
    port map (
            O => \N__28852\,
            I => \un1_M_this_external_address_q_cry_12\
        );

    \I__6715\ : IoInMux
    port map (
            O => \N__28849\,
            I => \N__28846\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__28846\,
            I => \N__28843\
        );

    \I__6713\ : Span4Mux_s3_h
    port map (
            O => \N__28843\,
            I => \N__28839\
        );

    \I__6712\ : InMux
    port map (
            O => \N__28842\,
            I => \N__28835\
        );

    \I__6711\ : Span4Mux_h
    port map (
            O => \N__28839\,
            I => \N__28832\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__28838\,
            I => \N__28829\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__28835\,
            I => \N__28826\
        );

    \I__6708\ : Span4Mux_h
    port map (
            O => \N__28832\,
            I => \N__28822\
        );

    \I__6707\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28819\
        );

    \I__6706\ : Span4Mux_h
    port map (
            O => \N__28826\,
            I => \N__28816\
        );

    \I__6705\ : InMux
    port map (
            O => \N__28825\,
            I => \N__28813\
        );

    \I__6704\ : Odrv4
    port map (
            O => \N__28822\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__28819\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__6702\ : Odrv4
    port map (
            O => \N__28816\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__28813\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__6700\ : InMux
    port map (
            O => \N__28804\,
            I => \N__28801\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__28801\,
            I => \N__28798\
        );

    \I__6698\ : Span4Mux_h
    port map (
            O => \N__28798\,
            I => \N__28795\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__28795\,
            I => \un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0\
        );

    \I__6696\ : InMux
    port map (
            O => \N__28792\,
            I => \un1_M_this_external_address_q_cry_13\
        );

    \I__6695\ : InMux
    port map (
            O => \N__28789\,
            I => \un1_M_this_external_address_q_cry_14\
        );

    \I__6694\ : CascadeMux
    port map (
            O => \N__28786\,
            I => \N__28781\
        );

    \I__6693\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28778\
        );

    \I__6692\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28775\
        );

    \I__6691\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28772\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__28778\,
            I => \un1_M_this_state_q_16_0\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__28775\,
            I => \un1_M_this_state_q_16_0\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__28772\,
            I => \un1_M_this_state_q_16_0\
        );

    \I__6687\ : InMux
    port map (
            O => \N__28765\,
            I => \un1_M_this_external_address_q_cry_0\
        );

    \I__6686\ : InMux
    port map (
            O => \N__28762\,
            I => \un1_M_this_external_address_q_cry_1\
        );

    \I__6685\ : InMux
    port map (
            O => \N__28759\,
            I => \un1_M_this_external_address_q_cry_2\
        );

    \I__6684\ : InMux
    port map (
            O => \N__28756\,
            I => \un1_M_this_external_address_q_cry_3\
        );

    \I__6683\ : IoInMux
    port map (
            O => \N__28753\,
            I => \N__28750\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__28750\,
            I => \N__28745\
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__28749\,
            I => \N__28741\
        );

    \I__6680\ : CascadeMux
    port map (
            O => \N__28748\,
            I => \N__28738\
        );

    \I__6679\ : Span12Mux_s4_h
    port map (
            O => \N__28745\,
            I => \N__28735\
        );

    \I__6678\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28732\
        );

    \I__6677\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28729\
        );

    \I__6676\ : InMux
    port map (
            O => \N__28738\,
            I => \N__28726\
        );

    \I__6675\ : Odrv12
    port map (
            O => \N__28735\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__28732\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__28729\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__28726\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__6671\ : InMux
    port map (
            O => \N__28717\,
            I => \N__28714\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__28714\,
            I => \un1_M_this_external_address_q_cry_4_c_RNIOSKBZ0\
        );

    \I__6669\ : InMux
    port map (
            O => \N__28711\,
            I => \un1_M_this_external_address_q_cry_4\
        );

    \I__6668\ : IoInMux
    port map (
            O => \N__28708\,
            I => \N__28705\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28702\
        );

    \I__6666\ : Span4Mux_s2_h
    port map (
            O => \N__28702\,
            I => \N__28699\
        );

    \I__6665\ : Span4Mux_v
    port map (
            O => \N__28699\,
            I => \N__28695\
        );

    \I__6664\ : InMux
    port map (
            O => \N__28698\,
            I => \N__28691\
        );

    \I__6663\ : Sp12to4
    port map (
            O => \N__28695\,
            I => \N__28687\
        );

    \I__6662\ : InMux
    port map (
            O => \N__28694\,
            I => \N__28684\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__28691\,
            I => \N__28681\
        );

    \I__6660\ : InMux
    port map (
            O => \N__28690\,
            I => \N__28678\
        );

    \I__6659\ : Odrv12
    port map (
            O => \N__28687\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__28684\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__6657\ : Odrv12
    port map (
            O => \N__28681\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__28678\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__6655\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28666\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__28666\,
            I => \un1_M_this_external_address_q_cry_5_c_RNIQVLBZ0\
        );

    \I__6653\ : InMux
    port map (
            O => \N__28663\,
            I => \un1_M_this_external_address_q_cry_5\
        );

    \I__6652\ : InMux
    port map (
            O => \N__28660\,
            I => \un1_M_this_external_address_q_cry_6\
        );

    \I__6651\ : CascadeMux
    port map (
            O => \N__28657\,
            I => \N_508_cascade_\
        );

    \I__6650\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28651\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28648\
        );

    \I__6648\ : Odrv4
    port map (
            O => \N__28648\,
            I => \M_this_state_d88_11\
        );

    \I__6647\ : CascadeMux
    port map (
            O => \N__28645\,
            I => \M_this_state_d88_11_cascade_\
        );

    \I__6646\ : InMux
    port map (
            O => \N__28642\,
            I => \N__28639\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__28639\,
            I => \N__28636\
        );

    \I__6644\ : Odrv12
    port map (
            O => \N__28636\,
            I => \M_this_state_d88_12\
        );

    \I__6643\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28630\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__28630\,
            I => \N__28627\
        );

    \I__6641\ : Odrv4
    port map (
            O => \N__28627\,
            I => \N_436\
        );

    \I__6640\ : InMux
    port map (
            O => \N__28624\,
            I => \N__28621\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__28621\,
            I => \N__28618\
        );

    \I__6638\ : Span4Mux_v
    port map (
            O => \N__28618\,
            I => \N__28615\
        );

    \I__6637\ : Span4Mux_h
    port map (
            O => \N__28615\,
            I => \N__28612\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__28612\,
            I => \N_465\
        );

    \I__6635\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28606\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__28606\,
            I => \N__28603\
        );

    \I__6633\ : Span4Mux_h
    port map (
            O => \N__28603\,
            I => \N__28600\
        );

    \I__6632\ : Odrv4
    port map (
            O => \N__28600\,
            I => \N_435\
        );

    \I__6631\ : CascadeMux
    port map (
            O => \N__28597\,
            I => \M_this_state_qsr_0_cascade_\
        );

    \I__6630\ : InMux
    port map (
            O => \N__28594\,
            I => \N__28591\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__28591\,
            I => \N__28588\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__28588\,
            I => \N_466\
        );

    \I__6627\ : IoInMux
    port map (
            O => \N__28585\,
            I => \N__28582\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__28582\,
            I => \N__28579\
        );

    \I__6625\ : Span4Mux_s2_h
    port map (
            O => \N__28579\,
            I => \N__28575\
        );

    \I__6624\ : CascadeMux
    port map (
            O => \N__28578\,
            I => \N__28571\
        );

    \I__6623\ : Span4Mux_h
    port map (
            O => \N__28575\,
            I => \N__28568\
        );

    \I__6622\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28565\
        );

    \I__6621\ : InMux
    port map (
            O => \N__28571\,
            I => \N__28562\
        );

    \I__6620\ : Sp12to4
    port map (
            O => \N__28568\,
            I => \N__28556\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__28565\,
            I => \N__28551\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__28562\,
            I => \N__28551\
        );

    \I__6617\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28544\
        );

    \I__6616\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28544\
        );

    \I__6615\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28544\
        );

    \I__6614\ : Span12Mux_v
    port map (
            O => \N__28556\,
            I => \N__28541\
        );

    \I__6613\ : Span4Mux_h
    port map (
            O => \N__28551\,
            I => \N__28538\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__28544\,
            I => \N__28535\
        );

    \I__6611\ : Odrv12
    port map (
            O => \N__28541\,
            I => led_c_1
        );

    \I__6610\ : Odrv4
    port map (
            O => \N__28538\,
            I => led_c_1
        );

    \I__6609\ : Odrv4
    port map (
            O => \N__28535\,
            I => led_c_1
        );

    \I__6608\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28525\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__28525\,
            I => \N__28520\
        );

    \I__6606\ : InMux
    port map (
            O => \N__28524\,
            I => \N__28517\
        );

    \I__6605\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28514\
        );

    \I__6604\ : Span4Mux_v
    port map (
            O => \N__28520\,
            I => \N__28509\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__28517\,
            I => \N__28509\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__28514\,
            I => \N__28506\
        );

    \I__6601\ : Span4Mux_h
    port map (
            O => \N__28509\,
            I => \N__28501\
        );

    \I__6600\ : Span4Mux_h
    port map (
            O => \N__28506\,
            I => \N__28498\
        );

    \I__6599\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28495\
        );

    \I__6598\ : InMux
    port map (
            O => \N__28504\,
            I => \N__28492\
        );

    \I__6597\ : Odrv4
    port map (
            O => \N__28501\,
            I => \M_this_state_d88\
        );

    \I__6596\ : Odrv4
    port map (
            O => \N__28498\,
            I => \M_this_state_d88\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__28495\,
            I => \M_this_state_d88\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__28492\,
            I => \M_this_state_d88\
        );

    \I__6593\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28478\
        );

    \I__6592\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28475\
        );

    \I__6591\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28472\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__28478\,
            I => \N__28462\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__28475\,
            I => \N__28457\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__28472\,
            I => \N__28457\
        );

    \I__6587\ : InMux
    port map (
            O => \N__28471\,
            I => \N__28452\
        );

    \I__6586\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28452\
        );

    \I__6585\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28445\
        );

    \I__6584\ : InMux
    port map (
            O => \N__28468\,
            I => \N__28445\
        );

    \I__6583\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28445\
        );

    \I__6582\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28440\
        );

    \I__6581\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28440\
        );

    \I__6580\ : Span4Mux_h
    port map (
            O => \N__28462\,
            I => \N__28435\
        );

    \I__6579\ : Span4Mux_h
    port map (
            O => \N__28457\,
            I => \N__28435\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__28452\,
            I => \N__28432\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__28445\,
            I => \N__28429\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__28440\,
            I => \N__28426\
        );

    \I__6575\ : Span4Mux_v
    port map (
            O => \N__28435\,
            I => \N__28423\
        );

    \I__6574\ : Span4Mux_h
    port map (
            O => \N__28432\,
            I => \N__28420\
        );

    \I__6573\ : Span4Mux_v
    port map (
            O => \N__28429\,
            I => \N__28417\
        );

    \I__6572\ : Span12Mux_h
    port map (
            O => \N__28426\,
            I => \N__28414\
        );

    \I__6571\ : Span4Mux_v
    port map (
            O => \N__28423\,
            I => \N__28411\
        );

    \I__6570\ : Span4Mux_v
    port map (
            O => \N__28420\,
            I => \N__28408\
        );

    \I__6569\ : Span4Mux_v
    port map (
            O => \N__28417\,
            I => \N__28405\
        );

    \I__6568\ : Span12Mux_v
    port map (
            O => \N__28414\,
            I => \N__28402\
        );

    \I__6567\ : Span4Mux_v
    port map (
            O => \N__28411\,
            I => \N__28399\
        );

    \I__6566\ : Span4Mux_v
    port map (
            O => \N__28408\,
            I => \N__28396\
        );

    \I__6565\ : IoSpan4Mux
    port map (
            O => \N__28405\,
            I => \N__28393\
        );

    \I__6564\ : Odrv12
    port map (
            O => \N__28402\,
            I => rst_n_c
        );

    \I__6563\ : Odrv4
    port map (
            O => \N__28399\,
            I => rst_n_c
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__28396\,
            I => rst_n_c
        );

    \I__6561\ : Odrv4
    port map (
            O => \N__28393\,
            I => rst_n_c
        );

    \I__6560\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28381\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__28381\,
            I => \N__28378\
        );

    \I__6558\ : Span4Mux_h
    port map (
            O => \N__28378\,
            I => \N__28375\
        );

    \I__6557\ : Odrv4
    port map (
            O => \N__28375\,
            I => \this_reset_cond.M_stage_qZ0Z_7\
        );

    \I__6556\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28369\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__28369\,
            I => \this_reset_cond.M_stage_qZ0Z_8\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__28366\,
            I => \N__28363\
        );

    \I__6553\ : CascadeBuf
    port map (
            O => \N__28363\,
            I => \N__28360\
        );

    \I__6552\ : CascadeMux
    port map (
            O => \N__28360\,
            I => \N__28357\
        );

    \I__6551\ : CascadeBuf
    port map (
            O => \N__28357\,
            I => \N__28354\
        );

    \I__6550\ : CascadeMux
    port map (
            O => \N__28354\,
            I => \N__28351\
        );

    \I__6549\ : CascadeBuf
    port map (
            O => \N__28351\,
            I => \N__28348\
        );

    \I__6548\ : CascadeMux
    port map (
            O => \N__28348\,
            I => \N__28345\
        );

    \I__6547\ : CascadeBuf
    port map (
            O => \N__28345\,
            I => \N__28342\
        );

    \I__6546\ : CascadeMux
    port map (
            O => \N__28342\,
            I => \N__28339\
        );

    \I__6545\ : CascadeBuf
    port map (
            O => \N__28339\,
            I => \N__28336\
        );

    \I__6544\ : CascadeMux
    port map (
            O => \N__28336\,
            I => \N__28333\
        );

    \I__6543\ : CascadeBuf
    port map (
            O => \N__28333\,
            I => \N__28330\
        );

    \I__6542\ : CascadeMux
    port map (
            O => \N__28330\,
            I => \N__28327\
        );

    \I__6541\ : CascadeBuf
    port map (
            O => \N__28327\,
            I => \N__28324\
        );

    \I__6540\ : CascadeMux
    port map (
            O => \N__28324\,
            I => \N__28321\
        );

    \I__6539\ : CascadeBuf
    port map (
            O => \N__28321\,
            I => \N__28318\
        );

    \I__6538\ : CascadeMux
    port map (
            O => \N__28318\,
            I => \N__28315\
        );

    \I__6537\ : CascadeBuf
    port map (
            O => \N__28315\,
            I => \N__28312\
        );

    \I__6536\ : CascadeMux
    port map (
            O => \N__28312\,
            I => \N__28309\
        );

    \I__6535\ : CascadeBuf
    port map (
            O => \N__28309\,
            I => \N__28306\
        );

    \I__6534\ : CascadeMux
    port map (
            O => \N__28306\,
            I => \N__28303\
        );

    \I__6533\ : CascadeBuf
    port map (
            O => \N__28303\,
            I => \N__28300\
        );

    \I__6532\ : CascadeMux
    port map (
            O => \N__28300\,
            I => \N__28297\
        );

    \I__6531\ : CascadeBuf
    port map (
            O => \N__28297\,
            I => \N__28294\
        );

    \I__6530\ : CascadeMux
    port map (
            O => \N__28294\,
            I => \N__28291\
        );

    \I__6529\ : CascadeBuf
    port map (
            O => \N__28291\,
            I => \N__28288\
        );

    \I__6528\ : CascadeMux
    port map (
            O => \N__28288\,
            I => \N__28285\
        );

    \I__6527\ : CascadeBuf
    port map (
            O => \N__28285\,
            I => \N__28282\
        );

    \I__6526\ : CascadeMux
    port map (
            O => \N__28282\,
            I => \N__28279\
        );

    \I__6525\ : CascadeBuf
    port map (
            O => \N__28279\,
            I => \N__28276\
        );

    \I__6524\ : CascadeMux
    port map (
            O => \N__28276\,
            I => \N__28273\
        );

    \I__6523\ : InMux
    port map (
            O => \N__28273\,
            I => \N__28270\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__28270\,
            I => \N__28267\
        );

    \I__6521\ : Span4Mux_s1_v
    port map (
            O => \N__28267\,
            I => \N__28263\
        );

    \I__6520\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28259\
        );

    \I__6519\ : Sp12to4
    port map (
            O => \N__28263\,
            I => \N__28255\
        );

    \I__6518\ : InMux
    port map (
            O => \N__28262\,
            I => \N__28252\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__28259\,
            I => \N__28249\
        );

    \I__6516\ : InMux
    port map (
            O => \N__28258\,
            I => \N__28246\
        );

    \I__6515\ : Span12Mux_h
    port map (
            O => \N__28255\,
            I => \N__28243\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__28252\,
            I => \N__28238\
        );

    \I__6513\ : Span4Mux_h
    port map (
            O => \N__28249\,
            I => \N__28238\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__28246\,
            I => \N__28233\
        );

    \I__6511\ : Span12Mux_v
    port map (
            O => \N__28243\,
            I => \N__28233\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__28238\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__6509\ : Odrv12
    port map (
            O => \N__28233\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__6508\ : CascadeMux
    port map (
            O => \N__28228\,
            I => \N__28223\
        );

    \I__6507\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28217\
        );

    \I__6506\ : InMux
    port map (
            O => \N__28226\,
            I => \N__28214\
        );

    \I__6505\ : InMux
    port map (
            O => \N__28223\,
            I => \N__28208\
        );

    \I__6504\ : CascadeMux
    port map (
            O => \N__28222\,
            I => \N__28204\
        );

    \I__6503\ : InMux
    port map (
            O => \N__28221\,
            I => \N__28200\
        );

    \I__6502\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28195\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__28217\,
            I => \N__28190\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__28214\,
            I => \N__28190\
        );

    \I__6499\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28185\
        );

    \I__6498\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28185\
        );

    \I__6497\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28182\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__28208\,
            I => \N__28179\
        );

    \I__6495\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28176\
        );

    \I__6494\ : InMux
    port map (
            O => \N__28204\,
            I => \N__28171\
        );

    \I__6493\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28171\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__28200\,
            I => \N__28167\
        );

    \I__6491\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28164\
        );

    \I__6490\ : InMux
    port map (
            O => \N__28198\,
            I => \N__28157\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__28195\,
            I => \N__28150\
        );

    \I__6488\ : Span4Mux_v
    port map (
            O => \N__28190\,
            I => \N__28150\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__28185\,
            I => \N__28150\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__28182\,
            I => \N__28145\
        );

    \I__6485\ : Span4Mux_h
    port map (
            O => \N__28179\,
            I => \N__28145\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__28176\,
            I => \N__28140\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__28171\,
            I => \N__28140\
        );

    \I__6482\ : InMux
    port map (
            O => \N__28170\,
            I => \N__28137\
        );

    \I__6481\ : Span4Mux_v
    port map (
            O => \N__28167\,
            I => \N__28132\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__28164\,
            I => \N__28132\
        );

    \I__6479\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28127\
        );

    \I__6478\ : InMux
    port map (
            O => \N__28162\,
            I => \N__28127\
        );

    \I__6477\ : InMux
    port map (
            O => \N__28161\,
            I => \N__28124\
        );

    \I__6476\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28121\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__28157\,
            I => \N__28116\
        );

    \I__6474\ : Span4Mux_v
    port map (
            O => \N__28150\,
            I => \N__28116\
        );

    \I__6473\ : Sp12to4
    port map (
            O => \N__28145\,
            I => \N__28111\
        );

    \I__6472\ : Span12Mux_h
    port map (
            O => \N__28140\,
            I => \N__28111\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__28137\,
            I => \N__28104\
        );

    \I__6470\ : Span4Mux_h
    port map (
            O => \N__28132\,
            I => \N__28104\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__28127\,
            I => \N__28104\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__28124\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__28121\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__6466\ : Odrv4
    port map (
            O => \N__28116\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__6465\ : Odrv12
    port map (
            O => \N__28111\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__6464\ : Odrv4
    port map (
            O => \N__28104\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__6463\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28090\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__28090\,
            I => \N__28087\
        );

    \I__6461\ : Span4Mux_h
    port map (
            O => \N__28087\,
            I => \N__28084\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__28084\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__28081\,
            I => \M_this_state_d88_1_cascade_\
        );

    \I__6458\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28069\
        );

    \I__6457\ : InMux
    port map (
            O => \N__28077\,
            I => \N__28069\
        );

    \I__6456\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28064\
        );

    \I__6455\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28064\
        );

    \I__6454\ : InMux
    port map (
            O => \N__28074\,
            I => \N__28061\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__28069\,
            I => \N__28056\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__28064\,
            I => \N__28056\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__28061\,
            I => \N__28053\
        );

    \I__6450\ : Odrv4
    port map (
            O => \N__28056\,
            I => \this_vga_signals.N_390_0\
        );

    \I__6449\ : Odrv12
    port map (
            O => \N__28053\,
            I => \this_vga_signals.N_390_0\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__28048\,
            I => \M_this_state_d88_12_cascade_\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__28045\,
            I => \N_507_cascade_\
        );

    \I__6446\ : InMux
    port map (
            O => \N__28042\,
            I => \N__28037\
        );

    \I__6445\ : InMux
    port map (
            O => \N__28041\,
            I => \N__28032\
        );

    \I__6444\ : CascadeMux
    port map (
            O => \N__28040\,
            I => \N__28028\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__28037\,
            I => \N__28024\
        );

    \I__6442\ : InMux
    port map (
            O => \N__28036\,
            I => \N__28021\
        );

    \I__6441\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28018\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__28032\,
            I => \N__28014\
        );

    \I__6439\ : InMux
    port map (
            O => \N__28031\,
            I => \N__28011\
        );

    \I__6438\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28006\
        );

    \I__6437\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28006\
        );

    \I__6436\ : Span4Mux_h
    port map (
            O => \N__28024\,
            I => \N__28001\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__28021\,
            I => \N__28001\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__28018\,
            I => \N__27998\
        );

    \I__6433\ : InMux
    port map (
            O => \N__28017\,
            I => \N__27995\
        );

    \I__6432\ : Span4Mux_h
    port map (
            O => \N__28014\,
            I => \N__27991\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__28011\,
            I => \N__27982\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__28006\,
            I => \N__27982\
        );

    \I__6429\ : Span4Mux_v
    port map (
            O => \N__28001\,
            I => \N__27982\
        );

    \I__6428\ : Span4Mux_h
    port map (
            O => \N__27998\,
            I => \N__27982\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__27995\,
            I => \N__27979\
        );

    \I__6426\ : InMux
    port map (
            O => \N__27994\,
            I => \N__27976\
        );

    \I__6425\ : Span4Mux_h
    port map (
            O => \N__27991\,
            I => \N__27973\
        );

    \I__6424\ : Span4Mux_h
    port map (
            O => \N__27982\,
            I => \N__27970\
        );

    \I__6423\ : Odrv12
    port map (
            O => \N__27979\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__27976\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6421\ : Odrv4
    port map (
            O => \N__27973\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6420\ : Odrv4
    port map (
            O => \N__27970\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6419\ : InMux
    port map (
            O => \N__27961\,
            I => \N__27957\
        );

    \I__6418\ : InMux
    port map (
            O => \N__27960\,
            I => \N__27954\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__27957\,
            I => \N__27951\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__27954\,
            I => \this_vga_signals.N_293_1\
        );

    \I__6415\ : Odrv4
    port map (
            O => \N__27951\,
            I => \this_vga_signals.N_293_1\
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__27946\,
            I => \N__27941\
        );

    \I__6413\ : InMux
    port map (
            O => \N__27945\,
            I => \N__27937\
        );

    \I__6412\ : CascadeMux
    port map (
            O => \N__27944\,
            I => \N__27932\
        );

    \I__6411\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27929\
        );

    \I__6410\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27926\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27921\
        );

    \I__6408\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27916\
        );

    \I__6407\ : InMux
    port map (
            O => \N__27935\,
            I => \N__27916\
        );

    \I__6406\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27913\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27910\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27907\
        );

    \I__6403\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27902\
        );

    \I__6402\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27902\
        );

    \I__6401\ : Span4Mux_v
    port map (
            O => \N__27921\,
            I => \N__27899\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__27916\,
            I => \N__27894\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__27913\,
            I => \N__27894\
        );

    \I__6398\ : Span4Mux_v
    port map (
            O => \N__27910\,
            I => \N__27891\
        );

    \I__6397\ : Span4Mux_v
    port map (
            O => \N__27907\,
            I => \N__27888\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__27902\,
            I => \N__27885\
        );

    \I__6395\ : Span4Mux_h
    port map (
            O => \N__27899\,
            I => \N__27878\
        );

    \I__6394\ : Span4Mux_v
    port map (
            O => \N__27894\,
            I => \N__27878\
        );

    \I__6393\ : Span4Mux_h
    port map (
            O => \N__27891\,
            I => \N__27878\
        );

    \I__6392\ : Odrv4
    port map (
            O => \N__27888\,
            I => \M_this_state_qZ0Z_15\
        );

    \I__6391\ : Odrv12
    port map (
            O => \N__27885\,
            I => \M_this_state_qZ0Z_15\
        );

    \I__6390\ : Odrv4
    port map (
            O => \N__27878\,
            I => \M_this_state_qZ0Z_15\
        );

    \I__6389\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27868\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__27868\,
            I => \N__27865\
        );

    \I__6387\ : Span4Mux_h
    port map (
            O => \N__27865\,
            I => \N__27861\
        );

    \I__6386\ : InMux
    port map (
            O => \N__27864\,
            I => \N__27858\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__27861\,
            I => \N__27855\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27852\
        );

    \I__6383\ : Odrv4
    port map (
            O => \N__27855\,
            I => \this_vga_signals.M_this_map_ram_write_data_1_sqmuxa\
        );

    \I__6382\ : Odrv12
    port map (
            O => \N__27852\,
            I => \this_vga_signals.M_this_map_ram_write_data_1_sqmuxa\
        );

    \I__6381\ : CascadeMux
    port map (
            O => \N__27847\,
            I => \this_vga_signals.N_293_cascade_\
        );

    \I__6380\ : InMux
    port map (
            O => \N__27844\,
            I => \N__27841\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__27841\,
            I => \N__27838\
        );

    \I__6378\ : Span4Mux_v
    port map (
            O => \N__27838\,
            I => \N__27835\
        );

    \I__6377\ : Span4Mux_v
    port map (
            O => \N__27835\,
            I => \N__27832\
        );

    \I__6376\ : Span4Mux_h
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__6375\ : Odrv4
    port map (
            O => \N__27829\,
            I => \M_this_map_ram_read_data_7\
        );

    \I__6374\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27815\
        );

    \I__6373\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27812\
        );

    \I__6372\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27809\
        );

    \I__6371\ : InMux
    port map (
            O => \N__27823\,
            I => \N__27806\
        );

    \I__6370\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27795\
        );

    \I__6369\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27795\
        );

    \I__6368\ : InMux
    port map (
            O => \N__27820\,
            I => \N__27792\
        );

    \I__6367\ : InMux
    port map (
            O => \N__27819\,
            I => \N__27789\
        );

    \I__6366\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27786\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__27815\,
            I => \N__27781\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__27812\,
            I => \N__27781\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__27809\,
            I => \N__27776\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__27806\,
            I => \N__27776\
        );

    \I__6361\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27773\
        );

    \I__6360\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27770\
        );

    \I__6359\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27763\
        );

    \I__6358\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27763\
        );

    \I__6357\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27763\
        );

    \I__6356\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27759\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__27795\,
            I => \N__27754\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__27792\,
            I => \N__27754\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__27789\,
            I => \N__27747\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__27786\,
            I => \N__27747\
        );

    \I__6351\ : Span4Mux_v
    port map (
            O => \N__27781\,
            I => \N__27747\
        );

    \I__6350\ : Span4Mux_h
    port map (
            O => \N__27776\,
            I => \N__27744\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__27773\,
            I => \N__27737\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__27770\,
            I => \N__27737\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__27763\,
            I => \N__27737\
        );

    \I__6346\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27734\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__27759\,
            I => \N__27729\
        );

    \I__6344\ : Span4Mux_v
    port map (
            O => \N__27754\,
            I => \N__27729\
        );

    \I__6343\ : Span4Mux_h
    port map (
            O => \N__27747\,
            I => \N__27724\
        );

    \I__6342\ : Span4Mux_v
    port map (
            O => \N__27744\,
            I => \N__27724\
        );

    \I__6341\ : Span12Mux_v
    port map (
            O => \N__27737\,
            I => \N__27719\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__27734\,
            I => \N__27719\
        );

    \I__6339\ : Sp12to4
    port map (
            O => \N__27729\,
            I => \N__27716\
        );

    \I__6338\ : Span4Mux_h
    port map (
            O => \N__27724\,
            I => \N__27713\
        );

    \I__6337\ : Span12Mux_h
    port map (
            O => \N__27719\,
            I => \N__27710\
        );

    \I__6336\ : Odrv12
    port map (
            O => \N__27716\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__6335\ : Odrv4
    port map (
            O => \N__27713\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__6334\ : Odrv12
    port map (
            O => \N__27710\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__6333\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27700\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__27700\,
            I => \this_vga_signals.M_this_external_address_d_8_mZ0Z_5\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__27697\,
            I => \N__27694\
        );

    \I__6330\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27691\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__27691\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_5\
        );

    \I__6328\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27685\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__27685\,
            I => \N__27682\
        );

    \I__6326\ : Odrv12
    port map (
            O => \N__27682\,
            I => \this_vga_signals.M_this_external_address_q_mZ0Z_6\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__27679\,
            I => \this_vga_signals.M_this_external_address_d_8_mZ0Z_6_cascade_\
        );

    \I__6324\ : CascadeMux
    port map (
            O => \N__27676\,
            I => \N__27673\
        );

    \I__6323\ : CascadeBuf
    port map (
            O => \N__27673\,
            I => \N__27670\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__27670\,
            I => \N__27667\
        );

    \I__6321\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27664\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__27664\,
            I => \N__27661\
        );

    \I__6319\ : Span4Mux_s1_v
    port map (
            O => \N__27661\,
            I => \N__27658\
        );

    \I__6318\ : Span4Mux_h
    port map (
            O => \N__27658\,
            I => \N__27652\
        );

    \I__6317\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27649\
        );

    \I__6316\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27646\
        );

    \I__6315\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27643\
        );

    \I__6314\ : Span4Mux_v
    port map (
            O => \N__27652\,
            I => \N__27640\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__27649\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__27646\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__27643\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__27640\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__6309\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27628\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__27628\,
            I => \N__27618\
        );

    \I__6307\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27615\
        );

    \I__6306\ : InMux
    port map (
            O => \N__27626\,
            I => \N__27612\
        );

    \I__6305\ : CascadeMux
    port map (
            O => \N__27625\,
            I => \N__27608\
        );

    \I__6304\ : InMux
    port map (
            O => \N__27624\,
            I => \N__27604\
        );

    \I__6303\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27600\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__27622\,
            I => \N__27594\
        );

    \I__6301\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27591\
        );

    \I__6300\ : Span4Mux_v
    port map (
            O => \N__27618\,
            I => \N__27586\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__27615\,
            I => \N__27586\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__27612\,
            I => \N__27583\
        );

    \I__6297\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27578\
        );

    \I__6296\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27578\
        );

    \I__6295\ : CascadeMux
    port map (
            O => \N__27607\,
            I => \N__27575\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__27604\,
            I => \N__27572\
        );

    \I__6293\ : InMux
    port map (
            O => \N__27603\,
            I => \N__27569\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__27600\,
            I => \N__27566\
        );

    \I__6291\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27563\
        );

    \I__6290\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27558\
        );

    \I__6289\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27558\
        );

    \I__6288\ : InMux
    port map (
            O => \N__27594\,
            I => \N__27555\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__27591\,
            I => \N__27545\
        );

    \I__6286\ : Span4Mux_h
    port map (
            O => \N__27586\,
            I => \N__27545\
        );

    \I__6285\ : Span4Mux_v
    port map (
            O => \N__27583\,
            I => \N__27545\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__27578\,
            I => \N__27545\
        );

    \I__6283\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27542\
        );

    \I__6282\ : Sp12to4
    port map (
            O => \N__27572\,
            I => \N__27529\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__27569\,
            I => \N__27529\
        );

    \I__6280\ : Sp12to4
    port map (
            O => \N__27566\,
            I => \N__27529\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__27563\,
            I => \N__27529\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__27558\,
            I => \N__27529\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__27555\,
            I => \N__27529\
        );

    \I__6276\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27526\
        );

    \I__6275\ : Span4Mux_v
    port map (
            O => \N__27545\,
            I => \N__27523\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__27542\,
            I => \N__27518\
        );

    \I__6273\ : Span12Mux_v
    port map (
            O => \N__27529\,
            I => \N__27518\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__27526\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__6271\ : Odrv4
    port map (
            O => \N__27523\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__6270\ : Odrv12
    port map (
            O => \N__27518\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__27511\,
            I => \N__27508\
        );

    \I__6268\ : InMux
    port map (
            O => \N__27508\,
            I => \N__27505\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__27505\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_8\
        );

    \I__6266\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27498\
        );

    \I__6265\ : CascadeMux
    port map (
            O => \N__27501\,
            I => \N__27490\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__27498\,
            I => \N__27486\
        );

    \I__6263\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27483\
        );

    \I__6262\ : InMux
    port map (
            O => \N__27496\,
            I => \N__27477\
        );

    \I__6261\ : InMux
    port map (
            O => \N__27495\,
            I => \N__27474\
        );

    \I__6260\ : InMux
    port map (
            O => \N__27494\,
            I => \N__27471\
        );

    \I__6259\ : IoInMux
    port map (
            O => \N__27493\,
            I => \N__27468\
        );

    \I__6258\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27465\
        );

    \I__6257\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27462\
        );

    \I__6256\ : Span4Mux_v
    port map (
            O => \N__27486\,
            I => \N__27454\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__27483\,
            I => \N__27454\
        );

    \I__6254\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27445\
        );

    \I__6253\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27445\
        );

    \I__6252\ : InMux
    port map (
            O => \N__27480\,
            I => \N__27442\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__27477\,
            I => \N__27437\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__27474\,
            I => \N__27437\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__27471\,
            I => \N__27434\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__27468\,
            I => \N__27431\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__27465\,
            I => \N__27426\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__27462\,
            I => \N__27426\
        );

    \I__6245\ : InMux
    port map (
            O => \N__27461\,
            I => \N__27419\
        );

    \I__6244\ : InMux
    port map (
            O => \N__27460\,
            I => \N__27419\
        );

    \I__6243\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27419\
        );

    \I__6242\ : Sp12to4
    port map (
            O => \N__27454\,
            I => \N__27416\
        );

    \I__6241\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27409\
        );

    \I__6240\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27409\
        );

    \I__6239\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27409\
        );

    \I__6238\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27406\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N__27403\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27400\
        );

    \I__6235\ : Span4Mux_v
    port map (
            O => \N__27437\,
            I => \N__27397\
        );

    \I__6234\ : Span4Mux_v
    port map (
            O => \N__27434\,
            I => \N__27394\
        );

    \I__6233\ : IoSpan4Mux
    port map (
            O => \N__27431\,
            I => \N__27391\
        );

    \I__6232\ : Span12Mux_v
    port map (
            O => \N__27426\,
            I => \N__27388\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__27419\,
            I => \N__27383\
        );

    \I__6230\ : Span12Mux_s9_h
    port map (
            O => \N__27416\,
            I => \N__27383\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__27409\,
            I => \N__27374\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__27406\,
            I => \N__27374\
        );

    \I__6227\ : Sp12to4
    port map (
            O => \N__27403\,
            I => \N__27374\
        );

    \I__6226\ : Sp12to4
    port map (
            O => \N__27400\,
            I => \N__27374\
        );

    \I__6225\ : Span4Mux_h
    port map (
            O => \N__27397\,
            I => \N__27371\
        );

    \I__6224\ : Span4Mux_h
    port map (
            O => \N__27394\,
            I => \N__27368\
        );

    \I__6223\ : Span4Mux_s2_h
    port map (
            O => \N__27391\,
            I => \N__27365\
        );

    \I__6222\ : Span12Mux_h
    port map (
            O => \N__27388\,
            I => \N__27362\
        );

    \I__6221\ : Span12Mux_h
    port map (
            O => \N__27383\,
            I => \N__27359\
        );

    \I__6220\ : Span12Mux_v
    port map (
            O => \N__27374\,
            I => \N__27356\
        );

    \I__6219\ : Span4Mux_h
    port map (
            O => \N__27371\,
            I => \N__27351\
        );

    \I__6218\ : Span4Mux_v
    port map (
            O => \N__27368\,
            I => \N__27351\
        );

    \I__6217\ : Span4Mux_h
    port map (
            O => \N__27365\,
            I => \N__27348\
        );

    \I__6216\ : Odrv12
    port map (
            O => \N__27362\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6215\ : Odrv12
    port map (
            O => \N__27359\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6214\ : Odrv12
    port map (
            O => \N__27356\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6213\ : Odrv4
    port map (
            O => \N__27351\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__27348\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6211\ : CascadeMux
    port map (
            O => \N__27337\,
            I => \this_vga_signals.M_this_external_address_d_5Z0Z_13_cascade_\
        );

    \I__6210\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27331\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__27331\,
            I => \N__27327\
        );

    \I__6208\ : CascadeMux
    port map (
            O => \N__27330\,
            I => \N__27324\
        );

    \I__6207\ : Span4Mux_h
    port map (
            O => \N__27327\,
            I => \N__27321\
        );

    \I__6206\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27318\
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__27321\,
            I => \this_vga_signals.M_this_state_d_1_sqmuxaZ0\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__27318\,
            I => \this_vga_signals.M_this_state_d_1_sqmuxaZ0\
        );

    \I__6203\ : CascadeMux
    port map (
            O => \N__27313\,
            I => \N__27310\
        );

    \I__6202\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27304\
        );

    \I__6201\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27304\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__27304\,
            I => \this_vga_signals.M_this_state_d_0_sqmuxaZ0Z_1\
        );

    \I__6199\ : CascadeMux
    port map (
            O => \N__27301\,
            I => \this_vga_signals.un1_M_this_state_q_21_0_cascade_\
        );

    \I__6198\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27295\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__27295\,
            I => \this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_13\
        );

    \I__6196\ : SRMux
    port map (
            O => \N__27292\,
            I => \N__27256\
        );

    \I__6195\ : SRMux
    port map (
            O => \N__27291\,
            I => \N__27256\
        );

    \I__6194\ : SRMux
    port map (
            O => \N__27290\,
            I => \N__27256\
        );

    \I__6193\ : SRMux
    port map (
            O => \N__27289\,
            I => \N__27256\
        );

    \I__6192\ : SRMux
    port map (
            O => \N__27288\,
            I => \N__27256\
        );

    \I__6191\ : SRMux
    port map (
            O => \N__27287\,
            I => \N__27256\
        );

    \I__6190\ : SRMux
    port map (
            O => \N__27286\,
            I => \N__27256\
        );

    \I__6189\ : SRMux
    port map (
            O => \N__27285\,
            I => \N__27256\
        );

    \I__6188\ : SRMux
    port map (
            O => \N__27284\,
            I => \N__27256\
        );

    \I__6187\ : SRMux
    port map (
            O => \N__27283\,
            I => \N__27256\
        );

    \I__6186\ : SRMux
    port map (
            O => \N__27282\,
            I => \N__27256\
        );

    \I__6185\ : SRMux
    port map (
            O => \N__27281\,
            I => \N__27256\
        );

    \I__6184\ : GlobalMux
    port map (
            O => \N__27256\,
            I => \N__27253\
        );

    \I__6183\ : gio2CtrlBuf
    port map (
            O => \N__27253\,
            I => \N_989_g\
        );

    \I__6182\ : InMux
    port map (
            O => \N__27250\,
            I => \N__27247\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__27247\,
            I => \N__27243\
        );

    \I__6180\ : InMux
    port map (
            O => \N__27246\,
            I => \N__27240\
        );

    \I__6179\ : Odrv4
    port map (
            O => \N__27243\,
            I => \this_vga_signals.N_469\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__27240\,
            I => \this_vga_signals.N_469\
        );

    \I__6177\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27232\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__27232\,
            I => \N__27228\
        );

    \I__6175\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27223\
        );

    \I__6174\ : Span4Mux_v
    port map (
            O => \N__27228\,
            I => \N__27220\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__27227\,
            I => \N__27217\
        );

    \I__6172\ : InMux
    port map (
            O => \N__27226\,
            I => \N__27212\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__27223\,
            I => \N__27209\
        );

    \I__6170\ : Span4Mux_h
    port map (
            O => \N__27220\,
            I => \N__27203\
        );

    \I__6169\ : InMux
    port map (
            O => \N__27217\,
            I => \N__27200\
        );

    \I__6168\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27195\
        );

    \I__6167\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27195\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__27212\,
            I => \N__27190\
        );

    \I__6165\ : Span4Mux_h
    port map (
            O => \N__27209\,
            I => \N__27190\
        );

    \I__6164\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27185\
        );

    \I__6163\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27185\
        );

    \I__6162\ : InMux
    port map (
            O => \N__27206\,
            I => \N__27182\
        );

    \I__6161\ : Odrv4
    port map (
            O => \N__27203\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__27200\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__27195\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__27190\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__27185\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__27182\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__6155\ : InMux
    port map (
            O => \N__27169\,
            I => \N__27162\
        );

    \I__6154\ : InMux
    port map (
            O => \N__27168\,
            I => \N__27162\
        );

    \I__6153\ : InMux
    port map (
            O => \N__27167\,
            I => \N__27155\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__27162\,
            I => \N__27152\
        );

    \I__6151\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27149\
        );

    \I__6150\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27146\
        );

    \I__6149\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27143\
        );

    \I__6148\ : InMux
    port map (
            O => \N__27158\,
            I => \N__27140\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__27155\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__6146\ : Odrv12
    port map (
            O => \N__27152\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__27149\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__27146\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__27143\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__27140\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__6141\ : CascadeMux
    port map (
            O => \N__27127\,
            I => \N__27123\
        );

    \I__6140\ : CascadeMux
    port map (
            O => \N__27126\,
            I => \N__27120\
        );

    \I__6139\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27115\
        );

    \I__6138\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27112\
        );

    \I__6137\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27107\
        );

    \I__6136\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27107\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__27115\,
            I => \N__27104\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__27112\,
            I => \N__27099\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27099\
        );

    \I__6132\ : Span4Mux_v
    port map (
            O => \N__27104\,
            I => \N__27093\
        );

    \I__6131\ : Span4Mux_v
    port map (
            O => \N__27099\,
            I => \N__27090\
        );

    \I__6130\ : CascadeMux
    port map (
            O => \N__27098\,
            I => \N__27087\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__27097\,
            I => \N__27083\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__27096\,
            I => \N__27080\
        );

    \I__6127\ : Span4Mux_h
    port map (
            O => \N__27093\,
            I => \N__27075\
        );

    \I__6126\ : Span4Mux_h
    port map (
            O => \N__27090\,
            I => \N__27075\
        );

    \I__6125\ : InMux
    port map (
            O => \N__27087\,
            I => \N__27070\
        );

    \I__6124\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27070\
        );

    \I__6123\ : InMux
    port map (
            O => \N__27083\,
            I => \N__27065\
        );

    \I__6122\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27065\
        );

    \I__6121\ : Sp12to4
    port map (
            O => \N__27075\,
            I => \N__27058\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__27070\,
            I => \N__27058\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__27065\,
            I => \N__27058\
        );

    \I__6118\ : Span12Mux_h
    port map (
            O => \N__27058\,
            I => \N__27055\
        );

    \I__6117\ : Odrv12
    port map (
            O => \N__27055\,
            I => port_enb_c
        );

    \I__6116\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27046\
        );

    \I__6115\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27046\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__27046\,
            I => \N__27039\
        );

    \I__6113\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27036\
        );

    \I__6112\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27031\
        );

    \I__6111\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27031\
        );

    \I__6110\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27026\
        );

    \I__6109\ : Span4Mux_h
    port map (
            O => \N__27039\,
            I => \N__27023\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__27036\,
            I => \N__27018\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__27031\,
            I => \N__27018\
        );

    \I__6106\ : InMux
    port map (
            O => \N__27030\,
            I => \N__27013\
        );

    \I__6105\ : InMux
    port map (
            O => \N__27029\,
            I => \N__27013\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__27026\,
            I => \M_this_delay_clk_out_0\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__27023\,
            I => \M_this_delay_clk_out_0\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__27018\,
            I => \M_this_delay_clk_out_0\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__27013\,
            I => \M_this_delay_clk_out_0\
        );

    \I__6100\ : InMux
    port map (
            O => \N__27004\,
            I => \N__26999\
        );

    \I__6099\ : InMux
    port map (
            O => \N__27003\,
            I => \N__26996\
        );

    \I__6098\ : CascadeMux
    port map (
            O => \N__27002\,
            I => \N__26992\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__26999\,
            I => \N__26988\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__26996\,
            I => \N__26985\
        );

    \I__6095\ : CascadeMux
    port map (
            O => \N__26995\,
            I => \N__26982\
        );

    \I__6094\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26979\
        );

    \I__6093\ : CascadeMux
    port map (
            O => \N__26991\,
            I => \N__26975\
        );

    \I__6092\ : Span4Mux_v
    port map (
            O => \N__26988\,
            I => \N__26969\
        );

    \I__6091\ : Span4Mux_v
    port map (
            O => \N__26985\,
            I => \N__26969\
        );

    \I__6090\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26966\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__26979\,
            I => \N__26963\
        );

    \I__6088\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26960\
        );

    \I__6087\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26957\
        );

    \I__6086\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26954\
        );

    \I__6085\ : Span4Mux_h
    port map (
            O => \N__26969\,
            I => \N__26948\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__26966\,
            I => \N__26948\
        );

    \I__6083\ : Span4Mux_v
    port map (
            O => \N__26963\,
            I => \N__26944\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__26960\,
            I => \N__26937\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__26957\,
            I => \N__26937\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__26954\,
            I => \N__26937\
        );

    \I__6079\ : InMux
    port map (
            O => \N__26953\,
            I => \N__26934\
        );

    \I__6078\ : Span4Mux_v
    port map (
            O => \N__26948\,
            I => \N__26931\
        );

    \I__6077\ : InMux
    port map (
            O => \N__26947\,
            I => \N__26928\
        );

    \I__6076\ : Span4Mux_h
    port map (
            O => \N__26944\,
            I => \N__26921\
        );

    \I__6075\ : Span4Mux_v
    port map (
            O => \N__26937\,
            I => \N__26921\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__26934\,
            I => \N__26921\
        );

    \I__6073\ : Sp12to4
    port map (
            O => \N__26931\,
            I => \N__26918\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__26928\,
            I => \N__26915\
        );

    \I__6071\ : Span4Mux_v
    port map (
            O => \N__26921\,
            I => \N__26912\
        );

    \I__6070\ : Span12Mux_s10_h
    port map (
            O => \N__26918\,
            I => \N__26909\
        );

    \I__6069\ : Sp12to4
    port map (
            O => \N__26915\,
            I => \N__26906\
        );

    \I__6068\ : Sp12to4
    port map (
            O => \N__26912\,
            I => \N__26903\
        );

    \I__6067\ : Span12Mux_v
    port map (
            O => \N__26909\,
            I => \N__26900\
        );

    \I__6066\ : Span12Mux_v
    port map (
            O => \N__26906\,
            I => \N__26895\
        );

    \I__6065\ : Span12Mux_h
    port map (
            O => \N__26903\,
            I => \N__26895\
        );

    \I__6064\ : Odrv12
    port map (
            O => \N__26900\,
            I => port_address_in_2
        );

    \I__6063\ : Odrv12
    port map (
            O => \N__26895\,
            I => port_address_in_2
        );

    \I__6062\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26886\
        );

    \I__6061\ : CascadeMux
    port map (
            O => \N__26889\,
            I => \N__26883\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__26886\,
            I => \N__26879\
        );

    \I__6059\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26874\
        );

    \I__6058\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26870\
        );

    \I__6057\ : Span4Mux_v
    port map (
            O => \N__26879\,
            I => \N__26867\
        );

    \I__6056\ : InMux
    port map (
            O => \N__26878\,
            I => \N__26864\
        );

    \I__6055\ : CascadeMux
    port map (
            O => \N__26877\,
            I => \N__26860\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__26874\,
            I => \N__26857\
        );

    \I__6053\ : InMux
    port map (
            O => \N__26873\,
            I => \N__26853\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__26870\,
            I => \N__26846\
        );

    \I__6051\ : Sp12to4
    port map (
            O => \N__26867\,
            I => \N__26846\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__26864\,
            I => \N__26846\
        );

    \I__6049\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26843\
        );

    \I__6048\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26840\
        );

    \I__6047\ : Span4Mux_v
    port map (
            O => \N__26857\,
            I => \N__26837\
        );

    \I__6046\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26834\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__26853\,
            I => \N__26831\
        );

    \I__6044\ : Span12Mux_h
    port map (
            O => \N__26846\,
            I => \N__26826\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__26843\,
            I => \N__26826\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26823\
        );

    \I__6041\ : Span4Mux_h
    port map (
            O => \N__26837\,
            I => \N__26818\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__26834\,
            I => \N__26818\
        );

    \I__6039\ : Span12Mux_v
    port map (
            O => \N__26831\,
            I => \N__26815\
        );

    \I__6038\ : Span12Mux_v
    port map (
            O => \N__26826\,
            I => \N__26812\
        );

    \I__6037\ : Span12Mux_v
    port map (
            O => \N__26823\,
            I => \N__26807\
        );

    \I__6036\ : Sp12to4
    port map (
            O => \N__26818\,
            I => \N__26807\
        );

    \I__6035\ : Odrv12
    port map (
            O => \N__26815\,
            I => port_address_in_0
        );

    \I__6034\ : Odrv12
    port map (
            O => \N__26812\,
            I => port_address_in_0
        );

    \I__6033\ : Odrv12
    port map (
            O => \N__26807\,
            I => port_address_in_0
        );

    \I__6032\ : CascadeMux
    port map (
            O => \N__26800\,
            I => \N__26797\
        );

    \I__6031\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26793\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__26796\,
            I => \N__26787\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__26793\,
            I => \N__26783\
        );

    \I__6028\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26776\
        );

    \I__6027\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26776\
        );

    \I__6026\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26776\
        );

    \I__6025\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26773\
        );

    \I__6024\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26770\
        );

    \I__6023\ : Span4Mux_v
    port map (
            O => \N__26783\,
            I => \N__26766\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__26776\,
            I => \N__26759\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__26773\,
            I => \N__26759\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__26770\,
            I => \N__26759\
        );

    \I__6019\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26756\
        );

    \I__6018\ : Sp12to4
    port map (
            O => \N__26766\,
            I => \N__26753\
        );

    \I__6017\ : Sp12to4
    port map (
            O => \N__26759\,
            I => \N__26748\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__26756\,
            I => \N__26748\
        );

    \I__6015\ : Span12Mux_h
    port map (
            O => \N__26753\,
            I => \N__26745\
        );

    \I__6014\ : Span12Mux_v
    port map (
            O => \N__26748\,
            I => \N__26742\
        );

    \I__6013\ : Span12Mux_v
    port map (
            O => \N__26745\,
            I => \N__26737\
        );

    \I__6012\ : Span12Mux_h
    port map (
            O => \N__26742\,
            I => \N__26737\
        );

    \I__6011\ : Odrv12
    port map (
            O => \N__26737\,
            I => port_address_in_3
        );

    \I__6010\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26725\
        );

    \I__6009\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26725\
        );

    \I__6008\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26725\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__26725\,
            I => \N__26721\
        );

    \I__6006\ : InMux
    port map (
            O => \N__26724\,
            I => \N__26718\
        );

    \I__6005\ : Span4Mux_h
    port map (
            O => \N__26721\,
            I => \N__26710\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__26718\,
            I => \N__26710\
        );

    \I__6003\ : InMux
    port map (
            O => \N__26717\,
            I => \N__26707\
        );

    \I__6002\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26704\
        );

    \I__6001\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26701\
        );

    \I__6000\ : Span4Mux_h
    port map (
            O => \N__26710\,
            I => \N__26696\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__26707\,
            I => \N__26696\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__26704\,
            I => \N__26691\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__26701\,
            I => \N__26691\
        );

    \I__5996\ : Span4Mux_v
    port map (
            O => \N__26696\,
            I => \N__26688\
        );

    \I__5995\ : Span4Mux_v
    port map (
            O => \N__26691\,
            I => \N__26685\
        );

    \I__5994\ : Sp12to4
    port map (
            O => \N__26688\,
            I => \N__26680\
        );

    \I__5993\ : Sp12to4
    port map (
            O => \N__26685\,
            I => \N__26680\
        );

    \I__5992\ : Span12Mux_h
    port map (
            O => \N__26680\,
            I => \N__26677\
        );

    \I__5991\ : Odrv12
    port map (
            O => \N__26677\,
            I => port_address_in_1
        );

    \I__5990\ : CascadeMux
    port map (
            O => \N__26674\,
            I => \N__26671\
        );

    \I__5989\ : InMux
    port map (
            O => \N__26671\,
            I => \N__26668\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__26668\,
            I => \N__26665\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__26665\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_10\
        );

    \I__5986\ : InMux
    port map (
            O => \N__26662\,
            I => \N__26659\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__26659\,
            I => \this_vga_signals.M_this_map_address_d_8_mZ0Z_1\
        );

    \I__5984\ : CascadeMux
    port map (
            O => \N__26656\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_1_cascade_\
        );

    \I__5983\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26650\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__26650\,
            I => \un1_M_this_map_address_q_cry_0_c_RNI6GRRZ0\
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__26647\,
            I => \N__26644\
        );

    \I__5980\ : CascadeBuf
    port map (
            O => \N__26644\,
            I => \N__26641\
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__26641\,
            I => \N__26638\
        );

    \I__5978\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26635\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__26635\,
            I => \N__26632\
        );

    \I__5976\ : Span4Mux_v
    port map (
            O => \N__26632\,
            I => \N__26629\
        );

    \I__5975\ : Span4Mux_h
    port map (
            O => \N__26629\,
            I => \N__26623\
        );

    \I__5974\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26620\
        );

    \I__5973\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26617\
        );

    \I__5972\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26614\
        );

    \I__5971\ : Span4Mux_v
    port map (
            O => \N__26623\,
            I => \N__26611\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__26620\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__26617\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__26614\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__5967\ : Odrv4
    port map (
            O => \N__26611\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__5966\ : CascadeMux
    port map (
            O => \N__26602\,
            I => \this_vga_signals.M_this_map_address_d_8_mZ0Z_3_cascade_\
        );

    \I__5965\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26596\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__26596\,
            I => \un1_M_this_map_address_q_cry_2_c_RNIAMTRZ0\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__26593\,
            I => \N__26590\
        );

    \I__5962\ : CascadeBuf
    port map (
            O => \N__26590\,
            I => \N__26587\
        );

    \I__5961\ : CascadeMux
    port map (
            O => \N__26587\,
            I => \N__26584\
        );

    \I__5960\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26581\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__26581\,
            I => \N__26578\
        );

    \I__5958\ : Span4Mux_s3_v
    port map (
            O => \N__26578\,
            I => \N__26575\
        );

    \I__5957\ : Span4Mux_h
    port map (
            O => \N__26575\,
            I => \N__26569\
        );

    \I__5956\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26566\
        );

    \I__5955\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26563\
        );

    \I__5954\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26560\
        );

    \I__5953\ : Span4Mux_v
    port map (
            O => \N__26569\,
            I => \N__26557\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__26566\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__26563\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__26560\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__26557\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__5948\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26545\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__26545\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_3\
        );

    \I__5946\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26539\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__26539\,
            I => \this_vga_signals.M_this_map_address_d_8_mZ0Z_4\
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__26536\,
            I => \N__26533\
        );

    \I__5943\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26530\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__26530\,
            I => \N__26527\
        );

    \I__5941\ : Odrv4
    port map (
            O => \N__26527\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_4\
        );

    \I__5940\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26521\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__26521\,
            I => \un1_M_this_map_address_q_cry_3_c_RNICPURZ0\
        );

    \I__5938\ : CascadeMux
    port map (
            O => \N__26518\,
            I => \N__26515\
        );

    \I__5937\ : CascadeBuf
    port map (
            O => \N__26515\,
            I => \N__26512\
        );

    \I__5936\ : CascadeMux
    port map (
            O => \N__26512\,
            I => \N__26509\
        );

    \I__5935\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26506\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__26506\,
            I => \N__26503\
        );

    \I__5933\ : Span4Mux_s3_v
    port map (
            O => \N__26503\,
            I => \N__26500\
        );

    \I__5932\ : Span4Mux_h
    port map (
            O => \N__26500\,
            I => \N__26494\
        );

    \I__5931\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26489\
        );

    \I__5930\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26489\
        );

    \I__5929\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26486\
        );

    \I__5928\ : Span4Mux_v
    port map (
            O => \N__26494\,
            I => \N__26483\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__26489\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__26486\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__26483\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__5924\ : InMux
    port map (
            O => \N__26476\,
            I => \N__26468\
        );

    \I__5923\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26465\
        );

    \I__5922\ : InMux
    port map (
            O => \N__26474\,
            I => \N__26459\
        );

    \I__5921\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26454\
        );

    \I__5920\ : InMux
    port map (
            O => \N__26472\,
            I => \N__26454\
        );

    \I__5919\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26450\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__26468\,
            I => \N__26445\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__26465\,
            I => \N__26445\
        );

    \I__5916\ : InMux
    port map (
            O => \N__26464\,
            I => \N__26442\
        );

    \I__5915\ : InMux
    port map (
            O => \N__26463\,
            I => \N__26437\
        );

    \I__5914\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26437\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__26459\,
            I => \N__26433\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__26454\,
            I => \N__26430\
        );

    \I__5911\ : InMux
    port map (
            O => \N__26453\,
            I => \N__26427\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__26450\,
            I => \N__26420\
        );

    \I__5909\ : Span4Mux_h
    port map (
            O => \N__26445\,
            I => \N__26420\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__26442\,
            I => \N__26417\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__26437\,
            I => \N__26414\
        );

    \I__5906\ : InMux
    port map (
            O => \N__26436\,
            I => \N__26411\
        );

    \I__5905\ : Span4Mux_h
    port map (
            O => \N__26433\,
            I => \N__26404\
        );

    \I__5904\ : Span4Mux_v
    port map (
            O => \N__26430\,
            I => \N__26404\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__26427\,
            I => \N__26404\
        );

    \I__5902\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26401\
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__26425\,
            I => \N__26396\
        );

    \I__5900\ : Span4Mux_v
    port map (
            O => \N__26420\,
            I => \N__26393\
        );

    \I__5899\ : Span4Mux_v
    port map (
            O => \N__26417\,
            I => \N__26386\
        );

    \I__5898\ : Span4Mux_h
    port map (
            O => \N__26414\,
            I => \N__26386\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__26411\,
            I => \N__26386\
        );

    \I__5896\ : Span4Mux_v
    port map (
            O => \N__26404\,
            I => \N__26381\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__26401\,
            I => \N__26381\
        );

    \I__5894\ : InMux
    port map (
            O => \N__26400\,
            I => \N__26378\
        );

    \I__5893\ : InMux
    port map (
            O => \N__26399\,
            I => \N__26373\
        );

    \I__5892\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26373\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__26393\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5890\ : Odrv4
    port map (
            O => \N__26386\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__26381\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__26378\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__26373\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__26362\,
            I => \N__26357\
        );

    \I__5885\ : InMux
    port map (
            O => \N__26361\,
            I => \N__26354\
        );

    \I__5884\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26351\
        );

    \I__5883\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26348\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__26354\,
            I => \N__26345\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__26351\,
            I => \N__26340\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__26348\,
            I => \N__26340\
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__26345\,
            I => \un1_M_this_state_q_12_0\
        );

    \I__5878\ : Odrv4
    port map (
            O => \N__26340\,
            I => \un1_M_this_state_q_12_0\
        );

    \I__5877\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26332\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__26332\,
            I => \this_vga_signals.M_this_map_address_d_5_mZ0Z_8\
        );

    \I__5875\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26317\
        );

    \I__5874\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26317\
        );

    \I__5873\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26317\
        );

    \I__5872\ : InMux
    port map (
            O => \N__26326\,
            I => \N__26310\
        );

    \I__5871\ : InMux
    port map (
            O => \N__26325\,
            I => \N__26310\
        );

    \I__5870\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26310\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__26317\,
            I => \N__26303\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__26310\,
            I => \N__26300\
        );

    \I__5867\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26297\
        );

    \I__5866\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26290\
        );

    \I__5865\ : InMux
    port map (
            O => \N__26307\,
            I => \N__26290\
        );

    \I__5864\ : InMux
    port map (
            O => \N__26306\,
            I => \N__26290\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__26303\,
            I => \this_vga_signals.un1_M_this_map_ram_write_en_0\
        );

    \I__5862\ : Odrv4
    port map (
            O => \N__26300\,
            I => \this_vga_signals.un1_M_this_map_ram_write_en_0\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__26297\,
            I => \this_vga_signals.un1_M_this_map_ram_write_en_0\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__26290\,
            I => \this_vga_signals.un1_M_this_map_ram_write_en_0\
        );

    \I__5859\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26278\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__26278\,
            I => \un1_M_this_map_address_q_cry_7_c_RNIK53SZ0\
        );

    \I__5857\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26272\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__26272\,
            I => \this_vga_signals.M_this_external_address_d_5Z0Z_14\
        );

    \I__5855\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26266\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__26266\,
            I => \this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_14\
        );

    \I__5853\ : CascadeMux
    port map (
            O => \N__26263\,
            I => \N__26260\
        );

    \I__5852\ : CascadeBuf
    port map (
            O => \N__26260\,
            I => \N__26257\
        );

    \I__5851\ : CascadeMux
    port map (
            O => \N__26257\,
            I => \N__26254\
        );

    \I__5850\ : CascadeBuf
    port map (
            O => \N__26254\,
            I => \N__26251\
        );

    \I__5849\ : CascadeMux
    port map (
            O => \N__26251\,
            I => \N__26248\
        );

    \I__5848\ : CascadeBuf
    port map (
            O => \N__26248\,
            I => \N__26245\
        );

    \I__5847\ : CascadeMux
    port map (
            O => \N__26245\,
            I => \N__26242\
        );

    \I__5846\ : CascadeBuf
    port map (
            O => \N__26242\,
            I => \N__26239\
        );

    \I__5845\ : CascadeMux
    port map (
            O => \N__26239\,
            I => \N__26236\
        );

    \I__5844\ : CascadeBuf
    port map (
            O => \N__26236\,
            I => \N__26233\
        );

    \I__5843\ : CascadeMux
    port map (
            O => \N__26233\,
            I => \N__26230\
        );

    \I__5842\ : CascadeBuf
    port map (
            O => \N__26230\,
            I => \N__26227\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__26227\,
            I => \N__26224\
        );

    \I__5840\ : CascadeBuf
    port map (
            O => \N__26224\,
            I => \N__26221\
        );

    \I__5839\ : CascadeMux
    port map (
            O => \N__26221\,
            I => \N__26218\
        );

    \I__5838\ : CascadeBuf
    port map (
            O => \N__26218\,
            I => \N__26215\
        );

    \I__5837\ : CascadeMux
    port map (
            O => \N__26215\,
            I => \N__26212\
        );

    \I__5836\ : CascadeBuf
    port map (
            O => \N__26212\,
            I => \N__26209\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__26209\,
            I => \N__26206\
        );

    \I__5834\ : CascadeBuf
    port map (
            O => \N__26206\,
            I => \N__26203\
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__26203\,
            I => \N__26200\
        );

    \I__5832\ : CascadeBuf
    port map (
            O => \N__26200\,
            I => \N__26197\
        );

    \I__5831\ : CascadeMux
    port map (
            O => \N__26197\,
            I => \N__26194\
        );

    \I__5830\ : CascadeBuf
    port map (
            O => \N__26194\,
            I => \N__26191\
        );

    \I__5829\ : CascadeMux
    port map (
            O => \N__26191\,
            I => \N__26188\
        );

    \I__5828\ : CascadeBuf
    port map (
            O => \N__26188\,
            I => \N__26185\
        );

    \I__5827\ : CascadeMux
    port map (
            O => \N__26185\,
            I => \N__26182\
        );

    \I__5826\ : CascadeBuf
    port map (
            O => \N__26182\,
            I => \N__26179\
        );

    \I__5825\ : CascadeMux
    port map (
            O => \N__26179\,
            I => \N__26176\
        );

    \I__5824\ : CascadeBuf
    port map (
            O => \N__26176\,
            I => \N__26173\
        );

    \I__5823\ : CascadeMux
    port map (
            O => \N__26173\,
            I => \N__26170\
        );

    \I__5822\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26167\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__26167\,
            I => \N__26162\
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__26166\,
            I => \N__26159\
        );

    \I__5819\ : InMux
    port map (
            O => \N__26165\,
            I => \N__26156\
        );

    \I__5818\ : Span4Mux_s1_v
    port map (
            O => \N__26162\,
            I => \N__26153\
        );

    \I__5817\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26149\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__26156\,
            I => \N__26146\
        );

    \I__5815\ : Sp12to4
    port map (
            O => \N__26153\,
            I => \N__26143\
        );

    \I__5814\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26140\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__26149\,
            I => \N__26135\
        );

    \I__5812\ : Span4Mux_h
    port map (
            O => \N__26146\,
            I => \N__26135\
        );

    \I__5811\ : Span12Mux_v
    port map (
            O => \N__26143\,
            I => \N__26132\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__26140\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__5809\ : Odrv4
    port map (
            O => \N__26135\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__5808\ : Odrv12
    port map (
            O => \N__26132\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__5807\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26122\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__26122\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__26119\,
            I => \N__26116\
        );

    \I__5804\ : CascadeBuf
    port map (
            O => \N__26116\,
            I => \N__26113\
        );

    \I__5803\ : CascadeMux
    port map (
            O => \N__26113\,
            I => \N__26110\
        );

    \I__5802\ : InMux
    port map (
            O => \N__26110\,
            I => \N__26107\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__26104\
        );

    \I__5800\ : Span4Mux_h
    port map (
            O => \N__26104\,
            I => \N__26101\
        );

    \I__5799\ : Span4Mux_h
    port map (
            O => \N__26101\,
            I => \N__26097\
        );

    \I__5798\ : InMux
    port map (
            O => \N__26100\,
            I => \N__26093\
        );

    \I__5797\ : Span4Mux_v
    port map (
            O => \N__26097\,
            I => \N__26089\
        );

    \I__5796\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26086\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26083\
        );

    \I__5794\ : InMux
    port map (
            O => \N__26092\,
            I => \N__26080\
        );

    \I__5793\ : Span4Mux_v
    port map (
            O => \N__26089\,
            I => \N__26077\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__26086\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__26083\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__26080\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__26077\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__5788\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26065\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__26065\,
            I => \this_vga_signals.M_this_map_address_d_8_mZ0Z_0\
        );

    \I__5786\ : CascadeMux
    port map (
            O => \N__26062\,
            I => \N__26059\
        );

    \I__5785\ : CascadeBuf
    port map (
            O => \N__26059\,
            I => \N__26056\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__26056\,
            I => \N__26053\
        );

    \I__5783\ : CascadeBuf
    port map (
            O => \N__26053\,
            I => \N__26050\
        );

    \I__5782\ : CascadeMux
    port map (
            O => \N__26050\,
            I => \N__26047\
        );

    \I__5781\ : CascadeBuf
    port map (
            O => \N__26047\,
            I => \N__26044\
        );

    \I__5780\ : CascadeMux
    port map (
            O => \N__26044\,
            I => \N__26041\
        );

    \I__5779\ : CascadeBuf
    port map (
            O => \N__26041\,
            I => \N__26038\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__26038\,
            I => \N__26035\
        );

    \I__5777\ : CascadeBuf
    port map (
            O => \N__26035\,
            I => \N__26032\
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__5775\ : CascadeBuf
    port map (
            O => \N__26029\,
            I => \N__26026\
        );

    \I__5774\ : CascadeMux
    port map (
            O => \N__26026\,
            I => \N__26023\
        );

    \I__5773\ : CascadeBuf
    port map (
            O => \N__26023\,
            I => \N__26020\
        );

    \I__5772\ : CascadeMux
    port map (
            O => \N__26020\,
            I => \N__26017\
        );

    \I__5771\ : CascadeBuf
    port map (
            O => \N__26017\,
            I => \N__26014\
        );

    \I__5770\ : CascadeMux
    port map (
            O => \N__26014\,
            I => \N__26011\
        );

    \I__5769\ : CascadeBuf
    port map (
            O => \N__26011\,
            I => \N__26008\
        );

    \I__5768\ : CascadeMux
    port map (
            O => \N__26008\,
            I => \N__26005\
        );

    \I__5767\ : CascadeBuf
    port map (
            O => \N__26005\,
            I => \N__26002\
        );

    \I__5766\ : CascadeMux
    port map (
            O => \N__26002\,
            I => \N__25999\
        );

    \I__5765\ : CascadeBuf
    port map (
            O => \N__25999\,
            I => \N__25996\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__25996\,
            I => \N__25993\
        );

    \I__5763\ : CascadeBuf
    port map (
            O => \N__25993\,
            I => \N__25990\
        );

    \I__5762\ : CascadeMux
    port map (
            O => \N__25990\,
            I => \N__25987\
        );

    \I__5761\ : CascadeBuf
    port map (
            O => \N__25987\,
            I => \N__25984\
        );

    \I__5760\ : CascadeMux
    port map (
            O => \N__25984\,
            I => \N__25981\
        );

    \I__5759\ : CascadeBuf
    port map (
            O => \N__25981\,
            I => \N__25978\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__25978\,
            I => \N__25975\
        );

    \I__5757\ : CascadeBuf
    port map (
            O => \N__25975\,
            I => \N__25972\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__25972\,
            I => \N__25969\
        );

    \I__5755\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25966\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__25966\,
            I => \N__25963\
        );

    \I__5753\ : Span4Mux_s3_v
    port map (
            O => \N__25963\,
            I => \N__25958\
        );

    \I__5752\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25955\
        );

    \I__5751\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25952\
        );

    \I__5750\ : Span4Mux_v
    port map (
            O => \N__25958\,
            I => \N__25948\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__25955\,
            I => \N__25943\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__25952\,
            I => \N__25943\
        );

    \I__5747\ : InMux
    port map (
            O => \N__25951\,
            I => \N__25940\
        );

    \I__5746\ : Span4Mux_v
    port map (
            O => \N__25948\,
            I => \N__25937\
        );

    \I__5745\ : Span4Mux_v
    port map (
            O => \N__25943\,
            I => \N__25934\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__25940\,
            I => \N__25929\
        );

    \I__5743\ : Sp12to4
    port map (
            O => \N__25937\,
            I => \N__25929\
        );

    \I__5742\ : Odrv4
    port map (
            O => \N__25934\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5741\ : Odrv12
    port map (
            O => \N__25929\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5740\ : InMux
    port map (
            O => \N__25924\,
            I => \N__25921\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__25921\,
            I => \N__25918\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__25918\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0\
        );

    \I__5737\ : InMux
    port map (
            O => \N__25915\,
            I => \N__25912\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__25912\,
            I => \N__25909\
        );

    \I__5735\ : Span4Mux_h
    port map (
            O => \N__25909\,
            I => \N__25906\
        );

    \I__5734\ : Odrv4
    port map (
            O => \N__25906\,
            I => \this_vga_signals.N_291\
        );

    \I__5733\ : CascadeMux
    port map (
            O => \N__25903\,
            I => \N__25899\
        );

    \I__5732\ : InMux
    port map (
            O => \N__25902\,
            I => \N__25895\
        );

    \I__5731\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25892\
        );

    \I__5730\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25889\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__25895\,
            I => \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__25892\,
            I => \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__25889\,
            I => \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__25882\,
            I => \N__25878\
        );

    \I__5725\ : InMux
    port map (
            O => \N__25881\,
            I => \N__25873\
        );

    \I__5724\ : InMux
    port map (
            O => \N__25878\,
            I => \N__25866\
        );

    \I__5723\ : InMux
    port map (
            O => \N__25877\,
            I => \N__25866\
        );

    \I__5722\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25866\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__25873\,
            I => \N__25861\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__25866\,
            I => \N__25861\
        );

    \I__5719\ : Span12Mux_v
    port map (
            O => \N__25861\,
            I => \N__25858\
        );

    \I__5718\ : Span12Mux_h
    port map (
            O => \N__25858\,
            I => \N__25855\
        );

    \I__5717\ : Odrv12
    port map (
            O => \N__25855\,
            I => port_address_in_5
        );

    \I__5716\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25843\
        );

    \I__5715\ : InMux
    port map (
            O => \N__25851\,
            I => \N__25843\
        );

    \I__5714\ : InMux
    port map (
            O => \N__25850\,
            I => \N__25843\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__25843\,
            I => \N__25840\
        );

    \I__5712\ : Span4Mux_v
    port map (
            O => \N__25840\,
            I => \N__25836\
        );

    \I__5711\ : InMux
    port map (
            O => \N__25839\,
            I => \N__25833\
        );

    \I__5710\ : Span4Mux_h
    port map (
            O => \N__25836\,
            I => \N__25830\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__25833\,
            I => \N__25827\
        );

    \I__5708\ : Span4Mux_h
    port map (
            O => \N__25830\,
            I => \N__25824\
        );

    \I__5707\ : Span12Mux_h
    port map (
            O => \N__25827\,
            I => \N__25821\
        );

    \I__5706\ : Odrv4
    port map (
            O => \N__25824\,
            I => port_address_in_6
        );

    \I__5705\ : Odrv12
    port map (
            O => \N__25821\,
            I => port_address_in_6
        );

    \I__5704\ : CascadeMux
    port map (
            O => \N__25816\,
            I => \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_4_cascade_\
        );

    \I__5703\ : InMux
    port map (
            O => \N__25813\,
            I => \N__25804\
        );

    \I__5702\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25804\
        );

    \I__5701\ : InMux
    port map (
            O => \N__25811\,
            I => \N__25801\
        );

    \I__5700\ : InMux
    port map (
            O => \N__25810\,
            I => \N__25796\
        );

    \I__5699\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25796\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__25804\,
            I => \this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__25801\,
            I => \this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__25796\,
            I => \this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0\
        );

    \I__5695\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25786\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__25786\,
            I => \N__25783\
        );

    \I__5693\ : Span4Mux_v
    port map (
            O => \N__25783\,
            I => \N__25779\
        );

    \I__5692\ : InMux
    port map (
            O => \N__25782\,
            I => \N__25776\
        );

    \I__5691\ : Span4Mux_h
    port map (
            O => \N__25779\,
            I => \N__25771\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__25776\,
            I => \N__25771\
        );

    \I__5689\ : Odrv4
    port map (
            O => \N__25771\,
            I => \this_vga_signals.N_444_1\
        );

    \I__5688\ : InMux
    port map (
            O => \N__25768\,
            I => \N__25765\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__25765\,
            I => \N__25761\
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__25764\,
            I => \N__25758\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__25761\,
            I => \N__25755\
        );

    \I__5684\ : InMux
    port map (
            O => \N__25758\,
            I => \N__25752\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__25755\,
            I => \this_vga_signals_M_this_state_q_ns_i_o2_0_14\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__25752\,
            I => \this_vga_signals_M_this_state_q_ns_i_o2_0_14\
        );

    \I__5681\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25743\
        );

    \I__5680\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25740\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__25743\,
            I => \N__25735\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__25740\,
            I => \N__25735\
        );

    \I__5677\ : Odrv4
    port map (
            O => \N__25735\,
            I => \M_this_state_q_fastZ0Z_14\
        );

    \I__5676\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25729\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__25729\,
            I => \N__25720\
        );

    \I__5674\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25717\
        );

    \I__5673\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25709\
        );

    \I__5672\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25709\
        );

    \I__5671\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25709\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__25724\,
            I => \N__25705\
        );

    \I__5669\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25702\
        );

    \I__5668\ : Span4Mux_v
    port map (
            O => \N__25720\,
            I => \N__25699\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__25717\,
            I => \N__25696\
        );

    \I__5666\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25693\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__25709\,
            I => \N__25690\
        );

    \I__5664\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25687\
        );

    \I__5663\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25684\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__25702\,
            I => \N__25680\
        );

    \I__5661\ : Sp12to4
    port map (
            O => \N__25699\,
            I => \N__25673\
        );

    \I__5660\ : Sp12to4
    port map (
            O => \N__25696\,
            I => \N__25673\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__25693\,
            I => \N__25673\
        );

    \I__5658\ : Span4Mux_v
    port map (
            O => \N__25690\,
            I => \N__25670\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__25687\,
            I => \N__25667\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__25684\,
            I => \N__25664\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__25683\,
            I => \N__25660\
        );

    \I__5654\ : Span12Mux_v
    port map (
            O => \N__25680\,
            I => \N__25655\
        );

    \I__5653\ : Span12Mux_v
    port map (
            O => \N__25673\,
            I => \N__25655\
        );

    \I__5652\ : Span4Mux_h
    port map (
            O => \N__25670\,
            I => \N__25648\
        );

    \I__5651\ : Span4Mux_h
    port map (
            O => \N__25667\,
            I => \N__25648\
        );

    \I__5650\ : Span4Mux_v
    port map (
            O => \N__25664\,
            I => \N__25648\
        );

    \I__5649\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25645\
        );

    \I__5648\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25642\
        );

    \I__5647\ : Odrv12
    port map (
            O => \N__25655\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__5646\ : Odrv4
    port map (
            O => \N__25648\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__25645\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__25642\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__25633\,
            I => \N__25630\
        );

    \I__5642\ : InMux
    port map (
            O => \N__25630\,
            I => \N__25627\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__25627\,
            I => \N__25624\
        );

    \I__5640\ : Span4Mux_v
    port map (
            O => \N__25624\,
            I => \N__25621\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__25621\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_12\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__25618\,
            I => \N__25615\
        );

    \I__5637\ : CascadeBuf
    port map (
            O => \N__25615\,
            I => \N__25612\
        );

    \I__5636\ : CascadeMux
    port map (
            O => \N__25612\,
            I => \N__25609\
        );

    \I__5635\ : CascadeBuf
    port map (
            O => \N__25609\,
            I => \N__25606\
        );

    \I__5634\ : CascadeMux
    port map (
            O => \N__25606\,
            I => \N__25603\
        );

    \I__5633\ : CascadeBuf
    port map (
            O => \N__25603\,
            I => \N__25600\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__25600\,
            I => \N__25597\
        );

    \I__5631\ : CascadeBuf
    port map (
            O => \N__25597\,
            I => \N__25594\
        );

    \I__5630\ : CascadeMux
    port map (
            O => \N__25594\,
            I => \N__25591\
        );

    \I__5629\ : CascadeBuf
    port map (
            O => \N__25591\,
            I => \N__25588\
        );

    \I__5628\ : CascadeMux
    port map (
            O => \N__25588\,
            I => \N__25585\
        );

    \I__5627\ : CascadeBuf
    port map (
            O => \N__25585\,
            I => \N__25582\
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__25582\,
            I => \N__25579\
        );

    \I__5625\ : CascadeBuf
    port map (
            O => \N__25579\,
            I => \N__25576\
        );

    \I__5624\ : CascadeMux
    port map (
            O => \N__25576\,
            I => \N__25573\
        );

    \I__5623\ : CascadeBuf
    port map (
            O => \N__25573\,
            I => \N__25570\
        );

    \I__5622\ : CascadeMux
    port map (
            O => \N__25570\,
            I => \N__25567\
        );

    \I__5621\ : CascadeBuf
    port map (
            O => \N__25567\,
            I => \N__25564\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__25564\,
            I => \N__25561\
        );

    \I__5619\ : CascadeBuf
    port map (
            O => \N__25561\,
            I => \N__25558\
        );

    \I__5618\ : CascadeMux
    port map (
            O => \N__25558\,
            I => \N__25555\
        );

    \I__5617\ : CascadeBuf
    port map (
            O => \N__25555\,
            I => \N__25552\
        );

    \I__5616\ : CascadeMux
    port map (
            O => \N__25552\,
            I => \N__25549\
        );

    \I__5615\ : CascadeBuf
    port map (
            O => \N__25549\,
            I => \N__25546\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__25546\,
            I => \N__25543\
        );

    \I__5613\ : CascadeBuf
    port map (
            O => \N__25543\,
            I => \N__25540\
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__25540\,
            I => \N__25537\
        );

    \I__5611\ : CascadeBuf
    port map (
            O => \N__25537\,
            I => \N__25534\
        );

    \I__5610\ : CascadeMux
    port map (
            O => \N__25534\,
            I => \N__25531\
        );

    \I__5609\ : CascadeBuf
    port map (
            O => \N__25531\,
            I => \N__25528\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__25528\,
            I => \N__25525\
        );

    \I__5607\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25522\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__25522\,
            I => \N__25519\
        );

    \I__5605\ : Span4Mux_h
    port map (
            O => \N__25519\,
            I => \N__25515\
        );

    \I__5604\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25511\
        );

    \I__5603\ : Sp12to4
    port map (
            O => \N__25515\,
            I => \N__25508\
        );

    \I__5602\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25505\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__25511\,
            I => \N__25502\
        );

    \I__5600\ : Span12Mux_s6_v
    port map (
            O => \N__25508\,
            I => \N__25498\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__25505\,
            I => \N__25495\
        );

    \I__5598\ : Span4Mux_v
    port map (
            O => \N__25502\,
            I => \N__25492\
        );

    \I__5597\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25489\
        );

    \I__5596\ : Span12Mux_v
    port map (
            O => \N__25498\,
            I => \N__25486\
        );

    \I__5595\ : Odrv12
    port map (
            O => \N__25495\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5594\ : Odrv4
    port map (
            O => \N__25492\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__25489\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5592\ : Odrv12
    port map (
            O => \N__25486\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5591\ : CascadeMux
    port map (
            O => \N__25477\,
            I => \N_389_0_cascade_\
        );

    \I__5590\ : InMux
    port map (
            O => \N__25474\,
            I => \N__25471\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__25471\,
            I => \N__25468\
        );

    \I__5588\ : Span4Mux_h
    port map (
            O => \N__25468\,
            I => \N__25465\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__25465\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1\
        );

    \I__5586\ : InMux
    port map (
            O => \N__25462\,
            I => \N__25458\
        );

    \I__5585\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25455\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__25458\,
            I => \N__25452\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__25455\,
            I => \M_this_state_q_fastZ0Z_15\
        );

    \I__5582\ : Odrv12
    port map (
            O => \N__25452\,
            I => \M_this_state_q_fastZ0Z_15\
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__25447\,
            I => \N__25442\
        );

    \I__5580\ : InMux
    port map (
            O => \N__25446\,
            I => \N__25439\
        );

    \I__5579\ : InMux
    port map (
            O => \N__25445\,
            I => \N__25436\
        );

    \I__5578\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25433\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__25439\,
            I => \N__25428\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__25436\,
            I => \N__25428\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__25433\,
            I => \N__25425\
        );

    \I__5574\ : Span4Mux_v
    port map (
            O => \N__25428\,
            I => \N__25420\
        );

    \I__5573\ : Span4Mux_h
    port map (
            O => \N__25425\,
            I => \N__25417\
        );

    \I__5572\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25412\
        );

    \I__5571\ : InMux
    port map (
            O => \N__25423\,
            I => \N__25412\
        );

    \I__5570\ : Odrv4
    port map (
            O => \N__25420\,
            I => \N_297\
        );

    \I__5569\ : Odrv4
    port map (
            O => \N__25417\,
            I => \N_297\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__25412\,
            I => \N_297\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__25405\,
            I => \N__25402\
        );

    \I__5566\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25399\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__25399\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_9\
        );

    \I__5564\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25393\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__25393\,
            I => \N__25387\
        );

    \I__5562\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25384\
        );

    \I__5561\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25374\
        );

    \I__5560\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25374\
        );

    \I__5559\ : Span4Mux_h
    port map (
            O => \N__25387\,
            I => \N__25369\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__25384\,
            I => \N__25369\
        );

    \I__5557\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25364\
        );

    \I__5556\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25364\
        );

    \I__5555\ : CascadeMux
    port map (
            O => \N__25381\,
            I => \N__25361\
        );

    \I__5554\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25358\
        );

    \I__5553\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25355\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__25374\,
            I => \N__25348\
        );

    \I__5551\ : Span4Mux_v
    port map (
            O => \N__25369\,
            I => \N__25348\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__25364\,
            I => \N__25348\
        );

    \I__5549\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25345\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__25358\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__25355\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__25348\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__25345\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__25336\,
            I => \this_vga_signals.M_this_state_q_ns_0_a3_sxZ0Z_9_cascade_\
        );

    \I__5543\ : InMux
    port map (
            O => \N__25333\,
            I => \N__25327\
        );

    \I__5542\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25327\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__25327\,
            I => \N__25324\
        );

    \I__5540\ : Span4Mux_v
    port map (
            O => \N__25324\,
            I => \N__25321\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__25321\,
            I => \N__25318\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__25318\,
            I => \N__25315\
        );

    \I__5537\ : Span4Mux_h
    port map (
            O => \N__25315\,
            I => \N__25312\
        );

    \I__5536\ : Odrv4
    port map (
            O => \N__25312\,
            I => port_address_in_4
        );

    \I__5535\ : InMux
    port map (
            O => \N__25309\,
            I => \N__25305\
        );

    \I__5534\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25302\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__25305\,
            I => \N__25299\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__25302\,
            I => \N__25296\
        );

    \I__5531\ : Span4Mux_h
    port map (
            O => \N__25299\,
            I => \N__25291\
        );

    \I__5530\ : Span4Mux_h
    port map (
            O => \N__25296\,
            I => \N__25291\
        );

    \I__5529\ : Span4Mux_v
    port map (
            O => \N__25291\,
            I => \N__25288\
        );

    \I__5528\ : Sp12to4
    port map (
            O => \N__25288\,
            I => \N__25284\
        );

    \I__5527\ : InMux
    port map (
            O => \N__25287\,
            I => \N__25281\
        );

    \I__5526\ : Span12Mux_h
    port map (
            O => \N__25284\,
            I => \N__25278\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__25281\,
            I => \N__25275\
        );

    \I__5524\ : Odrv12
    port map (
            O => \N__25278\,
            I => port_rw_in
        );

    \I__5523\ : Odrv12
    port map (
            O => \N__25275\,
            I => port_rw_in
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__25270\,
            I => \N__25266\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__25269\,
            I => \N__25263\
        );

    \I__5520\ : InMux
    port map (
            O => \N__25266\,
            I => \N__25258\
        );

    \I__5519\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25258\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__25258\,
            I => \N__25255\
        );

    \I__5517\ : Span12Mux_h
    port map (
            O => \N__25255\,
            I => \N__25252\
        );

    \I__5516\ : Span12Mux_v
    port map (
            O => \N__25252\,
            I => \N__25249\
        );

    \I__5515\ : Odrv12
    port map (
            O => \N__25249\,
            I => port_address_in_7
        );

    \I__5514\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25243\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__25243\,
            I => \un1_M_this_map_address_q_cry_6_c_RNII22SZ0\
        );

    \I__5512\ : InMux
    port map (
            O => \N__25240\,
            I => \un1_M_this_map_address_q_cry_6\
        );

    \I__5511\ : InMux
    port map (
            O => \N__25237\,
            I => \bfn_19_23_0_\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__25234\,
            I => \N__25231\
        );

    \I__5509\ : CascadeBuf
    port map (
            O => \N__25231\,
            I => \N__25228\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__25228\,
            I => \N__25225\
        );

    \I__5507\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25222\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__25222\,
            I => \N__25219\
        );

    \I__5505\ : Span4Mux_h
    port map (
            O => \N__25219\,
            I => \N__25215\
        );

    \I__5504\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25211\
        );

    \I__5503\ : Sp12to4
    port map (
            O => \N__25215\,
            I => \N__25207\
        );

    \I__5502\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25204\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__25211\,
            I => \N__25201\
        );

    \I__5500\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25198\
        );

    \I__5499\ : Span12Mux_s9_v
    port map (
            O => \N__25207\,
            I => \N__25195\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__25204\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__5497\ : Odrv12
    port map (
            O => \N__25201\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__25198\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__5495\ : Odrv12
    port map (
            O => \N__25195\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__5494\ : InMux
    port map (
            O => \N__25186\,
            I => \un1_M_this_map_address_q_cry_8\
        );

    \I__5493\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25180\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__25180\,
            I => \un1_M_this_map_address_q_cry_8_c_RNIM84SZ0\
        );

    \I__5491\ : InMux
    port map (
            O => \N__25177\,
            I => \N__25174\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__25174\,
            I => \this_vga_signals.M_this_map_address_d_5_mZ0Z_7\
        );

    \I__5489\ : CascadeMux
    port map (
            O => \N__25171\,
            I => \N__25168\
        );

    \I__5488\ : CascadeBuf
    port map (
            O => \N__25168\,
            I => \N__25165\
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__25165\,
            I => \N__25162\
        );

    \I__5486\ : InMux
    port map (
            O => \N__25162\,
            I => \N__25158\
        );

    \I__5485\ : CascadeMux
    port map (
            O => \N__25161\,
            I => \N__25153\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__25158\,
            I => \N__25150\
        );

    \I__5483\ : InMux
    port map (
            O => \N__25157\,
            I => \N__25147\
        );

    \I__5482\ : InMux
    port map (
            O => \N__25156\,
            I => \N__25144\
        );

    \I__5481\ : InMux
    port map (
            O => \N__25153\,
            I => \N__25141\
        );

    \I__5480\ : Span12Mux_s9_v
    port map (
            O => \N__25150\,
            I => \N__25138\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__25147\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__25144\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__25141\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__5476\ : Odrv12
    port map (
            O => \N__25138\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__5475\ : CascadeMux
    port map (
            O => \N__25129\,
            I => \N__25126\
        );

    \I__5474\ : InMux
    port map (
            O => \N__25126\,
            I => \N__25123\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__25123\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_7\
        );

    \I__5472\ : CascadeMux
    port map (
            O => \N__25120\,
            I => \N__25117\
        );

    \I__5471\ : CascadeBuf
    port map (
            O => \N__25117\,
            I => \N__25113\
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__25116\,
            I => \N__25110\
        );

    \I__5469\ : CascadeMux
    port map (
            O => \N__25113\,
            I => \N__25107\
        );

    \I__5468\ : InMux
    port map (
            O => \N__25110\,
            I => \N__25104\
        );

    \I__5467\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25101\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__25104\,
            I => \N__25098\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__25101\,
            I => \N__25094\
        );

    \I__5464\ : Span4Mux_h
    port map (
            O => \N__25098\,
            I => \N__25090\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__25097\,
            I => \N__25087\
        );

    \I__5462\ : Span4Mux_s2_v
    port map (
            O => \N__25094\,
            I => \N__25084\
        );

    \I__5461\ : CascadeMux
    port map (
            O => \N__25093\,
            I => \N__25081\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__25090\,
            I => \N__25077\
        );

    \I__5459\ : InMux
    port map (
            O => \N__25087\,
            I => \N__25074\
        );

    \I__5458\ : Span4Mux_h
    port map (
            O => \N__25084\,
            I => \N__25071\
        );

    \I__5457\ : InMux
    port map (
            O => \N__25081\,
            I => \N__25066\
        );

    \I__5456\ : InMux
    port map (
            O => \N__25080\,
            I => \N__25066\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__25077\,
            I => \N__25063\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__25074\,
            I => \N__25058\
        );

    \I__5453\ : Span4Mux_v
    port map (
            O => \N__25071\,
            I => \N__25058\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__25066\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__25063\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__5450\ : Odrv4
    port map (
            O => \N__25058\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__5449\ : InMux
    port map (
            O => \N__25051\,
            I => \N__25046\
        );

    \I__5448\ : InMux
    port map (
            O => \N__25050\,
            I => \N__25041\
        );

    \I__5447\ : InMux
    port map (
            O => \N__25049\,
            I => \N__25041\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__25046\,
            I => \this_ppu.un1_M_haddress_q_c5\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__25041\,
            I => \this_ppu.un1_M_haddress_q_c5\
        );

    \I__5444\ : SRMux
    port map (
            O => \N__25036\,
            I => \N__25031\
        );

    \I__5443\ : SRMux
    port map (
            O => \N__25035\,
            I => \N__25027\
        );

    \I__5442\ : SRMux
    port map (
            O => \N__25034\,
            I => \N__25024\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__25031\,
            I => \N__25021\
        );

    \I__5440\ : SRMux
    port map (
            O => \N__25030\,
            I => \N__25018\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__25027\,
            I => \N__25015\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__25024\,
            I => \N__25012\
        );

    \I__5437\ : Span4Mux_v
    port map (
            O => \N__25021\,
            I => \N__25007\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__25018\,
            I => \N__25007\
        );

    \I__5435\ : Span4Mux_h
    port map (
            O => \N__25015\,
            I => \N__25004\
        );

    \I__5434\ : Span4Mux_h
    port map (
            O => \N__25012\,
            I => \N__25001\
        );

    \I__5433\ : Span4Mux_v
    port map (
            O => \N__25007\,
            I => \N__24998\
        );

    \I__5432\ : Odrv4
    port map (
            O => \N__25004\,
            I => \this_ppu.M_last_q_RNI21NK5\
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__25001\,
            I => \this_ppu.M_last_q_RNI21NK5\
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__24998\,
            I => \this_ppu.M_last_q_RNI21NK5\
        );

    \I__5429\ : InMux
    port map (
            O => \N__24991\,
            I => \N__24988\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__24988\,
            I => \N__24985\
        );

    \I__5427\ : Odrv12
    port map (
            O => \N__24985\,
            I => \this_reset_cond.M_stage_qZ0Z_6\
        );

    \I__5426\ : InMux
    port map (
            O => \N__24982\,
            I => \N__24979\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__24979\,
            I => \N__24976\
        );

    \I__5424\ : Odrv12
    port map (
            O => \N__24976\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__24973\,
            I => \N__24970\
        );

    \I__5422\ : CascadeBuf
    port map (
            O => \N__24970\,
            I => \N__24967\
        );

    \I__5421\ : CascadeMux
    port map (
            O => \N__24967\,
            I => \N__24964\
        );

    \I__5420\ : CascadeBuf
    port map (
            O => \N__24964\,
            I => \N__24961\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__24961\,
            I => \N__24958\
        );

    \I__5418\ : CascadeBuf
    port map (
            O => \N__24958\,
            I => \N__24955\
        );

    \I__5417\ : CascadeMux
    port map (
            O => \N__24955\,
            I => \N__24952\
        );

    \I__5416\ : CascadeBuf
    port map (
            O => \N__24952\,
            I => \N__24949\
        );

    \I__5415\ : CascadeMux
    port map (
            O => \N__24949\,
            I => \N__24946\
        );

    \I__5414\ : CascadeBuf
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__5413\ : CascadeMux
    port map (
            O => \N__24943\,
            I => \N__24940\
        );

    \I__5412\ : CascadeBuf
    port map (
            O => \N__24940\,
            I => \N__24937\
        );

    \I__5411\ : CascadeMux
    port map (
            O => \N__24937\,
            I => \N__24934\
        );

    \I__5410\ : CascadeBuf
    port map (
            O => \N__24934\,
            I => \N__24931\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__24931\,
            I => \N__24928\
        );

    \I__5408\ : CascadeBuf
    port map (
            O => \N__24928\,
            I => \N__24925\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__24925\,
            I => \N__24922\
        );

    \I__5406\ : CascadeBuf
    port map (
            O => \N__24922\,
            I => \N__24919\
        );

    \I__5405\ : CascadeMux
    port map (
            O => \N__24919\,
            I => \N__24916\
        );

    \I__5404\ : CascadeBuf
    port map (
            O => \N__24916\,
            I => \N__24913\
        );

    \I__5403\ : CascadeMux
    port map (
            O => \N__24913\,
            I => \N__24910\
        );

    \I__5402\ : CascadeBuf
    port map (
            O => \N__24910\,
            I => \N__24907\
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__24907\,
            I => \N__24904\
        );

    \I__5400\ : CascadeBuf
    port map (
            O => \N__24904\,
            I => \N__24901\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__24901\,
            I => \N__24898\
        );

    \I__5398\ : CascadeBuf
    port map (
            O => \N__24898\,
            I => \N__24895\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__24895\,
            I => \N__24892\
        );

    \I__5396\ : CascadeBuf
    port map (
            O => \N__24892\,
            I => \N__24889\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__24889\,
            I => \N__24886\
        );

    \I__5394\ : CascadeBuf
    port map (
            O => \N__24886\,
            I => \N__24883\
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__24883\,
            I => \N__24880\
        );

    \I__5392\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24877\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__24877\,
            I => \N__24874\
        );

    \I__5390\ : Span4Mux_s1_v
    port map (
            O => \N__24874\,
            I => \N__24870\
        );

    \I__5389\ : CascadeMux
    port map (
            O => \N__24873\,
            I => \N__24867\
        );

    \I__5388\ : Sp12to4
    port map (
            O => \N__24870\,
            I => \N__24863\
        );

    \I__5387\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24860\
        );

    \I__5386\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24856\
        );

    \I__5385\ : Span12Mux_s5_v
    port map (
            O => \N__24863\,
            I => \N__24853\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__24860\,
            I => \N__24850\
        );

    \I__5383\ : InMux
    port map (
            O => \N__24859\,
            I => \N__24847\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__24856\,
            I => \N__24842\
        );

    \I__5381\ : Span12Mux_v
    port map (
            O => \N__24853\,
            I => \N__24842\
        );

    \I__5380\ : Odrv4
    port map (
            O => \N__24850\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__24847\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__5378\ : Odrv12
    port map (
            O => \N__24842\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__5377\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24832\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__24832\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5\
        );

    \I__5375\ : InMux
    port map (
            O => \N__24829\,
            I => \N__24826\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24823\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__24823\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_6\
        );

    \I__5372\ : CascadeMux
    port map (
            O => \N__24820\,
            I => \this_vga_signals.M_this_map_address_d_5_mZ0Z_6_cascade_\
        );

    \I__5371\ : InMux
    port map (
            O => \N__24817\,
            I => \N__24814\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__24814\,
            I => \M_this_map_address_q_RNICF7V6Z0Z_0\
        );

    \I__5369\ : InMux
    port map (
            O => \N__24811\,
            I => \un1_M_this_map_address_q_cry_0\
        );

    \I__5368\ : CascadeMux
    port map (
            O => \N__24808\,
            I => \N__24805\
        );

    \I__5367\ : CascadeBuf
    port map (
            O => \N__24805\,
            I => \N__24802\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__24802\,
            I => \N__24799\
        );

    \I__5365\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24796\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__24796\,
            I => \N__24793\
        );

    \I__5363\ : Span4Mux_s2_v
    port map (
            O => \N__24793\,
            I => \N__24790\
        );

    \I__5362\ : Span4Mux_h
    port map (
            O => \N__24790\,
            I => \N__24787\
        );

    \I__5361\ : Span4Mux_h
    port map (
            O => \N__24787\,
            I => \N__24781\
        );

    \I__5360\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24776\
        );

    \I__5359\ : InMux
    port map (
            O => \N__24785\,
            I => \N__24776\
        );

    \I__5358\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24773\
        );

    \I__5357\ : Span4Mux_v
    port map (
            O => \N__24781\,
            I => \N__24770\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__24776\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__24773\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__5354\ : Odrv4
    port map (
            O => \N__24770\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__5353\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24760\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__24760\,
            I => \un1_M_this_map_address_q_cry_1_c_RNI8JSRZ0\
        );

    \I__5351\ : InMux
    port map (
            O => \N__24757\,
            I => \un1_M_this_map_address_q_cry_1\
        );

    \I__5350\ : InMux
    port map (
            O => \N__24754\,
            I => \un1_M_this_map_address_q_cry_2\
        );

    \I__5349\ : InMux
    port map (
            O => \N__24751\,
            I => \un1_M_this_map_address_q_cry_3\
        );

    \I__5348\ : CascadeMux
    port map (
            O => \N__24748\,
            I => \N__24745\
        );

    \I__5347\ : CascadeBuf
    port map (
            O => \N__24745\,
            I => \N__24742\
        );

    \I__5346\ : CascadeMux
    port map (
            O => \N__24742\,
            I => \N__24739\
        );

    \I__5345\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24736\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__24736\,
            I => \N__24733\
        );

    \I__5343\ : Sp12to4
    port map (
            O => \N__24733\,
            I => \N__24727\
        );

    \I__5342\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24724\
        );

    \I__5341\ : InMux
    port map (
            O => \N__24731\,
            I => \N__24721\
        );

    \I__5340\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24718\
        );

    \I__5339\ : Span12Mux_s11_v
    port map (
            O => \N__24727\,
            I => \N__24715\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__24724\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__24721\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__24718\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__5335\ : Odrv12
    port map (
            O => \N__24715\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__5334\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24703\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__24703\,
            I => \un1_M_this_map_address_q_cry_4_c_RNIESVRZ0\
        );

    \I__5332\ : InMux
    port map (
            O => \N__24700\,
            I => \un1_M_this_map_address_q_cry_4\
        );

    \I__5331\ : CascadeMux
    port map (
            O => \N__24697\,
            I => \N__24694\
        );

    \I__5330\ : CascadeBuf
    port map (
            O => \N__24694\,
            I => \N__24691\
        );

    \I__5329\ : CascadeMux
    port map (
            O => \N__24691\,
            I => \N__24688\
        );

    \I__5328\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24685\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__24685\,
            I => \N__24682\
        );

    \I__5326\ : Span4Mux_v
    port map (
            O => \N__24682\,
            I => \N__24679\
        );

    \I__5325\ : Sp12to4
    port map (
            O => \N__24679\,
            I => \N__24673\
        );

    \I__5324\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24670\
        );

    \I__5323\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24667\
        );

    \I__5322\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24664\
        );

    \I__5321\ : Span12Mux_h
    port map (
            O => \N__24673\,
            I => \N__24661\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__24670\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__24667\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__24664\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__5317\ : Odrv12
    port map (
            O => \N__24661\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__5316\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24649\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__24649\,
            I => \un1_M_this_map_address_q_cry_5_c_RNIGV0SZ0\
        );

    \I__5314\ : InMux
    port map (
            O => \N__24646\,
            I => \un1_M_this_map_address_q_cry_5\
        );

    \I__5313\ : CascadeMux
    port map (
            O => \N__24643\,
            I => \this_vga_signals.M_this_state_d_1_sqmuxaZ0_cascade_\
        );

    \I__5312\ : CascadeMux
    port map (
            O => \N__24640\,
            I => \N__24637\
        );

    \I__5311\ : InMux
    port map (
            O => \N__24637\,
            I => \N__24634\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__24634\,
            I => \N__24631\
        );

    \I__5309\ : Span4Mux_v
    port map (
            O => \N__24631\,
            I => \N__24628\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__24628\,
            I => \this_vga_signals.N_399_0\
        );

    \I__5307\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24622\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__24622\,
            I => \this_vga_signals.M_this_map_address_d_5_mZ0Z_5\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__24619\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_5_cascade_\
        );

    \I__5304\ : CascadeMux
    port map (
            O => \N__24616\,
            I => \N__24613\
        );

    \I__5303\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24610\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__24610\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_0\
        );

    \I__5301\ : CascadeMux
    port map (
            O => \N__24607\,
            I => \N__24604\
        );

    \I__5300\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24601\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__24601\,
            I => \N__24598\
        );

    \I__5298\ : Odrv4
    port map (
            O => \N__24598\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_11\
        );

    \I__5297\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24591\
        );

    \I__5296\ : InMux
    port map (
            O => \N__24594\,
            I => \N__24588\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__24591\,
            I => \N__24585\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24582\
        );

    \I__5293\ : Odrv12
    port map (
            O => \N__24585\,
            I => \this_vga_signals.N_446_1\
        );

    \I__5292\ : Odrv4
    port map (
            O => \N__24582\,
            I => \this_vga_signals.N_446_1\
        );

    \I__5291\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24572\
        );

    \I__5290\ : InMux
    port map (
            O => \N__24576\,
            I => \N__24569\
        );

    \I__5289\ : CascadeMux
    port map (
            O => \N__24575\,
            I => \N__24563\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__24572\,
            I => \N__24556\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__24569\,
            I => \N__24556\
        );

    \I__5286\ : InMux
    port map (
            O => \N__24568\,
            I => \N__24553\
        );

    \I__5285\ : InMux
    port map (
            O => \N__24567\,
            I => \N__24550\
        );

    \I__5284\ : InMux
    port map (
            O => \N__24566\,
            I => \N__24543\
        );

    \I__5283\ : InMux
    port map (
            O => \N__24563\,
            I => \N__24543\
        );

    \I__5282\ : InMux
    port map (
            O => \N__24562\,
            I => \N__24543\
        );

    \I__5281\ : InMux
    port map (
            O => \N__24561\,
            I => \N__24540\
        );

    \I__5280\ : Span4Mux_h
    port map (
            O => \N__24556\,
            I => \N__24537\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__24553\,
            I => \N__24532\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__24550\,
            I => \N__24532\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__24543\,
            I => \N__24529\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__24540\,
            I => \N__24526\
        );

    \I__5275\ : Span4Mux_h
    port map (
            O => \N__24537\,
            I => \N__24520\
        );

    \I__5274\ : Span12Mux_h
    port map (
            O => \N__24532\,
            I => \N__24517\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__24529\,
            I => \N__24514\
        );

    \I__5272\ : Span4Mux_h
    port map (
            O => \N__24526\,
            I => \N__24511\
        );

    \I__5271\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24508\
        );

    \I__5270\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24505\
        );

    \I__5269\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24502\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__24520\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5267\ : Odrv12
    port map (
            O => \N__24517\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5266\ : Odrv4
    port map (
            O => \N__24514\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__24511\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__24508\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__24505\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__24502\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5261\ : InMux
    port map (
            O => \N__24487\,
            I => \N__24484\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__24484\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11\
        );

    \I__5259\ : CascadeMux
    port map (
            O => \N__24481\,
            I => \N__24477\
        );

    \I__5258\ : InMux
    port map (
            O => \N__24480\,
            I => \N__24470\
        );

    \I__5257\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24462\
        );

    \I__5256\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24459\
        );

    \I__5255\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24456\
        );

    \I__5254\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24449\
        );

    \I__5253\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24449\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__24470\,
            I => \N__24446\
        );

    \I__5251\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24443\
        );

    \I__5250\ : InMux
    port map (
            O => \N__24468\,
            I => \N__24440\
        );

    \I__5249\ : CascadeMux
    port map (
            O => \N__24467\,
            I => \N__24437\
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__24466\,
            I => \N__24432\
        );

    \I__5247\ : InMux
    port map (
            O => \N__24465\,
            I => \N__24428\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__24462\,
            I => \N__24423\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__24459\,
            I => \N__24423\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24420\
        );

    \I__5243\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24414\
        );

    \I__5242\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24414\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__24449\,
            I => \N__24407\
        );

    \I__5240\ : Span4Mux_h
    port map (
            O => \N__24446\,
            I => \N__24407\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__24443\,
            I => \N__24407\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__24440\,
            I => \N__24404\
        );

    \I__5237\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24400\
        );

    \I__5236\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24397\
        );

    \I__5235\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24390\
        );

    \I__5234\ : InMux
    port map (
            O => \N__24432\,
            I => \N__24390\
        );

    \I__5233\ : InMux
    port map (
            O => \N__24431\,
            I => \N__24390\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__24428\,
            I => \N__24387\
        );

    \I__5231\ : Span4Mux_h
    port map (
            O => \N__24423\,
            I => \N__24382\
        );

    \I__5230\ : Span4Mux_h
    port map (
            O => \N__24420\,
            I => \N__24382\
        );

    \I__5229\ : InMux
    port map (
            O => \N__24419\,
            I => \N__24379\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__24414\,
            I => \N__24372\
        );

    \I__5227\ : Span4Mux_v
    port map (
            O => \N__24407\,
            I => \N__24372\
        );

    \I__5226\ : Span4Mux_h
    port map (
            O => \N__24404\,
            I => \N__24372\
        );

    \I__5225\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24369\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__24400\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__24397\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__24390\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5221\ : Odrv4
    port map (
            O => \N__24387\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5220\ : Odrv4
    port map (
            O => \N__24382\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__24379\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5218\ : Odrv4
    port map (
            O => \N__24372\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__24369\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__24352\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_\
        );

    \I__5215\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24346\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__24346\,
            I => \N__24343\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__24343\,
            I => \un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__24340\,
            I => \N__24337\
        );

    \I__5211\ : CascadeBuf
    port map (
            O => \N__24337\,
            I => \N__24334\
        );

    \I__5210\ : CascadeMux
    port map (
            O => \N__24334\,
            I => \N__24331\
        );

    \I__5209\ : CascadeBuf
    port map (
            O => \N__24331\,
            I => \N__24328\
        );

    \I__5208\ : CascadeMux
    port map (
            O => \N__24328\,
            I => \N__24325\
        );

    \I__5207\ : CascadeBuf
    port map (
            O => \N__24325\,
            I => \N__24322\
        );

    \I__5206\ : CascadeMux
    port map (
            O => \N__24322\,
            I => \N__24319\
        );

    \I__5205\ : CascadeBuf
    port map (
            O => \N__24319\,
            I => \N__24316\
        );

    \I__5204\ : CascadeMux
    port map (
            O => \N__24316\,
            I => \N__24313\
        );

    \I__5203\ : CascadeBuf
    port map (
            O => \N__24313\,
            I => \N__24310\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__24310\,
            I => \N__24307\
        );

    \I__5201\ : CascadeBuf
    port map (
            O => \N__24307\,
            I => \N__24304\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__24304\,
            I => \N__24301\
        );

    \I__5199\ : CascadeBuf
    port map (
            O => \N__24301\,
            I => \N__24298\
        );

    \I__5198\ : CascadeMux
    port map (
            O => \N__24298\,
            I => \N__24295\
        );

    \I__5197\ : CascadeBuf
    port map (
            O => \N__24295\,
            I => \N__24292\
        );

    \I__5196\ : CascadeMux
    port map (
            O => \N__24292\,
            I => \N__24289\
        );

    \I__5195\ : CascadeBuf
    port map (
            O => \N__24289\,
            I => \N__24286\
        );

    \I__5194\ : CascadeMux
    port map (
            O => \N__24286\,
            I => \N__24283\
        );

    \I__5193\ : CascadeBuf
    port map (
            O => \N__24283\,
            I => \N__24280\
        );

    \I__5192\ : CascadeMux
    port map (
            O => \N__24280\,
            I => \N__24277\
        );

    \I__5191\ : CascadeBuf
    port map (
            O => \N__24277\,
            I => \N__24274\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__24274\,
            I => \N__24271\
        );

    \I__5189\ : CascadeBuf
    port map (
            O => \N__24271\,
            I => \N__24268\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__24268\,
            I => \N__24265\
        );

    \I__5187\ : CascadeBuf
    port map (
            O => \N__24265\,
            I => \N__24262\
        );

    \I__5186\ : CascadeMux
    port map (
            O => \N__24262\,
            I => \N__24259\
        );

    \I__5185\ : CascadeBuf
    port map (
            O => \N__24259\,
            I => \N__24256\
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__24256\,
            I => \N__24253\
        );

    \I__5183\ : CascadeBuf
    port map (
            O => \N__24253\,
            I => \N__24250\
        );

    \I__5182\ : CascadeMux
    port map (
            O => \N__24250\,
            I => \N__24247\
        );

    \I__5181\ : InMux
    port map (
            O => \N__24247\,
            I => \N__24244\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__24244\,
            I => \N__24241\
        );

    \I__5179\ : Span4Mux_h
    port map (
            O => \N__24241\,
            I => \N__24237\
        );

    \I__5178\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24234\
        );

    \I__5177\ : Sp12to4
    port map (
            O => \N__24237\,
            I => \N__24229\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__24234\,
            I => \N__24226\
        );

    \I__5175\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24221\
        );

    \I__5174\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24221\
        );

    \I__5173\ : Span12Mux_v
    port map (
            O => \N__24229\,
            I => \N__24218\
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__24226\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__24221\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5170\ : Odrv12
    port map (
            O => \N__24218\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5169\ : InMux
    port map (
            O => \N__24211\,
            I => \N__24208\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__24208\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_7\
        );

    \I__5167\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24202\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__24202\,
            I => \N__24199\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__24199\,
            I => \un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__24196\,
            I => \N__24193\
        );

    \I__5163\ : InMux
    port map (
            O => \N__24193\,
            I => \N__24190\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__24190\,
            I => \N__24187\
        );

    \I__5161\ : Span4Mux_h
    port map (
            O => \N__24187\,
            I => \N__24184\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__24184\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_4\
        );

    \I__5159\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24176\
        );

    \I__5158\ : InMux
    port map (
            O => \N__24180\,
            I => \N__24165\
        );

    \I__5157\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24165\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24162\
        );

    \I__5155\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24159\
        );

    \I__5154\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24152\
        );

    \I__5153\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24152\
        );

    \I__5152\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24152\
        );

    \I__5151\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24144\
        );

    \I__5150\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24144\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__24165\,
            I => \N__24139\
        );

    \I__5148\ : Span4Mux_v
    port map (
            O => \N__24162\,
            I => \N__24132\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__24159\,
            I => \N__24132\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__24152\,
            I => \N__24132\
        );

    \I__5145\ : InMux
    port map (
            O => \N__24151\,
            I => \N__24129\
        );

    \I__5144\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24124\
        );

    \I__5143\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24124\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__24144\,
            I => \N__24121\
        );

    \I__5141\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24116\
        );

    \I__5140\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24116\
        );

    \I__5139\ : Odrv4
    port map (
            O => \N__24139\,
            I => \this_vga_signals.un1_M_this_state_q_19_0\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__24132\,
            I => \this_vga_signals.un1_M_this_state_q_19_0\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__24129\,
            I => \this_vga_signals.un1_M_this_state_q_19_0\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__24124\,
            I => \this_vga_signals.un1_M_this_state_q_19_0\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__24121\,
            I => \this_vga_signals.un1_M_this_state_q_19_0\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__24116\,
            I => \this_vga_signals.un1_M_this_state_q_19_0\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__24103\,
            I => \this_vga_signals.N_294_cascade_\
        );

    \I__5132\ : CascadeMux
    port map (
            O => \N__24100\,
            I => \this_vga_signals.un1_M_this_state_q_14Z0Z_1_cascade_\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__24097\,
            I => \N__24092\
        );

    \I__5130\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24089\
        );

    \I__5129\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24086\
        );

    \I__5128\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24083\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__24089\,
            I => \un1_M_this_state_q_14_0\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__24086\,
            I => \un1_M_this_state_q_14_0\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__24083\,
            I => \un1_M_this_state_q_14_0\
        );

    \I__5124\ : CascadeMux
    port map (
            O => \N__24076\,
            I => \N__24073\
        );

    \I__5123\ : InMux
    port map (
            O => \N__24073\,
            I => \N__24069\
        );

    \I__5122\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24066\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__24069\,
            I => this_vga_signals_un23_i_a2_1_1
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__24066\,
            I => this_vga_signals_un23_i_a2_1_1
        );

    \I__5119\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24058\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__24058\,
            I => \N__24055\
        );

    \I__5117\ : Odrv4
    port map (
            O => \N__24055\,
            I => un23_i_a2_1
        );

    \I__5116\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24049\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__24049\,
            I => \N__24046\
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__24046\,
            I => \this_vga_signals.N_486\
        );

    \I__5113\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24039\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__24042\,
            I => \N__24036\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__24039\,
            I => \N__24033\
        );

    \I__5110\ : InMux
    port map (
            O => \N__24036\,
            I => \N__24030\
        );

    \I__5109\ : Span4Mux_v
    port map (
            O => \N__24033\,
            I => \N__24027\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__24030\,
            I => \N__24024\
        );

    \I__5107\ : Odrv4
    port map (
            O => \N__24027\,
            I => \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_5\
        );

    \I__5106\ : Odrv4
    port map (
            O => \N__24024\,
            I => \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_5\
        );

    \I__5105\ : CascadeMux
    port map (
            O => \N__24019\,
            I => \this_vga_signals.N_486_cascade_\
        );

    \I__5104\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24013\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__24013\,
            I => \N__24009\
        );

    \I__5102\ : InMux
    port map (
            O => \N__24012\,
            I => \N__24006\
        );

    \I__5101\ : Span4Mux_v
    port map (
            O => \N__24009\,
            I => \N__24001\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__24006\,
            I => \N__24001\
        );

    \I__5099\ : Span4Mux_v
    port map (
            O => \N__24001\,
            I => \N__23998\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__23998\,
            I => \this_vga_signals.N_438_1\
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__23995\,
            I => \N__23992\
        );

    \I__5096\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23989\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__23989\,
            I => \N__23986\
        );

    \I__5094\ : Odrv12
    port map (
            O => \N__23986\,
            I => \this_vga_signals_M_this_state_q_ns_i_o2_0_12\
        );

    \I__5093\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23977\
        );

    \I__5092\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23977\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__23977\,
            I => \N__23972\
        );

    \I__5090\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23969\
        );

    \I__5089\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23966\
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__23972\,
            I => \this_ppu.un1_M_haddress_q_c2\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__23969\,
            I => \this_ppu.un1_M_haddress_q_c2\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__23966\,
            I => \this_ppu.un1_M_haddress_q_c2\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__23959\,
            I => \N__23955\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__23958\,
            I => \N__23952\
        );

    \I__5083\ : CascadeBuf
    port map (
            O => \N__23955\,
            I => \N__23949\
        );

    \I__5082\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23946\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__23949\,
            I => \N__23943\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__23946\,
            I => \N__23940\
        );

    \I__5079\ : InMux
    port map (
            O => \N__23943\,
            I => \N__23937\
        );

    \I__5078\ : Span4Mux_h
    port map (
            O => \N__23940\,
            I => \N__23934\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__23937\,
            I => \N__23931\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__23934\,
            I => \N__23927\
        );

    \I__5075\ : Span4Mux_s2_v
    port map (
            O => \N__23931\,
            I => \N__23924\
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__23930\,
            I => \N__23921\
        );

    \I__5073\ : Span4Mux_v
    port map (
            O => \N__23927\,
            I => \N__23916\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__23924\,
            I => \N__23913\
        );

    \I__5071\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23908\
        );

    \I__5070\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23908\
        );

    \I__5069\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23905\
        );

    \I__5068\ : Span4Mux_h
    port map (
            O => \N__23916\,
            I => \N__23900\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__23913\,
            I => \N__23900\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__23908\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__23905\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__23900\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__5063\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23890\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__23890\,
            I => \N__23887\
        );

    \I__5061\ : Span4Mux_v
    port map (
            O => \N__23887\,
            I => \N__23882\
        );

    \I__5060\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23878\
        );

    \I__5059\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23875\
        );

    \I__5058\ : Span4Mux_h
    port map (
            O => \N__23882\,
            I => \N__23872\
        );

    \I__5057\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23869\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__23878\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__23875\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__5054\ : Odrv4
    port map (
            O => \N__23872\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__23869\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__5052\ : CascadeMux
    port map (
            O => \N__23860\,
            I => \N__23857\
        );

    \I__5051\ : CascadeBuf
    port map (
            O => \N__23857\,
            I => \N__23854\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__23854\,
            I => \N__23851\
        );

    \I__5049\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23848\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__23848\,
            I => \N__23845\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__23845\,
            I => \N__23842\
        );

    \I__5046\ : Span4Mux_h
    port map (
            O => \N__23842\,
            I => \N__23839\
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__23839\,
            I => \this_ppu_M_vaddress_q_i_6\
        );

    \I__5044\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23833\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__23833\,
            I => \N__23830\
        );

    \I__5042\ : Span4Mux_h
    port map (
            O => \N__23830\,
            I => \N__23827\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__23827\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_6\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__23824\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6_cascade_\
        );

    \I__5039\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23818\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__23818\,
            I => \N__23815\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__23815\,
            I => \un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0\
        );

    \I__5036\ : CascadeMux
    port map (
            O => \N__23812\,
            I => \N__23809\
        );

    \I__5035\ : CascadeBuf
    port map (
            O => \N__23809\,
            I => \N__23806\
        );

    \I__5034\ : CascadeMux
    port map (
            O => \N__23806\,
            I => \N__23803\
        );

    \I__5033\ : CascadeBuf
    port map (
            O => \N__23803\,
            I => \N__23800\
        );

    \I__5032\ : CascadeMux
    port map (
            O => \N__23800\,
            I => \N__23797\
        );

    \I__5031\ : CascadeBuf
    port map (
            O => \N__23797\,
            I => \N__23794\
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__23794\,
            I => \N__23791\
        );

    \I__5029\ : CascadeBuf
    port map (
            O => \N__23791\,
            I => \N__23788\
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__23788\,
            I => \N__23785\
        );

    \I__5027\ : CascadeBuf
    port map (
            O => \N__23785\,
            I => \N__23782\
        );

    \I__5026\ : CascadeMux
    port map (
            O => \N__23782\,
            I => \N__23779\
        );

    \I__5025\ : CascadeBuf
    port map (
            O => \N__23779\,
            I => \N__23776\
        );

    \I__5024\ : CascadeMux
    port map (
            O => \N__23776\,
            I => \N__23773\
        );

    \I__5023\ : CascadeBuf
    port map (
            O => \N__23773\,
            I => \N__23770\
        );

    \I__5022\ : CascadeMux
    port map (
            O => \N__23770\,
            I => \N__23767\
        );

    \I__5021\ : CascadeBuf
    port map (
            O => \N__23767\,
            I => \N__23764\
        );

    \I__5020\ : CascadeMux
    port map (
            O => \N__23764\,
            I => \N__23761\
        );

    \I__5019\ : CascadeBuf
    port map (
            O => \N__23761\,
            I => \N__23758\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__23758\,
            I => \N__23755\
        );

    \I__5017\ : CascadeBuf
    port map (
            O => \N__23755\,
            I => \N__23752\
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__23752\,
            I => \N__23749\
        );

    \I__5015\ : CascadeBuf
    port map (
            O => \N__23749\,
            I => \N__23746\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__23746\,
            I => \N__23743\
        );

    \I__5013\ : CascadeBuf
    port map (
            O => \N__23743\,
            I => \N__23740\
        );

    \I__5012\ : CascadeMux
    port map (
            O => \N__23740\,
            I => \N__23737\
        );

    \I__5011\ : CascadeBuf
    port map (
            O => \N__23737\,
            I => \N__23734\
        );

    \I__5010\ : CascadeMux
    port map (
            O => \N__23734\,
            I => \N__23731\
        );

    \I__5009\ : CascadeBuf
    port map (
            O => \N__23731\,
            I => \N__23728\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__23728\,
            I => \N__23725\
        );

    \I__5007\ : CascadeBuf
    port map (
            O => \N__23725\,
            I => \N__23722\
        );

    \I__5006\ : CascadeMux
    port map (
            O => \N__23722\,
            I => \N__23719\
        );

    \I__5005\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23716\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__23716\,
            I => \N__23713\
        );

    \I__5003\ : Span4Mux_v
    port map (
            O => \N__23713\,
            I => \N__23708\
        );

    \I__5002\ : InMux
    port map (
            O => \N__23712\,
            I => \N__23705\
        );

    \I__5001\ : InMux
    port map (
            O => \N__23711\,
            I => \N__23702\
        );

    \I__5000\ : Span4Mux_v
    port map (
            O => \N__23708\,
            I => \N__23699\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__23705\,
            I => \N__23696\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__23702\,
            I => \N__23692\
        );

    \I__4997\ : Sp12to4
    port map (
            O => \N__23699\,
            I => \N__23689\
        );

    \I__4996\ : Span4Mux_v
    port map (
            O => \N__23696\,
            I => \N__23686\
        );

    \I__4995\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23683\
        );

    \I__4994\ : Sp12to4
    port map (
            O => \N__23692\,
            I => \N__23678\
        );

    \I__4993\ : Span12Mux_h
    port map (
            O => \N__23689\,
            I => \N__23678\
        );

    \I__4992\ : Odrv4
    port map (
            O => \N__23686\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__23683\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__4990\ : Odrv12
    port map (
            O => \N__23678\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__4989\ : CascadeMux
    port map (
            O => \N__23671\,
            I => \N__23668\
        );

    \I__4988\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23665\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__23665\,
            I => \N__23662\
        );

    \I__4986\ : Span4Mux_v
    port map (
            O => \N__23662\,
            I => \N__23659\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__23659\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_0\
        );

    \I__4984\ : CascadeMux
    port map (
            O => \N__23656\,
            I => \N__23653\
        );

    \I__4983\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23650\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__23650\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_5\
        );

    \I__4981\ : InMux
    port map (
            O => \N__23647\,
            I => \N__23644\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__23644\,
            I => \N__23641\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__23641\,
            I => \un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0\
        );

    \I__4978\ : CascadeMux
    port map (
            O => \N__23638\,
            I => \N__23635\
        );

    \I__4977\ : InMux
    port map (
            O => \N__23635\,
            I => \N__23632\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__23632\,
            I => \N__23629\
        );

    \I__4975\ : Odrv4
    port map (
            O => \N__23629\,
            I => \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_6\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__23626\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_2_cascade_\
        );

    \I__4973\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23620\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__23620\,
            I => \this_vga_signals.M_this_map_address_d_8_mZ0Z_2\
        );

    \I__4971\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23614\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__23614\,
            I => \N__23611\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__23611\,
            I => \N__23608\
        );

    \I__4968\ : Odrv4
    port map (
            O => \N__23608\,
            I => \this_vga_signals.M_this_map_address_q_mZ0Z_9\
        );

    \I__4967\ : CascadeMux
    port map (
            O => \N__23605\,
            I => \N__23602\
        );

    \I__4966\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23599\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__23599\,
            I => \this_vga_signals.M_this_map_address_d_5_mZ0Z_9\
        );

    \I__4964\ : CascadeMux
    port map (
            O => \N__23596\,
            I => \N__23592\
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__23595\,
            I => \N__23589\
        );

    \I__4962\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23586\
        );

    \I__4961\ : CascadeBuf
    port map (
            O => \N__23589\,
            I => \N__23583\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__23586\,
            I => \N__23580\
        );

    \I__4959\ : CascadeMux
    port map (
            O => \N__23583\,
            I => \N__23577\
        );

    \I__4958\ : Span4Mux_h
    port map (
            O => \N__23580\,
            I => \N__23574\
        );

    \I__4957\ : InMux
    port map (
            O => \N__23577\,
            I => \N__23571\
        );

    \I__4956\ : Span4Mux_h
    port map (
            O => \N__23574\,
            I => \N__23566\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__23571\,
            I => \N__23563\
        );

    \I__4954\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23560\
        );

    \I__4953\ : InMux
    port map (
            O => \N__23569\,
            I => \N__23557\
        );

    \I__4952\ : Sp12to4
    port map (
            O => \N__23566\,
            I => \N__23552\
        );

    \I__4951\ : Span12Mux_h
    port map (
            O => \N__23563\,
            I => \N__23552\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__23560\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__23557\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4948\ : Odrv12
    port map (
            O => \N__23552\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4947\ : CascadeMux
    port map (
            O => \N__23545\,
            I => \N__23542\
        );

    \I__4946\ : CascadeBuf
    port map (
            O => \N__23542\,
            I => \N__23539\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__23539\,
            I => \N__23536\
        );

    \I__4944\ : CascadeBuf
    port map (
            O => \N__23536\,
            I => \N__23533\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__23533\,
            I => \N__23530\
        );

    \I__4942\ : CascadeBuf
    port map (
            O => \N__23530\,
            I => \N__23527\
        );

    \I__4941\ : CascadeMux
    port map (
            O => \N__23527\,
            I => \N__23524\
        );

    \I__4940\ : CascadeBuf
    port map (
            O => \N__23524\,
            I => \N__23521\
        );

    \I__4939\ : CascadeMux
    port map (
            O => \N__23521\,
            I => \N__23518\
        );

    \I__4938\ : CascadeBuf
    port map (
            O => \N__23518\,
            I => \N__23515\
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__23515\,
            I => \N__23512\
        );

    \I__4936\ : CascadeBuf
    port map (
            O => \N__23512\,
            I => \N__23509\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__23509\,
            I => \N__23506\
        );

    \I__4934\ : CascadeBuf
    port map (
            O => \N__23506\,
            I => \N__23503\
        );

    \I__4933\ : CascadeMux
    port map (
            O => \N__23503\,
            I => \N__23500\
        );

    \I__4932\ : CascadeBuf
    port map (
            O => \N__23500\,
            I => \N__23497\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__23497\,
            I => \N__23494\
        );

    \I__4930\ : CascadeBuf
    port map (
            O => \N__23494\,
            I => \N__23491\
        );

    \I__4929\ : CascadeMux
    port map (
            O => \N__23491\,
            I => \N__23488\
        );

    \I__4928\ : CascadeBuf
    port map (
            O => \N__23488\,
            I => \N__23485\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__23485\,
            I => \N__23482\
        );

    \I__4926\ : CascadeBuf
    port map (
            O => \N__23482\,
            I => \N__23479\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__23479\,
            I => \N__23476\
        );

    \I__4924\ : CascadeBuf
    port map (
            O => \N__23476\,
            I => \N__23473\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__23473\,
            I => \N__23470\
        );

    \I__4922\ : CascadeBuf
    port map (
            O => \N__23470\,
            I => \N__23467\
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__23467\,
            I => \N__23464\
        );

    \I__4920\ : CascadeBuf
    port map (
            O => \N__23464\,
            I => \N__23461\
        );

    \I__4919\ : CascadeMux
    port map (
            O => \N__23461\,
            I => \N__23458\
        );

    \I__4918\ : CascadeBuf
    port map (
            O => \N__23458\,
            I => \N__23455\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__23455\,
            I => \N__23451\
        );

    \I__4916\ : CascadeMux
    port map (
            O => \N__23454\,
            I => \N__23448\
        );

    \I__4915\ : InMux
    port map (
            O => \N__23451\,
            I => \N__23445\
        );

    \I__4914\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23442\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__23445\,
            I => \N__23439\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__23442\,
            I => \N__23435\
        );

    \I__4911\ : Span4Mux_v
    port map (
            O => \N__23439\,
            I => \N__23432\
        );

    \I__4910\ : CascadeMux
    port map (
            O => \N__23438\,
            I => \N__23429\
        );

    \I__4909\ : Sp12to4
    port map (
            O => \N__23435\,
            I => \N__23423\
        );

    \I__4908\ : Span4Mux_h
    port map (
            O => \N__23432\,
            I => \N__23420\
        );

    \I__4907\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23417\
        );

    \I__4906\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23414\
        );

    \I__4905\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23409\
        );

    \I__4904\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23409\
        );

    \I__4903\ : Span12Mux_v
    port map (
            O => \N__23423\,
            I => \N__23406\
        );

    \I__4902\ : Span4Mux_h
    port map (
            O => \N__23420\,
            I => \N__23403\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__23417\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__23414\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__23409\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__4898\ : Odrv12
    port map (
            O => \N__23406\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__4897\ : Odrv4
    port map (
            O => \N__23403\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__4896\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23389\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__23389\,
            I => \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\
        );

    \I__4894\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23383\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__23383\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12\
        );

    \I__4892\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23377\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__23377\,
            I => \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\
        );

    \I__4890\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23371\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__23371\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13\
        );

    \I__4888\ : CascadeMux
    port map (
            O => \N__23368\,
            I => \N__23365\
        );

    \I__4887\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23362\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__23362\,
            I => \N__23359\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__23359\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_13\
        );

    \I__4884\ : InMux
    port map (
            O => \N__23356\,
            I => \N__23353\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__23353\,
            I => \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\
        );

    \I__4882\ : CascadeMux
    port map (
            O => \N__23350\,
            I => \N__23344\
        );

    \I__4881\ : CascadeMux
    port map (
            O => \N__23349\,
            I => \N__23341\
        );

    \I__4880\ : CascadeMux
    port map (
            O => \N__23348\,
            I => \N__23336\
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__23347\,
            I => \N__23333\
        );

    \I__4878\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23330\
        );

    \I__4877\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23327\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__23340\,
            I => \N__23324\
        );

    \I__4875\ : CascadeMux
    port map (
            O => \N__23339\,
            I => \N__23320\
        );

    \I__4874\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23316\
        );

    \I__4873\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23313\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23310\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__23327\,
            I => \N__23307\
        );

    \I__4870\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23300\
        );

    \I__4869\ : InMux
    port map (
            O => \N__23323\,
            I => \N__23300\
        );

    \I__4868\ : InMux
    port map (
            O => \N__23320\,
            I => \N__23300\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__23319\,
            I => \N__23297\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__23316\,
            I => \N__23294\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__23313\,
            I => \N__23290\
        );

    \I__4864\ : Span4Mux_v
    port map (
            O => \N__23310\,
            I => \N__23285\
        );

    \I__4863\ : Span4Mux_v
    port map (
            O => \N__23307\,
            I => \N__23285\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__23300\,
            I => \N__23282\
        );

    \I__4861\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23279\
        );

    \I__4860\ : Span4Mux_h
    port map (
            O => \N__23294\,
            I => \N__23276\
        );

    \I__4859\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23273\
        );

    \I__4858\ : Span12Mux_v
    port map (
            O => \N__23290\,
            I => \N__23268\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__23285\,
            I => \N__23263\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__23282\,
            I => \N__23263\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23260\
        );

    \I__4854\ : Span4Mux_h
    port map (
            O => \N__23276\,
            I => \N__23255\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__23273\,
            I => \N__23255\
        );

    \I__4852\ : InMux
    port map (
            O => \N__23272\,
            I => \N__23252\
        );

    \I__4851\ : InMux
    port map (
            O => \N__23271\,
            I => \N__23249\
        );

    \I__4850\ : Odrv12
    port map (
            O => \N__23268\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__23263\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__23260\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__23255\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__23252\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__23249\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__4844\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23233\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__23233\,
            I => \N__23230\
        );

    \I__4842\ : Odrv12
    port map (
            O => \N__23230\,
            I => \this_vga_signals.M_this_state_q_ns_0_o2_0_0_0\
        );

    \I__4841\ : CascadeMux
    port map (
            O => \N__23227\,
            I => \this_vga_signals.M_this_state_q_ns_0_o2_0_1Z0Z_0_cascade_\
        );

    \I__4840\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23221\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__23221\,
            I => \N__23218\
        );

    \I__4838\ : Odrv12
    port map (
            O => \N__23218\,
            I => \M_this_sprites_address_q_RNI1DGI7Z0Z_0\
        );

    \I__4837\ : InMux
    port map (
            O => \N__23215\,
            I => \N__23212\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__23212\,
            I => \N__23209\
        );

    \I__4835\ : Span12Mux_h
    port map (
            O => \N__23209\,
            I => \N__23206\
        );

    \I__4834\ : Odrv12
    port map (
            O => \N__23206\,
            I => \M_this_map_ram_read_data_5\
        );

    \I__4833\ : CascadeMux
    port map (
            O => \N__23203\,
            I => \N__23200\
        );

    \I__4832\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23193\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__23199\,
            I => \N__23189\
        );

    \I__4830\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23186\
        );

    \I__4829\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23180\
        );

    \I__4828\ : InMux
    port map (
            O => \N__23196\,
            I => \N__23180\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__23193\,
            I => \N__23177\
        );

    \I__4826\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23174\
        );

    \I__4825\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23171\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__23186\,
            I => \N__23168\
        );

    \I__4823\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23165\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__23180\,
            I => \N__23162\
        );

    \I__4821\ : Span4Mux_h
    port map (
            O => \N__23177\,
            I => \N__23154\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__23174\,
            I => \N__23154\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__23171\,
            I => \N__23154\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__23168\,
            I => \N__23149\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__23165\,
            I => \N__23149\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__23162\,
            I => \N__23146\
        );

    \I__4815\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23143\
        );

    \I__4814\ : Span4Mux_h
    port map (
            O => \N__23154\,
            I => \N__23140\
        );

    \I__4813\ : Span4Mux_h
    port map (
            O => \N__23149\,
            I => \N__23137\
        );

    \I__4812\ : Sp12to4
    port map (
            O => \N__23146\,
            I => \N__23132\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__23143\,
            I => \N__23132\
        );

    \I__4810\ : Span4Mux_v
    port map (
            O => \N__23140\,
            I => \N__23129\
        );

    \I__4809\ : Sp12to4
    port map (
            O => \N__23137\,
            I => \N__23124\
        );

    \I__4808\ : Span12Mux_h
    port map (
            O => \N__23132\,
            I => \N__23124\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__23129\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__4806\ : Odrv12
    port map (
            O => \N__23124\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__4805\ : InMux
    port map (
            O => \N__23119\,
            I => \un1_M_this_sprites_address_q_cry_5\
        );

    \I__4804\ : InMux
    port map (
            O => \N__23116\,
            I => \un1_M_this_sprites_address_q_cry_6\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__23113\,
            I => \N__23110\
        );

    \I__4802\ : CascadeBuf
    port map (
            O => \N__23110\,
            I => \N__23107\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__23107\,
            I => \N__23104\
        );

    \I__4800\ : CascadeBuf
    port map (
            O => \N__23104\,
            I => \N__23101\
        );

    \I__4799\ : CascadeMux
    port map (
            O => \N__23101\,
            I => \N__23098\
        );

    \I__4798\ : CascadeBuf
    port map (
            O => \N__23098\,
            I => \N__23095\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__23095\,
            I => \N__23092\
        );

    \I__4796\ : CascadeBuf
    port map (
            O => \N__23092\,
            I => \N__23089\
        );

    \I__4795\ : CascadeMux
    port map (
            O => \N__23089\,
            I => \N__23086\
        );

    \I__4794\ : CascadeBuf
    port map (
            O => \N__23086\,
            I => \N__23083\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__23083\,
            I => \N__23080\
        );

    \I__4792\ : CascadeBuf
    port map (
            O => \N__23080\,
            I => \N__23077\
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__23077\,
            I => \N__23074\
        );

    \I__4790\ : CascadeBuf
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__23071\,
            I => \N__23068\
        );

    \I__4788\ : CascadeBuf
    port map (
            O => \N__23068\,
            I => \N__23065\
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__23065\,
            I => \N__23062\
        );

    \I__4786\ : CascadeBuf
    port map (
            O => \N__23062\,
            I => \N__23059\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__23059\,
            I => \N__23056\
        );

    \I__4784\ : CascadeBuf
    port map (
            O => \N__23056\,
            I => \N__23053\
        );

    \I__4783\ : CascadeMux
    port map (
            O => \N__23053\,
            I => \N__23050\
        );

    \I__4782\ : CascadeBuf
    port map (
            O => \N__23050\,
            I => \N__23047\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__23047\,
            I => \N__23044\
        );

    \I__4780\ : CascadeBuf
    port map (
            O => \N__23044\,
            I => \N__23041\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__23041\,
            I => \N__23038\
        );

    \I__4778\ : CascadeBuf
    port map (
            O => \N__23038\,
            I => \N__23035\
        );

    \I__4777\ : CascadeMux
    port map (
            O => \N__23035\,
            I => \N__23032\
        );

    \I__4776\ : CascadeBuf
    port map (
            O => \N__23032\,
            I => \N__23029\
        );

    \I__4775\ : CascadeMux
    port map (
            O => \N__23029\,
            I => \N__23026\
        );

    \I__4774\ : CascadeBuf
    port map (
            O => \N__23026\,
            I => \N__23023\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__23023\,
            I => \N__23020\
        );

    \I__4772\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23017\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__23014\
        );

    \I__4770\ : Span4Mux_s1_v
    port map (
            O => \N__23014\,
            I => \N__23011\
        );

    \I__4769\ : Sp12to4
    port map (
            O => \N__23011\,
            I => \N__23006\
        );

    \I__4768\ : InMux
    port map (
            O => \N__23010\,
            I => \N__23003\
        );

    \I__4767\ : InMux
    port map (
            O => \N__23009\,
            I => \N__22999\
        );

    \I__4766\ : Span12Mux_h
    port map (
            O => \N__23006\,
            I => \N__22996\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__23003\,
            I => \N__22993\
        );

    \I__4764\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22990\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__22999\,
            I => \N__22985\
        );

    \I__4762\ : Span12Mux_v
    port map (
            O => \N__22996\,
            I => \N__22985\
        );

    \I__4761\ : Odrv4
    port map (
            O => \N__22993\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__22990\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__4759\ : Odrv12
    port map (
            O => \N__22985\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__4758\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22975\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__22975\,
            I => \N__22972\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__22972\,
            I => \un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0\
        );

    \I__4755\ : InMux
    port map (
            O => \N__22969\,
            I => \bfn_18_18_0_\
        );

    \I__4754\ : CascadeMux
    port map (
            O => \N__22966\,
            I => \N__22963\
        );

    \I__4753\ : CascadeBuf
    port map (
            O => \N__22963\,
            I => \N__22960\
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__22960\,
            I => \N__22957\
        );

    \I__4751\ : CascadeBuf
    port map (
            O => \N__22957\,
            I => \N__22954\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__22954\,
            I => \N__22951\
        );

    \I__4749\ : CascadeBuf
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__22948\,
            I => \N__22945\
        );

    \I__4747\ : CascadeBuf
    port map (
            O => \N__22945\,
            I => \N__22942\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__22942\,
            I => \N__22939\
        );

    \I__4745\ : CascadeBuf
    port map (
            O => \N__22939\,
            I => \N__22936\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__22936\,
            I => \N__22933\
        );

    \I__4743\ : CascadeBuf
    port map (
            O => \N__22933\,
            I => \N__22930\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__22930\,
            I => \N__22927\
        );

    \I__4741\ : CascadeBuf
    port map (
            O => \N__22927\,
            I => \N__22924\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__22924\,
            I => \N__22921\
        );

    \I__4739\ : CascadeBuf
    port map (
            O => \N__22921\,
            I => \N__22918\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__4737\ : CascadeBuf
    port map (
            O => \N__22915\,
            I => \N__22912\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__22912\,
            I => \N__22909\
        );

    \I__4735\ : CascadeBuf
    port map (
            O => \N__22909\,
            I => \N__22906\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__22906\,
            I => \N__22903\
        );

    \I__4733\ : CascadeBuf
    port map (
            O => \N__22903\,
            I => \N__22900\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__22900\,
            I => \N__22897\
        );

    \I__4731\ : CascadeBuf
    port map (
            O => \N__22897\,
            I => \N__22894\
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__22894\,
            I => \N__22891\
        );

    \I__4729\ : CascadeBuf
    port map (
            O => \N__22891\,
            I => \N__22888\
        );

    \I__4728\ : CascadeMux
    port map (
            O => \N__22888\,
            I => \N__22885\
        );

    \I__4727\ : CascadeBuf
    port map (
            O => \N__22885\,
            I => \N__22882\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__22882\,
            I => \N__22879\
        );

    \I__4725\ : CascadeBuf
    port map (
            O => \N__22879\,
            I => \N__22876\
        );

    \I__4724\ : CascadeMux
    port map (
            O => \N__22876\,
            I => \N__22873\
        );

    \I__4723\ : InMux
    port map (
            O => \N__22873\,
            I => \N__22870\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__22870\,
            I => \N__22867\
        );

    \I__4721\ : Span4Mux_h
    port map (
            O => \N__22867\,
            I => \N__22864\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__22864\,
            I => \N__22861\
        );

    \I__4719\ : Span4Mux_h
    port map (
            O => \N__22861\,
            I => \N__22856\
        );

    \I__4718\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22852\
        );

    \I__4717\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22849\
        );

    \I__4716\ : Sp12to4
    port map (
            O => \N__22856\,
            I => \N__22846\
        );

    \I__4715\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22843\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__22852\,
            I => \N__22836\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__22849\,
            I => \N__22836\
        );

    \I__4712\ : Span12Mux_s11_v
    port map (
            O => \N__22846\,
            I => \N__22836\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__22843\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4710\ : Odrv12
    port map (
            O => \N__22836\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4709\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22828\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__22828\,
            I => \N__22825\
        );

    \I__4707\ : Odrv12
    port map (
            O => \N__22825\,
            I => \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\
        );

    \I__4706\ : InMux
    port map (
            O => \N__22822\,
            I => \un1_M_this_sprites_address_q_cry_8\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__22819\,
            I => \N__22816\
        );

    \I__4704\ : CascadeBuf
    port map (
            O => \N__22816\,
            I => \N__22813\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__22813\,
            I => \N__22810\
        );

    \I__4702\ : CascadeBuf
    port map (
            O => \N__22810\,
            I => \N__22807\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__22807\,
            I => \N__22804\
        );

    \I__4700\ : CascadeBuf
    port map (
            O => \N__22804\,
            I => \N__22801\
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \N__22798\
        );

    \I__4698\ : CascadeBuf
    port map (
            O => \N__22798\,
            I => \N__22795\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__22795\,
            I => \N__22792\
        );

    \I__4696\ : CascadeBuf
    port map (
            O => \N__22792\,
            I => \N__22789\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__22789\,
            I => \N__22786\
        );

    \I__4694\ : CascadeBuf
    port map (
            O => \N__22786\,
            I => \N__22783\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__22783\,
            I => \N__22780\
        );

    \I__4692\ : CascadeBuf
    port map (
            O => \N__22780\,
            I => \N__22777\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__22777\,
            I => \N__22774\
        );

    \I__4690\ : CascadeBuf
    port map (
            O => \N__22774\,
            I => \N__22771\
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__22771\,
            I => \N__22768\
        );

    \I__4688\ : CascadeBuf
    port map (
            O => \N__22768\,
            I => \N__22765\
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__22765\,
            I => \N__22762\
        );

    \I__4686\ : CascadeBuf
    port map (
            O => \N__22762\,
            I => \N__22759\
        );

    \I__4685\ : CascadeMux
    port map (
            O => \N__22759\,
            I => \N__22756\
        );

    \I__4684\ : CascadeBuf
    port map (
            O => \N__22756\,
            I => \N__22753\
        );

    \I__4683\ : CascadeMux
    port map (
            O => \N__22753\,
            I => \N__22750\
        );

    \I__4682\ : CascadeBuf
    port map (
            O => \N__22750\,
            I => \N__22747\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__22747\,
            I => \N__22744\
        );

    \I__4680\ : CascadeBuf
    port map (
            O => \N__22744\,
            I => \N__22741\
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__22741\,
            I => \N__22738\
        );

    \I__4678\ : CascadeBuf
    port map (
            O => \N__22738\,
            I => \N__22735\
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__22735\,
            I => \N__22732\
        );

    \I__4676\ : CascadeBuf
    port map (
            O => \N__22732\,
            I => \N__22729\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__22729\,
            I => \N__22726\
        );

    \I__4674\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22723\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__22723\,
            I => \N__22720\
        );

    \I__4672\ : Span4Mux_s2_v
    port map (
            O => \N__22720\,
            I => \N__22716\
        );

    \I__4671\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22712\
        );

    \I__4670\ : Span4Mux_v
    port map (
            O => \N__22716\,
            I => \N__22709\
        );

    \I__4669\ : InMux
    port map (
            O => \N__22715\,
            I => \N__22705\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__22712\,
            I => \N__22702\
        );

    \I__4667\ : Sp12to4
    port map (
            O => \N__22709\,
            I => \N__22699\
        );

    \I__4666\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22696\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__22705\,
            I => \N__22691\
        );

    \I__4664\ : Span4Mux_h
    port map (
            O => \N__22702\,
            I => \N__22691\
        );

    \I__4663\ : Span12Mux_h
    port map (
            O => \N__22699\,
            I => \N__22688\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__22696\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__22691\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__4660\ : Odrv12
    port map (
            O => \N__22688\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__4659\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22678\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__22678\,
            I => \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0\
        );

    \I__4657\ : InMux
    port map (
            O => \N__22675\,
            I => \un1_M_this_sprites_address_q_cry_9\
        );

    \I__4656\ : InMux
    port map (
            O => \N__22672\,
            I => \un1_M_this_sprites_address_q_cry_10\
        );

    \I__4655\ : InMux
    port map (
            O => \N__22669\,
            I => \un1_M_this_sprites_address_q_cry_11\
        );

    \I__4654\ : InMux
    port map (
            O => \N__22666\,
            I => \un1_M_this_sprites_address_q_cry_12\
        );

    \I__4653\ : CascadeMux
    port map (
            O => \N__22663\,
            I => \N__22659\
        );

    \I__4652\ : InMux
    port map (
            O => \N__22662\,
            I => \N__22656\
        );

    \I__4651\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22650\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22647\
        );

    \I__4649\ : InMux
    port map (
            O => \N__22655\,
            I => \N__22640\
        );

    \I__4648\ : InMux
    port map (
            O => \N__22654\,
            I => \N__22640\
        );

    \I__4647\ : InMux
    port map (
            O => \N__22653\,
            I => \N__22640\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__22650\,
            I => \N__22637\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__22647\,
            I => \this_vga_signals.M_this_state_q_ns_15\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__22640\,
            I => \this_vga_signals.M_this_state_q_ns_15\
        );

    \I__4643\ : Odrv4
    port map (
            O => \N__22637\,
            I => \this_vga_signals.M_this_state_q_ns_15\
        );

    \I__4642\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22627\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N__22624\
        );

    \I__4640\ : Odrv4
    port map (
            O => \N__22624\,
            I => \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\
        );

    \I__4639\ : InMux
    port map (
            O => \N__22621\,
            I => \un1_M_this_sprites_address_q_cry_0\
        );

    \I__4638\ : CascadeMux
    port map (
            O => \N__22618\,
            I => \N__22615\
        );

    \I__4637\ : CascadeBuf
    port map (
            O => \N__22615\,
            I => \N__22612\
        );

    \I__4636\ : CascadeMux
    port map (
            O => \N__22612\,
            I => \N__22609\
        );

    \I__4635\ : CascadeBuf
    port map (
            O => \N__22609\,
            I => \N__22606\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__22606\,
            I => \N__22603\
        );

    \I__4633\ : CascadeBuf
    port map (
            O => \N__22603\,
            I => \N__22600\
        );

    \I__4632\ : CascadeMux
    port map (
            O => \N__22600\,
            I => \N__22597\
        );

    \I__4631\ : CascadeBuf
    port map (
            O => \N__22597\,
            I => \N__22594\
        );

    \I__4630\ : CascadeMux
    port map (
            O => \N__22594\,
            I => \N__22591\
        );

    \I__4629\ : CascadeBuf
    port map (
            O => \N__22591\,
            I => \N__22588\
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__22588\,
            I => \N__22585\
        );

    \I__4627\ : CascadeBuf
    port map (
            O => \N__22585\,
            I => \N__22582\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__22582\,
            I => \N__22579\
        );

    \I__4625\ : CascadeBuf
    port map (
            O => \N__22579\,
            I => \N__22576\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__22576\,
            I => \N__22573\
        );

    \I__4623\ : CascadeBuf
    port map (
            O => \N__22573\,
            I => \N__22570\
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__22570\,
            I => \N__22567\
        );

    \I__4621\ : CascadeBuf
    port map (
            O => \N__22567\,
            I => \N__22564\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__22564\,
            I => \N__22561\
        );

    \I__4619\ : CascadeBuf
    port map (
            O => \N__22561\,
            I => \N__22558\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__22558\,
            I => \N__22555\
        );

    \I__4617\ : CascadeBuf
    port map (
            O => \N__22555\,
            I => \N__22552\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__22552\,
            I => \N__22549\
        );

    \I__4615\ : CascadeBuf
    port map (
            O => \N__22549\,
            I => \N__22546\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__22546\,
            I => \N__22543\
        );

    \I__4613\ : CascadeBuf
    port map (
            O => \N__22543\,
            I => \N__22540\
        );

    \I__4612\ : CascadeMux
    port map (
            O => \N__22540\,
            I => \N__22537\
        );

    \I__4611\ : CascadeBuf
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__22534\,
            I => \N__22531\
        );

    \I__4609\ : CascadeBuf
    port map (
            O => \N__22531\,
            I => \N__22528\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__22528\,
            I => \N__22525\
        );

    \I__4607\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22522\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__22522\,
            I => \N__22519\
        );

    \I__4605\ : Span4Mux_v
    port map (
            O => \N__22519\,
            I => \N__22516\
        );

    \I__4604\ : Span4Mux_h
    port map (
            O => \N__22516\,
            I => \N__22512\
        );

    \I__4603\ : InMux
    port map (
            O => \N__22515\,
            I => \N__22509\
        );

    \I__4602\ : Sp12to4
    port map (
            O => \N__22512\,
            I => \N__22504\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__22509\,
            I => \N__22501\
        );

    \I__4600\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22496\
        );

    \I__4599\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22496\
        );

    \I__4598\ : Span12Mux_v
    port map (
            O => \N__22504\,
            I => \N__22493\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__22501\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__22496\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4595\ : Odrv12
    port map (
            O => \N__22493\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4594\ : InMux
    port map (
            O => \N__22486\,
            I => \N__22483\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__22483\,
            I => \N__22480\
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__22480\,
            I => \un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0\
        );

    \I__4591\ : InMux
    port map (
            O => \N__22477\,
            I => \un1_M_this_sprites_address_q_cry_1\
        );

    \I__4590\ : InMux
    port map (
            O => \N__22474\,
            I => \N__22471\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__22471\,
            I => \N__22468\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__22468\,
            I => \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\
        );

    \I__4587\ : InMux
    port map (
            O => \N__22465\,
            I => \un1_M_this_sprites_address_q_cry_2\
        );

    \I__4586\ : InMux
    port map (
            O => \N__22462\,
            I => \un1_M_this_sprites_address_q_cry_3\
        );

    \I__4585\ : InMux
    port map (
            O => \N__22459\,
            I => \un1_M_this_sprites_address_q_cry_4\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__22456\,
            I => \N__22453\
        );

    \I__4583\ : InMux
    port map (
            O => \N__22453\,
            I => \N__22450\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__22450\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_1\
        );

    \I__4581\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22444\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__22444\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__4578\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22435\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__22435\,
            I => \N__22432\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__22432\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_9\
        );

    \I__4575\ : CascadeMux
    port map (
            O => \N__22429\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2_cascade_\
        );

    \I__4574\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22423\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__22423\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_2\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__22420\,
            I => \N__22417\
        );

    \I__4571\ : InMux
    port map (
            O => \N__22417\,
            I => \N__22414\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__22414\,
            I => \N__22411\
        );

    \I__4569\ : Odrv4
    port map (
            O => \N__22411\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_3\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__22408\,
            I => \N__22405\
        );

    \I__4567\ : InMux
    port map (
            O => \N__22405\,
            I => \N__22402\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__22402\,
            I => \N__22399\
        );

    \I__4565\ : Span4Mux_v
    port map (
            O => \N__22399\,
            I => \N__22396\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__22396\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_10\
        );

    \I__4563\ : InMux
    port map (
            O => \N__22393\,
            I => \N__22390\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__22390\,
            I => \M_this_state_q_RNIMJ231Z0Z_8\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__22387\,
            I => \N__22384\
        );

    \I__4560\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22381\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__22381\,
            I => \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_3\
        );

    \I__4558\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22375\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__22375\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__22372\,
            I => \N__22369\
        );

    \I__4555\ : CascadeBuf
    port map (
            O => \N__22369\,
            I => \N__22366\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__22366\,
            I => \N__22363\
        );

    \I__4553\ : CascadeBuf
    port map (
            O => \N__22363\,
            I => \N__22360\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__22360\,
            I => \N__22357\
        );

    \I__4551\ : CascadeBuf
    port map (
            O => \N__22357\,
            I => \N__22354\
        );

    \I__4550\ : CascadeMux
    port map (
            O => \N__22354\,
            I => \N__22351\
        );

    \I__4549\ : CascadeBuf
    port map (
            O => \N__22351\,
            I => \N__22348\
        );

    \I__4548\ : CascadeMux
    port map (
            O => \N__22348\,
            I => \N__22345\
        );

    \I__4547\ : CascadeBuf
    port map (
            O => \N__22345\,
            I => \N__22342\
        );

    \I__4546\ : CascadeMux
    port map (
            O => \N__22342\,
            I => \N__22339\
        );

    \I__4545\ : CascadeBuf
    port map (
            O => \N__22339\,
            I => \N__22336\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__22336\,
            I => \N__22333\
        );

    \I__4543\ : CascadeBuf
    port map (
            O => \N__22333\,
            I => \N__22330\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__22330\,
            I => \N__22327\
        );

    \I__4541\ : CascadeBuf
    port map (
            O => \N__22327\,
            I => \N__22324\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__22324\,
            I => \N__22321\
        );

    \I__4539\ : CascadeBuf
    port map (
            O => \N__22321\,
            I => \N__22318\
        );

    \I__4538\ : CascadeMux
    port map (
            O => \N__22318\,
            I => \N__22315\
        );

    \I__4537\ : CascadeBuf
    port map (
            O => \N__22315\,
            I => \N__22312\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__22312\,
            I => \N__22309\
        );

    \I__4535\ : CascadeBuf
    port map (
            O => \N__22309\,
            I => \N__22306\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__22306\,
            I => \N__22303\
        );

    \I__4533\ : CascadeBuf
    port map (
            O => \N__22303\,
            I => \N__22300\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__22300\,
            I => \N__22297\
        );

    \I__4531\ : CascadeBuf
    port map (
            O => \N__22297\,
            I => \N__22294\
        );

    \I__4530\ : CascadeMux
    port map (
            O => \N__22294\,
            I => \N__22291\
        );

    \I__4529\ : CascadeBuf
    port map (
            O => \N__22291\,
            I => \N__22288\
        );

    \I__4528\ : CascadeMux
    port map (
            O => \N__22288\,
            I => \N__22285\
        );

    \I__4527\ : CascadeBuf
    port map (
            O => \N__22285\,
            I => \N__22281\
        );

    \I__4526\ : CascadeMux
    port map (
            O => \N__22284\,
            I => \N__22278\
        );

    \I__4525\ : CascadeMux
    port map (
            O => \N__22281\,
            I => \N__22275\
        );

    \I__4524\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22272\
        );

    \I__4523\ : InMux
    port map (
            O => \N__22275\,
            I => \N__22269\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__22272\,
            I => \N__22266\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__22269\,
            I => \N__22263\
        );

    \I__4520\ : Span4Mux_v
    port map (
            O => \N__22266\,
            I => \N__22259\
        );

    \I__4519\ : Span4Mux_v
    port map (
            O => \N__22263\,
            I => \N__22256\
        );

    \I__4518\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22253\
        );

    \I__4517\ : Sp12to4
    port map (
            O => \N__22259\,
            I => \N__22248\
        );

    \I__4516\ : Sp12to4
    port map (
            O => \N__22256\,
            I => \N__22245\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__22253\,
            I => \N__22242\
        );

    \I__4514\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22237\
        );

    \I__4513\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22237\
        );

    \I__4512\ : Span12Mux_h
    port map (
            O => \N__22248\,
            I => \N__22232\
        );

    \I__4511\ : Span12Mux_h
    port map (
            O => \N__22245\,
            I => \N__22232\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__22242\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__22237\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4508\ : Odrv12
    port map (
            O => \N__22232\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4507\ : CEMux
    port map (
            O => \N__22225\,
            I => \N__22221\
        );

    \I__4506\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22216\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__22221\,
            I => \N__22213\
        );

    \I__4504\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22210\
        );

    \I__4503\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22207\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__22216\,
            I => \N__22204\
        );

    \I__4501\ : Span4Mux_h
    port map (
            O => \N__22213\,
            I => \N__22201\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__22210\,
            I => \N__22196\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__22207\,
            I => \N__22196\
        );

    \I__4498\ : Span4Mux_h
    port map (
            O => \N__22204\,
            I => \N__22193\
        );

    \I__4497\ : Span4Mux_h
    port map (
            O => \N__22201\,
            I => \N__22190\
        );

    \I__4496\ : Span4Mux_v
    port map (
            O => \N__22196\,
            I => \N__22187\
        );

    \I__4495\ : Span4Mux_v
    port map (
            O => \N__22193\,
            I => \N__22184\
        );

    \I__4494\ : Odrv4
    port map (
            O => \N__22190\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__22187\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__22184\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__22177\,
            I => \N__22174\
        );

    \I__4490\ : CascadeBuf
    port map (
            O => \N__22174\,
            I => \N__22171\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__22171\,
            I => \N__22168\
        );

    \I__4488\ : CascadeBuf
    port map (
            O => \N__22168\,
            I => \N__22165\
        );

    \I__4487\ : CascadeMux
    port map (
            O => \N__22165\,
            I => \N__22162\
        );

    \I__4486\ : CascadeBuf
    port map (
            O => \N__22162\,
            I => \N__22159\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__22159\,
            I => \N__22156\
        );

    \I__4484\ : CascadeBuf
    port map (
            O => \N__22156\,
            I => \N__22153\
        );

    \I__4483\ : CascadeMux
    port map (
            O => \N__22153\,
            I => \N__22150\
        );

    \I__4482\ : CascadeBuf
    port map (
            O => \N__22150\,
            I => \N__22147\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__22147\,
            I => \N__22144\
        );

    \I__4480\ : CascadeBuf
    port map (
            O => \N__22144\,
            I => \N__22141\
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__22141\,
            I => \N__22138\
        );

    \I__4478\ : CascadeBuf
    port map (
            O => \N__22138\,
            I => \N__22135\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__4476\ : CascadeBuf
    port map (
            O => \N__22132\,
            I => \N__22129\
        );

    \I__4475\ : CascadeMux
    port map (
            O => \N__22129\,
            I => \N__22126\
        );

    \I__4474\ : CascadeBuf
    port map (
            O => \N__22126\,
            I => \N__22123\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__22123\,
            I => \N__22120\
        );

    \I__4472\ : CascadeBuf
    port map (
            O => \N__22120\,
            I => \N__22117\
        );

    \I__4471\ : CascadeMux
    port map (
            O => \N__22117\,
            I => \N__22114\
        );

    \I__4470\ : CascadeBuf
    port map (
            O => \N__22114\,
            I => \N__22111\
        );

    \I__4469\ : CascadeMux
    port map (
            O => \N__22111\,
            I => \N__22108\
        );

    \I__4468\ : CascadeBuf
    port map (
            O => \N__22108\,
            I => \N__22105\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__22105\,
            I => \N__22102\
        );

    \I__4466\ : CascadeBuf
    port map (
            O => \N__22102\,
            I => \N__22099\
        );

    \I__4465\ : CascadeMux
    port map (
            O => \N__22099\,
            I => \N__22096\
        );

    \I__4464\ : CascadeBuf
    port map (
            O => \N__22096\,
            I => \N__22093\
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__22093\,
            I => \N__22090\
        );

    \I__4462\ : CascadeBuf
    port map (
            O => \N__22090\,
            I => \N__22087\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__22087\,
            I => \N__22083\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__22086\,
            I => \N__22080\
        );

    \I__4459\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22077\
        );

    \I__4458\ : InMux
    port map (
            O => \N__22080\,
            I => \N__22073\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__22077\,
            I => \N__22070\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__22076\,
            I => \N__22067\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22063\
        );

    \I__4454\ : Span4Mux_s3_v
    port map (
            O => \N__22070\,
            I => \N__22060\
        );

    \I__4453\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22057\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__22066\,
            I => \N__22054\
        );

    \I__4451\ : Sp12to4
    port map (
            O => \N__22063\,
            I => \N__22051\
        );

    \I__4450\ : Sp12to4
    port map (
            O => \N__22060\,
            I => \N__22048\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__22057\,
            I => \N__22045\
        );

    \I__4448\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22042\
        );

    \I__4447\ : Span12Mux_v
    port map (
            O => \N__22051\,
            I => \N__22039\
        );

    \I__4446\ : Span12Mux_h
    port map (
            O => \N__22048\,
            I => \N__22036\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__22045\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__22042\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4443\ : Odrv12
    port map (
            O => \N__22039\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4442\ : Odrv12
    port map (
            O => \N__22036\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4441\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22017\
        );

    \I__4440\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22017\
        );

    \I__4439\ : InMux
    port map (
            O => \N__22025\,
            I => \N__22012\
        );

    \I__4438\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22012\
        );

    \I__4437\ : InMux
    port map (
            O => \N__22023\,
            I => \N__22005\
        );

    \I__4436\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22002\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__22017\,
            I => \N__21998\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__22012\,
            I => \N__21995\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__22011\,
            I => \N__21991\
        );

    \I__4432\ : InMux
    port map (
            O => \N__22010\,
            I => \N__21984\
        );

    \I__4431\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21979\
        );

    \I__4430\ : InMux
    port map (
            O => \N__22008\,
            I => \N__21979\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__22005\,
            I => \N__21976\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__22002\,
            I => \N__21973\
        );

    \I__4427\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21969\
        );

    \I__4426\ : Span4Mux_v
    port map (
            O => \N__21998\,
            I => \N__21964\
        );

    \I__4425\ : Span4Mux_v
    port map (
            O => \N__21995\,
            I => \N__21964\
        );

    \I__4424\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21961\
        );

    \I__4423\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21958\
        );

    \I__4422\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21955\
        );

    \I__4421\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21948\
        );

    \I__4420\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21948\
        );

    \I__4419\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21948\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__21984\,
            I => \N__21945\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__21979\,
            I => \N__21940\
        );

    \I__4416\ : Span4Mux_v
    port map (
            O => \N__21976\,
            I => \N__21940\
        );

    \I__4415\ : Span4Mux_v
    port map (
            O => \N__21973\,
            I => \N__21937\
        );

    \I__4414\ : InMux
    port map (
            O => \N__21972\,
            I => \N__21934\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__21969\,
            I => \N__21929\
        );

    \I__4412\ : Span4Mux_h
    port map (
            O => \N__21964\,
            I => \N__21929\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__21961\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__21958\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__21955\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__21948\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__21945\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__4406\ : Odrv4
    port map (
            O => \N__21940\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__21937\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__21934\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__21929\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__4402\ : InMux
    port map (
            O => \N__21910\,
            I => \N__21907\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__21907\,
            I => \N__21904\
        );

    \I__4400\ : Odrv4
    port map (
            O => \N__21904\,
            I => \M_this_state_q_RNI2S2SZ0Z_13\
        );

    \I__4399\ : CascadeMux
    port map (
            O => \N__21901\,
            I => \M_this_state_q_RNITS9I4Z0Z_7_cascade_\
        );

    \I__4398\ : IoInMux
    port map (
            O => \N__21898\,
            I => \N__21895\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__21895\,
            I => \N__21892\
        );

    \I__4396\ : IoSpan4Mux
    port map (
            O => \N__21892\,
            I => \N__21889\
        );

    \I__4395\ : Span4Mux_s3_h
    port map (
            O => \N__21889\,
            I => \N__21886\
        );

    \I__4394\ : Sp12to4
    port map (
            O => \N__21886\,
            I => \N__21883\
        );

    \I__4393\ : Span12Mux_s11_h
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__4392\ : Span12Mux_v
    port map (
            O => \N__21880\,
            I => \N__21877\
        );

    \I__4391\ : Odrv12
    port map (
            O => \N__21877\,
            I => dma_ac0_5_i
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__21874\,
            I => \dma_ac0_5_i_cascade_\
        );

    \I__4389\ : IoInMux
    port map (
            O => \N__21871\,
            I => \N__21868\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__21868\,
            I => \N__21862\
        );

    \I__4387\ : IoInMux
    port map (
            O => \N__21867\,
            I => \N__21859\
        );

    \I__4386\ : IoInMux
    port map (
            O => \N__21866\,
            I => \N__21855\
        );

    \I__4385\ : IoInMux
    port map (
            O => \N__21865\,
            I => \N__21849\
        );

    \I__4384\ : IoSpan4Mux
    port map (
            O => \N__21862\,
            I => \N__21843\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__21859\,
            I => \N__21843\
        );

    \I__4382\ : IoInMux
    port map (
            O => \N__21858\,
            I => \N__21840\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__21855\,
            I => \N__21836\
        );

    \I__4380\ : IoInMux
    port map (
            O => \N__21854\,
            I => \N__21833\
        );

    \I__4379\ : IoInMux
    port map (
            O => \N__21853\,
            I => \N__21830\
        );

    \I__4378\ : IoInMux
    port map (
            O => \N__21852\,
            I => \N__21827\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__21849\,
            I => \N__21823\
        );

    \I__4376\ : IoInMux
    port map (
            O => \N__21848\,
            I => \N__21819\
        );

    \I__4375\ : IoSpan4Mux
    port map (
            O => \N__21843\,
            I => \N__21814\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__21840\,
            I => \N__21814\
        );

    \I__4373\ : IoInMux
    port map (
            O => \N__21839\,
            I => \N__21811\
        );

    \I__4372\ : IoSpan4Mux
    port map (
            O => \N__21836\,
            I => \N__21802\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__21833\,
            I => \N__21802\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__21830\,
            I => \N__21802\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__21827\,
            I => \N__21799\
        );

    \I__4368\ : IoInMux
    port map (
            O => \N__21826\,
            I => \N__21796\
        );

    \I__4367\ : IoSpan4Mux
    port map (
            O => \N__21823\,
            I => \N__21793\
        );

    \I__4366\ : IoInMux
    port map (
            O => \N__21822\,
            I => \N__21790\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__21819\,
            I => \N__21787\
        );

    \I__4364\ : IoSpan4Mux
    port map (
            O => \N__21814\,
            I => \N__21782\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__21811\,
            I => \N__21782\
        );

    \I__4362\ : IoInMux
    port map (
            O => \N__21810\,
            I => \N__21779\
        );

    \I__4361\ : IoInMux
    port map (
            O => \N__21809\,
            I => \N__21776\
        );

    \I__4360\ : IoSpan4Mux
    port map (
            O => \N__21802\,
            I => \N__21768\
        );

    \I__4359\ : IoSpan4Mux
    port map (
            O => \N__21799\,
            I => \N__21768\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__21796\,
            I => \N__21768\
        );

    \I__4357\ : IoSpan4Mux
    port map (
            O => \N__21793\,
            I => \N__21763\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__21790\,
            I => \N__21763\
        );

    \I__4355\ : IoSpan4Mux
    port map (
            O => \N__21787\,
            I => \N__21760\
        );

    \I__4354\ : IoSpan4Mux
    port map (
            O => \N__21782\,
            I => \N__21755\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__21779\,
            I => \N__21755\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__21776\,
            I => \N__21752\
        );

    \I__4351\ : IoInMux
    port map (
            O => \N__21775\,
            I => \N__21749\
        );

    \I__4350\ : IoSpan4Mux
    port map (
            O => \N__21768\,
            I => \N__21744\
        );

    \I__4349\ : IoSpan4Mux
    port map (
            O => \N__21763\,
            I => \N__21744\
        );

    \I__4348\ : Span4Mux_s3_h
    port map (
            O => \N__21760\,
            I => \N__21740\
        );

    \I__4347\ : IoSpan4Mux
    port map (
            O => \N__21755\,
            I => \N__21735\
        );

    \I__4346\ : IoSpan4Mux
    port map (
            O => \N__21752\,
            I => \N__21735\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__21749\,
            I => \N__21731\
        );

    \I__4344\ : Span4Mux_s0_h
    port map (
            O => \N__21744\,
            I => \N__21728\
        );

    \I__4343\ : IoInMux
    port map (
            O => \N__21743\,
            I => \N__21725\
        );

    \I__4342\ : Span4Mux_v
    port map (
            O => \N__21740\,
            I => \N__21722\
        );

    \I__4341\ : Span4Mux_s3_v
    port map (
            O => \N__21735\,
            I => \N__21719\
        );

    \I__4340\ : IoInMux
    port map (
            O => \N__21734\,
            I => \N__21716\
        );

    \I__4339\ : Span12Mux_s9_h
    port map (
            O => \N__21731\,
            I => \N__21713\
        );

    \I__4338\ : Sp12to4
    port map (
            O => \N__21728\,
            I => \N__21708\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21708\
        );

    \I__4336\ : Sp12to4
    port map (
            O => \N__21722\,
            I => \N__21705\
        );

    \I__4335\ : Sp12to4
    port map (
            O => \N__21719\,
            I => \N__21700\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21700\
        );

    \I__4333\ : Span12Mux_v
    port map (
            O => \N__21713\,
            I => \N__21695\
        );

    \I__4332\ : Span12Mux_s9_h
    port map (
            O => \N__21708\,
            I => \N__21695\
        );

    \I__4331\ : Span12Mux_h
    port map (
            O => \N__21705\,
            I => \N__21690\
        );

    \I__4330\ : Span12Mux_s5_v
    port map (
            O => \N__21700\,
            I => \N__21690\
        );

    \I__4329\ : Odrv12
    port map (
            O => \N__21695\,
            I => dma_ac0_5_i_i
        );

    \I__4328\ : Odrv12
    port map (
            O => \N__21690\,
            I => dma_ac0_5_i_i
        );

    \I__4327\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21682\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__21682\,
            I => \this_vga_signals.un23_i_a2_4Z0Z_0\
        );

    \I__4325\ : InMux
    port map (
            O => \N__21679\,
            I => \N__21676\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__21676\,
            I => \M_this_state_q_RNI6Q0SZ0Z_7\
        );

    \I__4323\ : InMux
    port map (
            O => \N__21673\,
            I => \N__21670\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__21670\,
            I => \N__21667\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__21667\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__21664\,
            I => \N__21661\
        );

    \I__4319\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21658\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__21658\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_8\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__21655\,
            I => \this_vga_signals.un23_i_a2_x1Z0Z_0_cascade_\
        );

    \I__4316\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21649\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__21649\,
            I => \N__21646\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__21643\,
            I => \N__21638\
        );

    \I__4312\ : InMux
    port map (
            O => \N__21642\,
            I => \N__21635\
        );

    \I__4311\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21632\
        );

    \I__4310\ : Sp12to4
    port map (
            O => \N__21638\,
            I => \N__21627\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__21635\,
            I => \N__21627\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__21632\,
            I => \N__21624\
        );

    \I__4307\ : Span12Mux_s4_h
    port map (
            O => \N__21627\,
            I => \N__21621\
        );

    \I__4306\ : Span4Mux_v
    port map (
            O => \N__21624\,
            I => \N__21618\
        );

    \I__4305\ : Span12Mux_h
    port map (
            O => \N__21621\,
            I => \N__21615\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__21618\,
            I => \N__21612\
        );

    \I__4303\ : Odrv12
    port map (
            O => \N__21615\,
            I => \dma_ac0Z0Z_5\
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__21612\,
            I => \dma_ac0Z0Z_5\
        );

    \I__4301\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21604\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__21604\,
            I => this_vga_signals_un23_i_a2_1_3
        );

    \I__4299\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21598\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__21598\,
            I => this_vga_signals_un23_i_a2_4_2
        );

    \I__4297\ : CascadeMux
    port map (
            O => \N__21595\,
            I => \this_vga_signals_un23_i_a2_3_2_cascade_\
        );

    \I__4296\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__21589\,
            I => dma_c3_0
        );

    \I__4294\ : InMux
    port map (
            O => \N__21586\,
            I => \N__21582\
        );

    \I__4293\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21579\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__21582\,
            I => dma_axb0
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__21579\,
            I => dma_axb0
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__21574\,
            I => \N__21571\
        );

    \I__4289\ : CascadeBuf
    port map (
            O => \N__21571\,
            I => \N__21568\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__21568\,
            I => \N__21565\
        );

    \I__4287\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21562\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__21562\,
            I => \N__21559\
        );

    \I__4285\ : Span4Mux_s2_v
    port map (
            O => \N__21559\,
            I => \N__21556\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__21556\,
            I => \N__21552\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__21555\,
            I => \N__21548\
        );

    \I__4282\ : Span4Mux_h
    port map (
            O => \N__21552\,
            I => \N__21544\
        );

    \I__4281\ : InMux
    port map (
            O => \N__21551\,
            I => \N__21541\
        );

    \I__4280\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21538\
        );

    \I__4279\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21535\
        );

    \I__4278\ : Span4Mux_v
    port map (
            O => \N__21544\,
            I => \N__21532\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__21541\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__21538\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__21535\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__4274\ : Odrv4
    port map (
            O => \N__21532\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__4273\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21518\
        );

    \I__4272\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21515\
        );

    \I__4271\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21512\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__21518\,
            I => \this_ppu.un1_M_vaddress_q_c5\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__21515\,
            I => \this_ppu.un1_M_vaddress_q_c5\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__21512\,
            I => \this_ppu.un1_M_vaddress_q_c5\
        );

    \I__4267\ : SRMux
    port map (
            O => \N__21505\,
            I => \N__21500\
        );

    \I__4266\ : SRMux
    port map (
            O => \N__21504\,
            I => \N__21497\
        );

    \I__4265\ : SRMux
    port map (
            O => \N__21503\,
            I => \N__21494\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__21500\,
            I => \N__21489\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__21497\,
            I => \N__21484\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__21494\,
            I => \N__21484\
        );

    \I__4261\ : SRMux
    port map (
            O => \N__21493\,
            I => \N__21481\
        );

    \I__4260\ : SRMux
    port map (
            O => \N__21492\,
            I => \N__21478\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__21489\,
            I => \N__21471\
        );

    \I__4258\ : Span4Mux_v
    port map (
            O => \N__21484\,
            I => \N__21471\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__21481\,
            I => \N__21471\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__21478\,
            I => \N__21468\
        );

    \I__4255\ : Span4Mux_h
    port map (
            O => \N__21471\,
            I => \N__21463\
        );

    \I__4254\ : Span4Mux_v
    port map (
            O => \N__21468\,
            I => \N__21460\
        );

    \I__4253\ : SRMux
    port map (
            O => \N__21467\,
            I => \N__21457\
        );

    \I__4252\ : SRMux
    port map (
            O => \N__21466\,
            I => \N__21454\
        );

    \I__4251\ : Odrv4
    port map (
            O => \N__21463\,
            I => \this_ppu.M_last_q_RNIQKTIG\
        );

    \I__4250\ : Odrv4
    port map (
            O => \N__21460\,
            I => \this_ppu.M_last_q_RNIQKTIG\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__21457\,
            I => \this_ppu.M_last_q_RNIQKTIG\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__21454\,
            I => \this_ppu.M_last_q_RNIQKTIG\
        );

    \I__4247\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21441\
        );

    \I__4246\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21438\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__21441\,
            I => \this_ppu.M_vaddress_qZ0Z_7\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__21438\,
            I => \this_ppu.M_vaddress_qZ0Z_7\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__21433\,
            I => \N__21430\
        );

    \I__4242\ : CascadeBuf
    port map (
            O => \N__21430\,
            I => \N__21427\
        );

    \I__4241\ : CascadeMux
    port map (
            O => \N__21427\,
            I => \N__21424\
        );

    \I__4240\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21421\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21418\
        );

    \I__4238\ : Span12Mux_h
    port map (
            O => \N__21418\,
            I => \N__21415\
        );

    \I__4237\ : Odrv12
    port map (
            O => \N__21415\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__4236\ : IoInMux
    port map (
            O => \N__21412\,
            I => \N__21409\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__21409\,
            I => \N__21406\
        );

    \I__4234\ : IoSpan4Mux
    port map (
            O => \N__21406\,
            I => \N__21403\
        );

    \I__4233\ : Span4Mux_s0_v
    port map (
            O => \N__21403\,
            I => \N__21400\
        );

    \I__4232\ : Span4Mux_v
    port map (
            O => \N__21400\,
            I => \N__21397\
        );

    \I__4231\ : Span4Mux_v
    port map (
            O => \N__21397\,
            I => \N__21394\
        );

    \I__4230\ : Sp12to4
    port map (
            O => \N__21394\,
            I => \N__21391\
        );

    \I__4229\ : Odrv12
    port map (
            O => \N__21391\,
            I => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\
        );

    \I__4228\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21384\
        );

    \I__4227\ : InMux
    port map (
            O => \N__21387\,
            I => \N__21380\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__21384\,
            I => \N__21376\
        );

    \I__4225\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21373\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21369\
        );

    \I__4223\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21366\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__21376\,
            I => \N__21362\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__21373\,
            I => \N__21359\
        );

    \I__4220\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21356\
        );

    \I__4219\ : Span4Mux_v
    port map (
            O => \N__21369\,
            I => \N__21350\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__21366\,
            I => \N__21350\
        );

    \I__4217\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21347\
        );

    \I__4216\ : Span4Mux_v
    port map (
            O => \N__21362\,
            I => \N__21341\
        );

    \I__4215\ : Span4Mux_h
    port map (
            O => \N__21359\,
            I => \N__21341\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__21356\,
            I => \N__21338\
        );

    \I__4213\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21335\
        );

    \I__4212\ : Span4Mux_v
    port map (
            O => \N__21350\,
            I => \N__21330\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__21347\,
            I => \N__21330\
        );

    \I__4210\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21327\
        );

    \I__4209\ : Span4Mux_v
    port map (
            O => \N__21341\,
            I => \N__21322\
        );

    \I__4208\ : Span4Mux_h
    port map (
            O => \N__21338\,
            I => \N__21322\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21319\
        );

    \I__4206\ : Span4Mux_v
    port map (
            O => \N__21330\,
            I => \N__21314\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__21327\,
            I => \N__21314\
        );

    \I__4204\ : Span4Mux_v
    port map (
            O => \N__21322\,
            I => \N__21309\
        );

    \I__4203\ : Span4Mux_h
    port map (
            O => \N__21319\,
            I => \N__21309\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__21314\,
            I => \N__21306\
        );

    \I__4201\ : Span4Mux_h
    port map (
            O => \N__21309\,
            I => \N__21301\
        );

    \I__4200\ : Span4Mux_h
    port map (
            O => \N__21306\,
            I => \N__21301\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__21301\,
            I => \M_this_sprites_ram_write_data_0\
        );

    \I__4198\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21294\
        );

    \I__4197\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21290\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__21294\,
            I => \N__21286\
        );

    \I__4195\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21283\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__21290\,
            I => \N__21279\
        );

    \I__4193\ : InMux
    port map (
            O => \N__21289\,
            I => \N__21276\
        );

    \I__4192\ : Span4Mux_v
    port map (
            O => \N__21286\,
            I => \N__21270\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__21283\,
            I => \N__21270\
        );

    \I__4190\ : InMux
    port map (
            O => \N__21282\,
            I => \N__21267\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__21279\,
            I => \N__21264\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__21276\,
            I => \N__21261\
        );

    \I__4187\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21258\
        );

    \I__4186\ : Span4Mux_v
    port map (
            O => \N__21270\,
            I => \N__21253\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__21267\,
            I => \N__21253\
        );

    \I__4184\ : Span4Mux_v
    port map (
            O => \N__21264\,
            I => \N__21247\
        );

    \I__4183\ : Span4Mux_h
    port map (
            O => \N__21261\,
            I => \N__21247\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__21258\,
            I => \N__21244\
        );

    \I__4181\ : Span4Mux_v
    port map (
            O => \N__21253\,
            I => \N__21241\
        );

    \I__4180\ : InMux
    port map (
            O => \N__21252\,
            I => \N__21238\
        );

    \I__4179\ : Span4Mux_v
    port map (
            O => \N__21247\,
            I => \N__21232\
        );

    \I__4178\ : Span4Mux_h
    port map (
            O => \N__21244\,
            I => \N__21232\
        );

    \I__4177\ : Span4Mux_v
    port map (
            O => \N__21241\,
            I => \N__21227\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__21238\,
            I => \N__21227\
        );

    \I__4175\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21224\
        );

    \I__4174\ : Span4Mux_v
    port map (
            O => \N__21232\,
            I => \N__21219\
        );

    \I__4173\ : Span4Mux_h
    port map (
            O => \N__21227\,
            I => \N__21219\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21216\
        );

    \I__4171\ : Span4Mux_h
    port map (
            O => \N__21219\,
            I => \N__21213\
        );

    \I__4170\ : Span12Mux_s10_h
    port map (
            O => \N__21216\,
            I => \N__21210\
        );

    \I__4169\ : Odrv4
    port map (
            O => \N__21213\,
            I => \M_this_sprites_ram_write_data_1\
        );

    \I__4168\ : Odrv12
    port map (
            O => \N__21210\,
            I => \M_this_sprites_ram_write_data_1\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__21205\,
            I => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux_cascade_\
        );

    \I__4166\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21199\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21192\
        );

    \I__4164\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21189\
        );

    \I__4163\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21186\
        );

    \I__4162\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21183\
        );

    \I__4161\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21178\
        );

    \I__4160\ : Span4Mux_v
    port map (
            O => \N__21192\,
            I => \N__21174\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__21189\,
            I => \N__21171\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21168\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__21183\,
            I => \N__21165\
        );

    \I__4156\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21162\
        );

    \I__4155\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21159\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__21178\,
            I => \N__21156\
        );

    \I__4153\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21153\
        );

    \I__4152\ : Sp12to4
    port map (
            O => \N__21174\,
            I => \N__21146\
        );

    \I__4151\ : Sp12to4
    port map (
            O => \N__21171\,
            I => \N__21146\
        );

    \I__4150\ : Sp12to4
    port map (
            O => \N__21168\,
            I => \N__21146\
        );

    \I__4149\ : Sp12to4
    port map (
            O => \N__21165\,
            I => \N__21143\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__21162\,
            I => \N__21140\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__21159\,
            I => \N__21137\
        );

    \I__4146\ : Span12Mux_h
    port map (
            O => \N__21156\,
            I => \N__21134\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__21153\,
            I => \N__21131\
        );

    \I__4144\ : Span12Mux_v
    port map (
            O => \N__21146\,
            I => \N__21126\
        );

    \I__4143\ : Span12Mux_v
    port map (
            O => \N__21143\,
            I => \N__21126\
        );

    \I__4142\ : Span12Mux_h
    port map (
            O => \N__21140\,
            I => \N__21121\
        );

    \I__4141\ : Span12Mux_h
    port map (
            O => \N__21137\,
            I => \N__21121\
        );

    \I__4140\ : Span12Mux_v
    port map (
            O => \N__21134\,
            I => \N__21116\
        );

    \I__4139\ : Span12Mux_h
    port map (
            O => \N__21131\,
            I => \N__21116\
        );

    \I__4138\ : Odrv12
    port map (
            O => \N__21126\,
            I => \M_this_sprites_ram_write_data_2\
        );

    \I__4137\ : Odrv12
    port map (
            O => \N__21121\,
            I => \M_this_sprites_ram_write_data_2\
        );

    \I__4136\ : Odrv12
    port map (
            O => \N__21116\,
            I => \M_this_sprites_ram_write_data_2\
        );

    \I__4135\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21106\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__21106\,
            I => \N__21101\
        );

    \I__4133\ : InMux
    port map (
            O => \N__21105\,
            I => \N__21096\
        );

    \I__4132\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21096\
        );

    \I__4131\ : Odrv4
    port map (
            O => \N__21101\,
            I => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__21096\,
            I => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\
        );

    \I__4129\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21086\
        );

    \I__4128\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21082\
        );

    \I__4127\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21078\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__21086\,
            I => \N__21074\
        );

    \I__4125\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21071\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__21082\,
            I => \N__21067\
        );

    \I__4123\ : InMux
    port map (
            O => \N__21081\,
            I => \N__21064\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__21078\,
            I => \N__21061\
        );

    \I__4121\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21058\
        );

    \I__4120\ : Span4Mux_v
    port map (
            O => \N__21074\,
            I => \N__21053\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__21071\,
            I => \N__21053\
        );

    \I__4118\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21050\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__21067\,
            I => \N__21046\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__21064\,
            I => \N__21043\
        );

    \I__4115\ : Span4Mux_v
    port map (
            O => \N__21061\,
            I => \N__21038\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21038\
        );

    \I__4113\ : Span4Mux_v
    port map (
            O => \N__21053\,
            I => \N__21033\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__21050\,
            I => \N__21033\
        );

    \I__4111\ : InMux
    port map (
            O => \N__21049\,
            I => \N__21030\
        );

    \I__4110\ : Span4Mux_v
    port map (
            O => \N__21046\,
            I => \N__21025\
        );

    \I__4109\ : Span4Mux_h
    port map (
            O => \N__21043\,
            I => \N__21025\
        );

    \I__4108\ : Sp12to4
    port map (
            O => \N__21038\,
            I => \N__21022\
        );

    \I__4107\ : Span4Mux_v
    port map (
            O => \N__21033\,
            I => \N__21019\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__21030\,
            I => \N__21016\
        );

    \I__4105\ : Span4Mux_h
    port map (
            O => \N__21025\,
            I => \N__21013\
        );

    \I__4104\ : Span12Mux_v
    port map (
            O => \N__21022\,
            I => \N__21006\
        );

    \I__4103\ : Sp12to4
    port map (
            O => \N__21019\,
            I => \N__21006\
        );

    \I__4102\ : Span12Mux_s8_h
    port map (
            O => \N__21016\,
            I => \N__21006\
        );

    \I__4101\ : Odrv4
    port map (
            O => \N__21013\,
            I => \M_this_sprites_ram_write_data_3\
        );

    \I__4100\ : Odrv12
    port map (
            O => \N__21006\,
            I => \M_this_sprites_ram_write_data_3\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__21001\,
            I => \N__20995\
        );

    \I__4098\ : InMux
    port map (
            O => \N__21000\,
            I => \N__20992\
        );

    \I__4097\ : InMux
    port map (
            O => \N__20999\,
            I => \N__20988\
        );

    \I__4096\ : InMux
    port map (
            O => \N__20998\,
            I => \N__20983\
        );

    \I__4095\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20983\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__20992\,
            I => \N__20978\
        );

    \I__4093\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20975\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__20988\,
            I => \N__20972\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__20983\,
            I => \N__20969\
        );

    \I__4090\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20964\
        );

    \I__4089\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20964\
        );

    \I__4088\ : Span4Mux_v
    port map (
            O => \N__20978\,
            I => \N__20959\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20956\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__20972\,
            I => \N__20949\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__20969\,
            I => \N__20949\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__20964\,
            I => \N__20949\
        );

    \I__4083\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20946\
        );

    \I__4082\ : InMux
    port map (
            O => \N__20962\,
            I => \N__20943\
        );

    \I__4081\ : Sp12to4
    port map (
            O => \N__20959\,
            I => \N__20938\
        );

    \I__4080\ : Sp12to4
    port map (
            O => \N__20956\,
            I => \N__20938\
        );

    \I__4079\ : Span4Mux_h
    port map (
            O => \N__20949\,
            I => \N__20935\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__20946\,
            I => \N__20932\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20929\
        );

    \I__4076\ : Odrv12
    port map (
            O => \N__20938\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__4075\ : Odrv4
    port map (
            O => \N__20935\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__4074\ : Odrv12
    port map (
            O => \N__20932\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__20929\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__4072\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20917\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__20917\,
            I => \N__20914\
        );

    \I__4070\ : Span12Mux_h
    port map (
            O => \N__20914\,
            I => \N__20908\
        );

    \I__4069\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20903\
        );

    \I__4068\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20903\
        );

    \I__4067\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20900\
        );

    \I__4066\ : Odrv12
    port map (
            O => \N__20908\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__20903\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__20900\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__20893\,
            I => \N__20890\
        );

    \I__4062\ : InMux
    port map (
            O => \N__20890\,
            I => \N__20887\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__20887\,
            I => \N__20884\
        );

    \I__4060\ : Span12Mux_v
    port map (
            O => \N__20884\,
            I => \N__20881\
        );

    \I__4059\ : Odrv12
    port map (
            O => \N__20881\,
            I => \M_this_vga_signals_address_5\
        );

    \I__4058\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20875\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__20875\,
            I => \N__20872\
        );

    \I__4056\ : Span4Mux_h
    port map (
            O => \N__20872\,
            I => \N__20869\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__20869\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__4054\ : CEMux
    port map (
            O => \N__20866\,
            I => \N__20863\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__20863\,
            I => \N__20859\
        );

    \I__4052\ : CEMux
    port map (
            O => \N__20862\,
            I => \N__20856\
        );

    \I__4051\ : Span4Mux_s3_v
    port map (
            O => \N__20859\,
            I => \N__20851\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__20856\,
            I => \N__20851\
        );

    \I__4049\ : Span4Mux_h
    port map (
            O => \N__20851\,
            I => \N__20848\
        );

    \I__4048\ : Span4Mux_v
    port map (
            O => \N__20848\,
            I => \N__20845\
        );

    \I__4047\ : Span4Mux_v
    port map (
            O => \N__20845\,
            I => \N__20842\
        );

    \I__4046\ : Span4Mux_h
    port map (
            O => \N__20842\,
            I => \N__20839\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__20839\,
            I => \this_sprites_ram.mem_WE_14\
        );

    \I__4044\ : CEMux
    port map (
            O => \N__20836\,
            I => \N__20833\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20829\
        );

    \I__4042\ : CEMux
    port map (
            O => \N__20832\,
            I => \N__20826\
        );

    \I__4041\ : Span4Mux_v
    port map (
            O => \N__20829\,
            I => \N__20821\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__20826\,
            I => \N__20821\
        );

    \I__4039\ : Span4Mux_h
    port map (
            O => \N__20821\,
            I => \N__20818\
        );

    \I__4038\ : Span4Mux_v
    port map (
            O => \N__20818\,
            I => \N__20815\
        );

    \I__4037\ : Span4Mux_h
    port map (
            O => \N__20815\,
            I => \N__20812\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__20812\,
            I => \this_sprites_ram.mem_WE_12\
        );

    \I__4035\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20805\
        );

    \I__4034\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20802\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20795\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__20802\,
            I => \N__20795\
        );

    \I__4031\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20792\
        );

    \I__4030\ : InMux
    port map (
            O => \N__20800\,
            I => \N__20789\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__20795\,
            I => \N__20781\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__20792\,
            I => \N__20781\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__20789\,
            I => \N__20781\
        );

    \I__4026\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20778\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__20781\,
            I => \N__20775\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__20778\,
            I => \N__20772\
        );

    \I__4023\ : Span4Mux_h
    port map (
            O => \N__20775\,
            I => \N__20764\
        );

    \I__4022\ : Span4Mux_v
    port map (
            O => \N__20772\,
            I => \N__20764\
        );

    \I__4021\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20757\
        );

    \I__4020\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20757\
        );

    \I__4019\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20757\
        );

    \I__4018\ : Odrv4
    port map (
            O => \N__20764\,
            I => \M_this_sprites_ram_write_en_0\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__20757\,
            I => \M_this_sprites_ram_write_en_0\
        );

    \I__4016\ : CEMux
    port map (
            O => \N__20752\,
            I => \N__20748\
        );

    \I__4015\ : CEMux
    port map (
            O => \N__20751\,
            I => \N__20745\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__20748\,
            I => \N__20742\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__20745\,
            I => \N__20739\
        );

    \I__4012\ : Span4Mux_h
    port map (
            O => \N__20742\,
            I => \N__20736\
        );

    \I__4011\ : Span4Mux_h
    port map (
            O => \N__20739\,
            I => \N__20733\
        );

    \I__4010\ : Span4Mux_v
    port map (
            O => \N__20736\,
            I => \N__20730\
        );

    \I__4009\ : Span4Mux_h
    port map (
            O => \N__20733\,
            I => \N__20727\
        );

    \I__4008\ : Span4Mux_h
    port map (
            O => \N__20730\,
            I => \N__20724\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__20727\,
            I => \N__20721\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__20724\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__4005\ : Odrv4
    port map (
            O => \N__20721\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__4004\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__20713\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__4002\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20707\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__20707\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__4000\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20701\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__20701\,
            I => \N__20698\
        );

    \I__3998\ : Span4Mux_h
    port map (
            O => \N__20698\,
            I => \N__20695\
        );

    \I__3997\ : Span4Mux_v
    port map (
            O => \N__20695\,
            I => \N__20692\
        );

    \I__3996\ : Span4Mux_h
    port map (
            O => \N__20692\,
            I => \N__20689\
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__20689\,
            I => \this_sprites_ram.mem_out_bus6_1\
        );

    \I__3994\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20683\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__20683\,
            I => \N__20680\
        );

    \I__3992\ : Span4Mux_h
    port map (
            O => \N__20680\,
            I => \N__20677\
        );

    \I__3991\ : Span4Mux_v
    port map (
            O => \N__20677\,
            I => \N__20674\
        );

    \I__3990\ : Span4Mux_v
    port map (
            O => \N__20674\,
            I => \N__20671\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__20671\,
            I => \this_sprites_ram.mem_out_bus2_1\
        );

    \I__3988\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20665\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__20665\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\
        );

    \I__3986\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20659\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__20659\,
            I => \N__20656\
        );

    \I__3984\ : Odrv12
    port map (
            O => \N__20656\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\
        );

    \I__3983\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20650\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__20650\,
            I => \N__20647\
        );

    \I__3981\ : Span4Mux_h
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__3980\ : Odrv4
    port map (
            O => \N__20644\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\
        );

    \I__3979\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20638\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__20638\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2\
        );

    \I__3977\ : InMux
    port map (
            O => \N__20635\,
            I => \N__20632\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__20632\,
            I => \N__20629\
        );

    \I__3975\ : Span4Mux_v
    port map (
            O => \N__20629\,
            I => \N__20626\
        );

    \I__3974\ : Span4Mux_h
    port map (
            O => \N__20626\,
            I => \N__20623\
        );

    \I__3973\ : Span4Mux_h
    port map (
            O => \N__20623\,
            I => \N__20620\
        );

    \I__3972\ : Odrv4
    port map (
            O => \N__20620\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__3971\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20614\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__20614\,
            I => \N__20609\
        );

    \I__3969\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20605\
        );

    \I__3968\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20602\
        );

    \I__3967\ : Span4Mux_h
    port map (
            O => \N__20609\,
            I => \N__20598\
        );

    \I__3966\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20595\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__20605\,
            I => \N__20590\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__20602\,
            I => \N__20590\
        );

    \I__3963\ : InMux
    port map (
            O => \N__20601\,
            I => \N__20587\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__20598\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__20595\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3960\ : Odrv12
    port map (
            O => \N__20590\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__20587\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3958\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20573\
        );

    \I__3957\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20568\
        );

    \I__3956\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20568\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__20573\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__20568\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__3953\ : CEMux
    port map (
            O => \N__20563\,
            I => \N__20560\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__20560\,
            I => \N__20557\
        );

    \I__3951\ : Span4Mux_s2_v
    port map (
            O => \N__20557\,
            I => \N__20553\
        );

    \I__3950\ : CEMux
    port map (
            O => \N__20556\,
            I => \N__20550\
        );

    \I__3949\ : Sp12to4
    port map (
            O => \N__20553\,
            I => \N__20545\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__20550\,
            I => \N__20545\
        );

    \I__3947\ : Span12Mux_v
    port map (
            O => \N__20545\,
            I => \N__20542\
        );

    \I__3946\ : Odrv12
    port map (
            O => \N__20542\,
            I => \this_sprites_ram.mem_WE_0\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__20539\,
            I => \N__20536\
        );

    \I__3944\ : CascadeBuf
    port map (
            O => \N__20536\,
            I => \N__20533\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__20533\,
            I => \N__20530\
        );

    \I__3942\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20526\
        );

    \I__3941\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20522\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__20526\,
            I => \N__20519\
        );

    \I__3939\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20516\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__20522\,
            I => \N__20511\
        );

    \I__3937\ : Span12Mux_s9_v
    port map (
            O => \N__20519\,
            I => \N__20511\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__20516\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__3935\ : Odrv12
    port map (
            O => \N__20511\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__3934\ : CascadeMux
    port map (
            O => \N__20506\,
            I => \N__20503\
        );

    \I__3933\ : CascadeBuf
    port map (
            O => \N__20503\,
            I => \N__20500\
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__20500\,
            I => \N__20497\
        );

    \I__3931\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20494\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__20494\,
            I => \N__20490\
        );

    \I__3929\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20487\
        );

    \I__3928\ : Span4Mux_h
    port map (
            O => \N__20490\,
            I => \N__20484\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__20487\,
            I => \N__20479\
        );

    \I__3926\ : Sp12to4
    port map (
            O => \N__20484\,
            I => \N__20476\
        );

    \I__3925\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20473\
        );

    \I__3924\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20470\
        );

    \I__3923\ : Span4Mux_h
    port map (
            O => \N__20479\,
            I => \N__20467\
        );

    \I__3922\ : Span12Mux_s10_v
    port map (
            O => \N__20476\,
            I => \N__20464\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__20473\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__20470\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__20467\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__3918\ : Odrv12
    port map (
            O => \N__20464\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__20455\,
            I => \N__20452\
        );

    \I__3916\ : CascadeBuf
    port map (
            O => \N__20452\,
            I => \N__20449\
        );

    \I__3915\ : CascadeMux
    port map (
            O => \N__20449\,
            I => \N__20446\
        );

    \I__3914\ : CascadeBuf
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__20443\,
            I => \N__20440\
        );

    \I__3912\ : CascadeBuf
    port map (
            O => \N__20440\,
            I => \N__20437\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__20437\,
            I => \N__20434\
        );

    \I__3910\ : CascadeBuf
    port map (
            O => \N__20434\,
            I => \N__20431\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__20431\,
            I => \N__20428\
        );

    \I__3908\ : CascadeBuf
    port map (
            O => \N__20428\,
            I => \N__20425\
        );

    \I__3907\ : CascadeMux
    port map (
            O => \N__20425\,
            I => \N__20422\
        );

    \I__3906\ : CascadeBuf
    port map (
            O => \N__20422\,
            I => \N__20419\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__20419\,
            I => \N__20416\
        );

    \I__3904\ : CascadeBuf
    port map (
            O => \N__20416\,
            I => \N__20413\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__20413\,
            I => \N__20410\
        );

    \I__3902\ : CascadeBuf
    port map (
            O => \N__20410\,
            I => \N__20407\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__20407\,
            I => \N__20404\
        );

    \I__3900\ : CascadeBuf
    port map (
            O => \N__20404\,
            I => \N__20401\
        );

    \I__3899\ : CascadeMux
    port map (
            O => \N__20401\,
            I => \N__20398\
        );

    \I__3898\ : CascadeBuf
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__20395\,
            I => \N__20392\
        );

    \I__3896\ : CascadeBuf
    port map (
            O => \N__20392\,
            I => \N__20389\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__20389\,
            I => \N__20386\
        );

    \I__3894\ : CascadeBuf
    port map (
            O => \N__20386\,
            I => \N__20383\
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__20383\,
            I => \N__20380\
        );

    \I__3892\ : CascadeBuf
    port map (
            O => \N__20380\,
            I => \N__20377\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__20377\,
            I => \N__20374\
        );

    \I__3890\ : CascadeBuf
    port map (
            O => \N__20374\,
            I => \N__20371\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__20371\,
            I => \N__20368\
        );

    \I__3888\ : CascadeBuf
    port map (
            O => \N__20368\,
            I => \N__20365\
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__20365\,
            I => \N__20361\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__20364\,
            I => \N__20358\
        );

    \I__3885\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20353\
        );

    \I__3884\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20349\
        );

    \I__3883\ : InMux
    port map (
            O => \N__20357\,
            I => \N__20346\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__20356\,
            I => \N__20343\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__20353\,
            I => \N__20340\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__20352\,
            I => \N__20337\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__20349\,
            I => \N__20334\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__20346\,
            I => \N__20331\
        );

    \I__3877\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20328\
        );

    \I__3876\ : Span4Mux_v
    port map (
            O => \N__20340\,
            I => \N__20325\
        );

    \I__3875\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20322\
        );

    \I__3874\ : Span4Mux_h
    port map (
            O => \N__20334\,
            I => \N__20315\
        );

    \I__3873\ : Span4Mux_v
    port map (
            O => \N__20331\,
            I => \N__20315\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__20328\,
            I => \N__20315\
        );

    \I__3871\ : Span4Mux_v
    port map (
            O => \N__20325\,
            I => \N__20312\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__20322\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__20315\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__3868\ : Odrv4
    port map (
            O => \N__20312\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__3867\ : InMux
    port map (
            O => \N__20305\,
            I => \N__20300\
        );

    \I__3866\ : InMux
    port map (
            O => \N__20304\,
            I => \N__20297\
        );

    \I__3865\ : InMux
    port map (
            O => \N__20303\,
            I => \N__20294\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__20300\,
            I => \N__20289\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__20297\,
            I => \N__20289\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__20294\,
            I => \N__20286\
        );

    \I__3861\ : Span4Mux_v
    port map (
            O => \N__20289\,
            I => \N__20283\
        );

    \I__3860\ : Span4Mux_v
    port map (
            O => \N__20286\,
            I => \N__20280\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__20283\,
            I => \this_ppu.un1_M_vaddress_q_c2\
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__20280\,
            I => \this_ppu.un1_M_vaddress_q_c2\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__20275\,
            I => \this_ppu.M_state_q_i_1_cascade_\
        );

    \I__3856\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20269\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__20269\,
            I => \this_ppu.M_last_q_RNIMRAD5_2\
        );

    \I__3854\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20263\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__20263\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_3\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__20260\,
            I => \N__20256\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__20259\,
            I => \N__20253\
        );

    \I__3850\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20250\
        );

    \I__3849\ : InMux
    port map (
            O => \N__20253\,
            I => \N__20247\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__20250\,
            I => \this_ppu.M_count_qZ1Z_3\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__20247\,
            I => \this_ppu.M_count_qZ1Z_3\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__20242\,
            I => \N__20239\
        );

    \I__3845\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20235\
        );

    \I__3844\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20232\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__20235\,
            I => \this_ppu.M_count_qZ1Z_4\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__20232\,
            I => \this_ppu.M_count_qZ1Z_4\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__20227\,
            I => \N__20224\
        );

    \I__3840\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20221\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__20221\,
            I => \N__20217\
        );

    \I__3838\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20214\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__20217\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__20214\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__3835\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20206\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__20206\,
            I => \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4\
        );

    \I__3833\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20199\
        );

    \I__3832\ : InMux
    port map (
            O => \N__20202\,
            I => \N__20196\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__20199\,
            I => \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_5\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__20196\,
            I => \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_5\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__20191\,
            I => \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4_cascade_\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__20188\,
            I => \N__20185\
        );

    \I__3827\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20181\
        );

    \I__3826\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20178\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__20181\,
            I => \N__20170\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20170\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__20177\,
            I => \N__20167\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__20176\,
            I => \N__20164\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__20175\,
            I => \N__20161\
        );

    \I__3820\ : Span4Mux_v
    port map (
            O => \N__20170\,
            I => \N__20156\
        );

    \I__3819\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20153\
        );

    \I__3818\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20150\
        );

    \I__3817\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20145\
        );

    \I__3816\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20145\
        );

    \I__3815\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20142\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__20156\,
            I => \this_ppu.M_state_d_0_sqmuxa_1\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__20153\,
            I => \this_ppu.M_state_d_0_sqmuxa_1\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__20150\,
            I => \this_ppu.M_state_d_0_sqmuxa_1\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__20145\,
            I => \this_ppu.M_state_d_0_sqmuxa_1\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__20142\,
            I => \this_ppu.M_state_d_0_sqmuxa_1\
        );

    \I__3809\ : CascadeMux
    port map (
            O => \N__20131\,
            I => \this_ppu.M_state_d_0_sqmuxa_1_cascade_\
        );

    \I__3808\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20125\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__20125\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_5\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__20122\,
            I => \N__20119\
        );

    \I__3805\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20115\
        );

    \I__3804\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20112\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__20115\,
            I => \this_ppu.M_count_qZ1Z_5\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__20112\,
            I => \this_ppu.M_count_qZ1Z_5\
        );

    \I__3801\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20101\
        );

    \I__3800\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20101\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__20101\,
            I => \N__20088\
        );

    \I__3798\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20081\
        );

    \I__3797\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20081\
        );

    \I__3796\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20081\
        );

    \I__3795\ : InMux
    port map (
            O => \N__20097\,
            I => \N__20078\
        );

    \I__3794\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20075\
        );

    \I__3793\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20072\
        );

    \I__3792\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20069\
        );

    \I__3791\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20062\
        );

    \I__3790\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20062\
        );

    \I__3789\ : InMux
    port map (
            O => \N__20091\,
            I => \N__20062\
        );

    \I__3788\ : Span4Mux_h
    port map (
            O => \N__20088\,
            I => \N__20059\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20056\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__20078\,
            I => \this_ppu.M_state_q_i_1\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__20075\,
            I => \this_ppu.M_state_q_i_1\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__20072\,
            I => \this_ppu.M_state_q_i_1\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__20069\,
            I => \this_ppu.M_state_q_i_1\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__20062\,
            I => \this_ppu.M_state_q_i_1\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__20059\,
            I => \this_ppu.M_state_q_i_1\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__20056\,
            I => \this_ppu.M_state_q_i_1\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__20041\,
            I => \N__20037\
        );

    \I__3778\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20032\
        );

    \I__3777\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20032\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__20032\,
            I => \this_ppu.M_count_qZ0Z_7\
        );

    \I__3775\ : InMux
    port map (
            O => \N__20029\,
            I => \N__20019\
        );

    \I__3774\ : InMux
    port map (
            O => \N__20028\,
            I => \N__20016\
        );

    \I__3773\ : InMux
    port map (
            O => \N__20027\,
            I => \N__20013\
        );

    \I__3772\ : InMux
    port map (
            O => \N__20026\,
            I => \N__20006\
        );

    \I__3771\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20006\
        );

    \I__3770\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20006\
        );

    \I__3769\ : InMux
    port map (
            O => \N__20023\,
            I => \N__20001\
        );

    \I__3768\ : InMux
    port map (
            O => \N__20022\,
            I => \N__20001\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__20019\,
            I => \this_ppu.N_82_i\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__20016\,
            I => \this_ppu.N_82_i\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__20013\,
            I => \this_ppu.N_82_i\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__20006\,
            I => \this_ppu.N_82_i\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__20001\,
            I => \this_ppu.N_82_i\
        );

    \I__3762\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19987\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__19987\,
            I => \this_ppu.un1_M_count_q_1_axb_7\
        );

    \I__3760\ : InMux
    port map (
            O => \N__19984\,
            I => \N__19981\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__19981\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__3758\ : InMux
    port map (
            O => \N__19978\,
            I => \N__19975\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__19975\,
            I => \N__19972\
        );

    \I__3756\ : Span4Mux_h
    port map (
            O => \N__19972\,
            I => \N__19969\
        );

    \I__3755\ : Sp12to4
    port map (
            O => \N__19969\,
            I => \N__19966\
        );

    \I__3754\ : Span12Mux_v
    port map (
            O => \N__19966\,
            I => \N__19963\
        );

    \I__3753\ : Odrv12
    port map (
            O => \N__19963\,
            I => \this_sprites_ram.mem_out_bus6_2\
        );

    \I__3752\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19957\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__19957\,
            I => \N__19954\
        );

    \I__3750\ : Span4Mux_v
    port map (
            O => \N__19954\,
            I => \N__19951\
        );

    \I__3749\ : Sp12to4
    port map (
            O => \N__19951\,
            I => \N__19948\
        );

    \I__3748\ : Odrv12
    port map (
            O => \N__19948\,
            I => \this_sprites_ram.mem_out_bus2_2\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__19945\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_\
        );

    \I__3746\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19939\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__19939\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0\
        );

    \I__3744\ : InMux
    port map (
            O => \N__19936\,
            I => \N__19933\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__19933\,
            I => \N__19930\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__19930\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\
        );

    \I__3741\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19924\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__19924\,
            I => \N__19921\
        );

    \I__3739\ : Span4Mux_v
    port map (
            O => \N__19921\,
            I => \N__19918\
        );

    \I__3738\ : Odrv4
    port map (
            O => \N__19918\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__19915\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\
        );

    \I__3736\ : InMux
    port map (
            O => \N__19912\,
            I => \N__19909\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__19909\,
            I => \N__19906\
        );

    \I__3734\ : Span4Mux_v
    port map (
            O => \N__19906\,
            I => \N__19903\
        );

    \I__3733\ : Sp12to4
    port map (
            O => \N__19903\,
            I => \N__19900\
        );

    \I__3732\ : Odrv12
    port map (
            O => \N__19900\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__3731\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19894\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__19894\,
            I => \N__19891\
        );

    \I__3729\ : Span4Mux_h
    port map (
            O => \N__19891\,
            I => \N__19888\
        );

    \I__3728\ : Span4Mux_h
    port map (
            O => \N__19888\,
            I => \N__19885\
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__19885\,
            I => \this_sprites_ram.mem_out_bus5_1\
        );

    \I__3726\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19879\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__19879\,
            I => \N__19876\
        );

    \I__3724\ : Span4Mux_h
    port map (
            O => \N__19876\,
            I => \N__19873\
        );

    \I__3723\ : Span4Mux_v
    port map (
            O => \N__19873\,
            I => \N__19870\
        );

    \I__3722\ : Span4Mux_v
    port map (
            O => \N__19870\,
            I => \N__19867\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__19867\,
            I => \N__19864\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__19864\,
            I => \this_sprites_ram.mem_out_bus1_1\
        );

    \I__3719\ : InMux
    port map (
            O => \N__19861\,
            I => \N__19858\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__19858\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__19855\,
            I => \this_ppu.N_91_cascade_\
        );

    \I__3716\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19848\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__19851\,
            I => \N__19845\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__19848\,
            I => \N__19842\
        );

    \I__3713\ : InMux
    port map (
            O => \N__19845\,
            I => \N__19839\
        );

    \I__3712\ : Odrv4
    port map (
            O => \N__19842\,
            I => \this_ppu.M_count_qZ1Z_1\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__19839\,
            I => \this_ppu.M_count_qZ1Z_1\
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__19834\,
            I => \N__19830\
        );

    \I__3709\ : InMux
    port map (
            O => \N__19833\,
            I => \N__19827\
        );

    \I__3708\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19824\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__19827\,
            I => \N__19821\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__19824\,
            I => \N__19818\
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__19821\,
            I => \this_ppu.M_count_qZ1Z_2\
        );

    \I__3704\ : Odrv4
    port map (
            O => \N__19818\,
            I => \this_ppu.M_count_qZ1Z_2\
        );

    \I__3703\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19809\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__19812\,
            I => \N__19805\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__19809\,
            I => \N__19802\
        );

    \I__3700\ : InMux
    port map (
            O => \N__19808\,
            I => \N__19799\
        );

    \I__3699\ : InMux
    port map (
            O => \N__19805\,
            I => \N__19796\
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__19802\,
            I => \this_ppu.M_count_qZ1Z_0\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__19799\,
            I => \this_ppu.M_count_qZ1Z_0\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__19796\,
            I => \this_ppu.M_count_qZ1Z_0\
        );

    \I__3695\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19786\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__19786\,
            I => \N__19783\
        );

    \I__3693\ : Span4Mux_v
    port map (
            O => \N__19783\,
            I => \N__19780\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__19780\,
            I => \N__19777\
        );

    \I__3691\ : Sp12to4
    port map (
            O => \N__19777\,
            I => \N__19774\
        );

    \I__3690\ : Span12Mux_h
    port map (
            O => \N__19774\,
            I => \N__19771\
        );

    \I__3689\ : Odrv12
    port map (
            O => \N__19771\,
            I => \this_sprites_ram.mem_out_bus6_0\
        );

    \I__3688\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19765\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__19765\,
            I => \N__19762\
        );

    \I__3686\ : Span4Mux_h
    port map (
            O => \N__19762\,
            I => \N__19759\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__19759\,
            I => \N__19756\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__19756\,
            I => \this_sprites_ram.mem_out_bus2_0\
        );

    \I__3683\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19747\
        );

    \I__3682\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19742\
        );

    \I__3681\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19742\
        );

    \I__3680\ : InMux
    port map (
            O => \N__19750\,
            I => \N__19739\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__19747\,
            I => \N__19736\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__19742\,
            I => \N__19733\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__19739\,
            I => \N__19730\
        );

    \I__3676\ : Span4Mux_h
    port map (
            O => \N__19736\,
            I => \N__19727\
        );

    \I__3675\ : Span4Mux_v
    port map (
            O => \N__19733\,
            I => \N__19724\
        );

    \I__3674\ : Span4Mux_h
    port map (
            O => \N__19730\,
            I => \N__19721\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__19727\,
            I => \this_vga_signals.if_m8_0_a3_1_1_1\
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__19724\,
            I => \this_vga_signals.if_m8_0_a3_1_1_1\
        );

    \I__3671\ : Odrv4
    port map (
            O => \N__19721\,
            I => \this_vga_signals.if_m8_0_a3_1_1_1\
        );

    \I__3670\ : CascadeMux
    port map (
            O => \N__19714\,
            I => \N__19711\
        );

    \I__3669\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19697\
        );

    \I__3668\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19694\
        );

    \I__3667\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19687\
        );

    \I__3666\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19687\
        );

    \I__3665\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19684\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__19706\,
            I => \N__19681\
        );

    \I__3663\ : CascadeMux
    port map (
            O => \N__19705\,
            I => \N__19677\
        );

    \I__3662\ : CascadeMux
    port map (
            O => \N__19704\,
            I => \N__19672\
        );

    \I__3661\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19668\
        );

    \I__3660\ : InMux
    port map (
            O => \N__19702\,
            I => \N__19665\
        );

    \I__3659\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19660\
        );

    \I__3658\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19657\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__19697\,
            I => \N__19652\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__19694\,
            I => \N__19652\
        );

    \I__3655\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19649\
        );

    \I__3654\ : CascadeMux
    port map (
            O => \N__19692\,
            I => \N__19645\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__19687\,
            I => \N__19638\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19635\
        );

    \I__3651\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19630\
        );

    \I__3650\ : InMux
    port map (
            O => \N__19680\,
            I => \N__19630\
        );

    \I__3649\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19625\
        );

    \I__3648\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19625\
        );

    \I__3647\ : InMux
    port map (
            O => \N__19675\,
            I => \N__19618\
        );

    \I__3646\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19618\
        );

    \I__3645\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19618\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__19668\,
            I => \N__19612\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__19665\,
            I => \N__19609\
        );

    \I__3642\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19604\
        );

    \I__3641\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19604\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__19660\,
            I => \N__19601\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__19657\,
            I => \N__19594\
        );

    \I__3638\ : Span4Mux_v
    port map (
            O => \N__19652\,
            I => \N__19594\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__19649\,
            I => \N__19594\
        );

    \I__3636\ : InMux
    port map (
            O => \N__19648\,
            I => \N__19587\
        );

    \I__3635\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19587\
        );

    \I__3634\ : InMux
    port map (
            O => \N__19644\,
            I => \N__19587\
        );

    \I__3633\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19584\
        );

    \I__3632\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19579\
        );

    \I__3631\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19579\
        );

    \I__3630\ : Span4Mux_v
    port map (
            O => \N__19638\,
            I => \N__19574\
        );

    \I__3629\ : Span4Mux_v
    port map (
            O => \N__19635\,
            I => \N__19574\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__19630\,
            I => \N__19567\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__19625\,
            I => \N__19567\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__19618\,
            I => \N__19567\
        );

    \I__3625\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19562\
        );

    \I__3624\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19562\
        );

    \I__3623\ : InMux
    port map (
            O => \N__19615\,
            I => \N__19559\
        );

    \I__3622\ : Span4Mux_h
    port map (
            O => \N__19612\,
            I => \N__19546\
        );

    \I__3621\ : Span4Mux_v
    port map (
            O => \N__19609\,
            I => \N__19546\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__19604\,
            I => \N__19546\
        );

    \I__3619\ : Span4Mux_h
    port map (
            O => \N__19601\,
            I => \N__19546\
        );

    \I__3618\ : Span4Mux_h
    port map (
            O => \N__19594\,
            I => \N__19546\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__19587\,
            I => \N__19546\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__19584\,
            I => \N__19541\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__19579\,
            I => \N__19541\
        );

    \I__3614\ : Odrv4
    port map (
            O => \N__19574\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__3613\ : Odrv12
    port map (
            O => \N__19567\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__19562\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__19559\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__19546\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__3609\ : Odrv12
    port map (
            O => \N__19541\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__3608\ : InMux
    port map (
            O => \N__19528\,
            I => \N__19514\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__19527\,
            I => \N__19509\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__19526\,
            I => \N__19504\
        );

    \I__3605\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19501\
        );

    \I__3604\ : InMux
    port map (
            O => \N__19524\,
            I => \N__19492\
        );

    \I__3603\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19492\
        );

    \I__3602\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19492\
        );

    \I__3601\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19492\
        );

    \I__3600\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19489\
        );

    \I__3599\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19482\
        );

    \I__3598\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19482\
        );

    \I__3597\ : InMux
    port map (
            O => \N__19517\,
            I => \N__19482\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__19514\,
            I => \N__19479\
        );

    \I__3595\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19476\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__19512\,
            I => \N__19467\
        );

    \I__3593\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19464\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__19508\,
            I => \N__19459\
        );

    \I__3591\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19452\
        );

    \I__3590\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19449\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__19501\,
            I => \N__19444\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__19492\,
            I => \N__19444\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19439\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__19482\,
            I => \N__19439\
        );

    \I__3585\ : Span4Mux_v
    port map (
            O => \N__19479\,
            I => \N__19434\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__19476\,
            I => \N__19434\
        );

    \I__3583\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19431\
        );

    \I__3582\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19428\
        );

    \I__3581\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19423\
        );

    \I__3580\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19423\
        );

    \I__3579\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19416\
        );

    \I__3578\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19416\
        );

    \I__3577\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19416\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__19464\,
            I => \N__19413\
        );

    \I__3575\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19410\
        );

    \I__3574\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19403\
        );

    \I__3573\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19403\
        );

    \I__3572\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19403\
        );

    \I__3571\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19396\
        );

    \I__3570\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19396\
        );

    \I__3569\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19396\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__19452\,
            I => \N__19387\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__19449\,
            I => \N__19387\
        );

    \I__3566\ : Span4Mux_v
    port map (
            O => \N__19444\,
            I => \N__19387\
        );

    \I__3565\ : Span4Mux_v
    port map (
            O => \N__19439\,
            I => \N__19387\
        );

    \I__3564\ : Span4Mux_h
    port map (
            O => \N__19434\,
            I => \N__19380\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__19431\,
            I => \N__19380\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__19428\,
            I => \N__19380\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__19423\,
            I => \N__19375\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__19416\,
            I => \N__19375\
        );

    \I__3559\ : Odrv12
    port map (
            O => \N__19413\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__19410\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__19403\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__19396\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__3555\ : Odrv4
    port map (
            O => \N__19387\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__3554\ : Odrv4
    port map (
            O => \N__19380\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__19375\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__19360\,
            I => \N__19357\
        );

    \I__3551\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19353\
        );

    \I__3550\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19350\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__19353\,
            I => \N__19347\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__19350\,
            I => \N__19344\
        );

    \I__3547\ : Span4Mux_h
    port map (
            O => \N__19347\,
            I => \N__19341\
        );

    \I__3546\ : Span4Mux_h
    port map (
            O => \N__19344\,
            I => \N__19338\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__19341\,
            I => \this_vga_signals.if_N_5_0\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__19338\,
            I => \this_vga_signals.if_N_5_0\
        );

    \I__3543\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19330\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__19330\,
            I => \N__19327\
        );

    \I__3541\ : Odrv4
    port map (
            O => \N__19327\,
            I => \this_reset_cond.M_stage_qZ0Z_4\
        );

    \I__3540\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19321\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__19321\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\
        );

    \I__3538\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19315\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__19315\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\
        );

    \I__3536\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19309\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__19309\,
            I => \N__19306\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__19306\,
            I => \N__19303\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__19303\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\
        );

    \I__3532\ : InMux
    port map (
            O => \N__19300\,
            I => \N__19297\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__19297\,
            I => \this_reset_cond.M_stage_qZ0Z_5\
        );

    \I__3530\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19291\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__19291\,
            I => \N__19288\
        );

    \I__3528\ : Span4Mux_v
    port map (
            O => \N__19288\,
            I => \N__19285\
        );

    \I__3527\ : Span4Mux_h
    port map (
            O => \N__19285\,
            I => \N__19282\
        );

    \I__3526\ : Odrv4
    port map (
            O => \N__19282\,
            I => \this_sprites_ram.mem_out_bus4_1\
        );

    \I__3525\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19276\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__19276\,
            I => \N__19273\
        );

    \I__3523\ : Span4Mux_v
    port map (
            O => \N__19273\,
            I => \N__19270\
        );

    \I__3522\ : Sp12to4
    port map (
            O => \N__19270\,
            I => \N__19267\
        );

    \I__3521\ : Span12Mux_h
    port map (
            O => \N__19267\,
            I => \N__19264\
        );

    \I__3520\ : Span12Mux_v
    port map (
            O => \N__19264\,
            I => \N__19261\
        );

    \I__3519\ : Odrv12
    port map (
            O => \N__19261\,
            I => \this_sprites_ram.mem_out_bus0_1\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__19258\,
            I => \N__19250\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__19257\,
            I => \N__19243\
        );

    \I__3516\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19238\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__19255\,
            I => \N__19234\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__19254\,
            I => \N__19225\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__19253\,
            I => \N__19222\
        );

    \I__3512\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19218\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__19249\,
            I => \N__19213\
        );

    \I__3510\ : CascadeMux
    port map (
            O => \N__19248\,
            I => \N__19210\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__19247\,
            I => \N__19207\
        );

    \I__3508\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19204\
        );

    \I__3507\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19198\
        );

    \I__3506\ : InMux
    port map (
            O => \N__19242\,
            I => \N__19193\
        );

    \I__3505\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19193\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__19238\,
            I => \N__19190\
        );

    \I__3503\ : InMux
    port map (
            O => \N__19237\,
            I => \N__19185\
        );

    \I__3502\ : InMux
    port map (
            O => \N__19234\,
            I => \N__19185\
        );

    \I__3501\ : InMux
    port map (
            O => \N__19233\,
            I => \N__19182\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__19232\,
            I => \N__19179\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__19231\,
            I => \N__19176\
        );

    \I__3498\ : InMux
    port map (
            O => \N__19230\,
            I => \N__19173\
        );

    \I__3497\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19170\
        );

    \I__3496\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19167\
        );

    \I__3495\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19164\
        );

    \I__3494\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19159\
        );

    \I__3493\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19159\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__19218\,
            I => \N__19156\
        );

    \I__3491\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19153\
        );

    \I__3490\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19150\
        );

    \I__3489\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19147\
        );

    \I__3488\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19142\
        );

    \I__3487\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19142\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__19204\,
            I => \N__19135\
        );

    \I__3485\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19132\
        );

    \I__3484\ : InMux
    port map (
            O => \N__19202\,
            I => \N__19125\
        );

    \I__3483\ : InMux
    port map (
            O => \N__19201\,
            I => \N__19125\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__19198\,
            I => \N__19122\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__19193\,
            I => \N__19115\
        );

    \I__3480\ : Span4Mux_h
    port map (
            O => \N__19190\,
            I => \N__19115\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__19185\,
            I => \N__19115\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__19182\,
            I => \N__19112\
        );

    \I__3477\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19107\
        );

    \I__3476\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19107\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__19173\,
            I => \N__19104\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__19170\,
            I => \N__19099\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__19167\,
            I => \N__19099\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__19164\,
            I => \N__19094\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__19159\,
            I => \N__19094\
        );

    \I__3470\ : Span4Mux_v
    port map (
            O => \N__19156\,
            I => \N__19089\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__19153\,
            I => \N__19089\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__19150\,
            I => \N__19082\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__19147\,
            I => \N__19082\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__19142\,
            I => \N__19082\
        );

    \I__3465\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19073\
        );

    \I__3464\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19073\
        );

    \I__3463\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19073\
        );

    \I__3462\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19073\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__19135\,
            I => \N__19070\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__19132\,
            I => \N__19067\
        );

    \I__3459\ : InMux
    port map (
            O => \N__19131\,
            I => \N__19064\
        );

    \I__3458\ : InMux
    port map (
            O => \N__19130\,
            I => \N__19061\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__19125\,
            I => \N__19058\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__19122\,
            I => \N__19053\
        );

    \I__3455\ : Span4Mux_v
    port map (
            O => \N__19115\,
            I => \N__19053\
        );

    \I__3454\ : Span4Mux_h
    port map (
            O => \N__19112\,
            I => \N__19048\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__19107\,
            I => \N__19048\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__19104\,
            I => \N__19035\
        );

    \I__3451\ : Span4Mux_v
    port map (
            O => \N__19099\,
            I => \N__19035\
        );

    \I__3450\ : Span4Mux_v
    port map (
            O => \N__19094\,
            I => \N__19035\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__19089\,
            I => \N__19035\
        );

    \I__3448\ : Span4Mux_v
    port map (
            O => \N__19082\,
            I => \N__19035\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__19073\,
            I => \N__19035\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__19070\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__19067\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__19064\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__19061\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__3442\ : Odrv12
    port map (
            O => \N__19058\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__19053\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__19048\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__19035\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__19018\,
            I => \N__19015\
        );

    \I__3437\ : InMux
    port map (
            O => \N__19015\,
            I => \N__19001\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__19014\,
            I => \N__18997\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__19013\,
            I => \N__18992\
        );

    \I__3434\ : InMux
    port map (
            O => \N__19012\,
            I => \N__18986\
        );

    \I__3433\ : InMux
    port map (
            O => \N__19011\,
            I => \N__18986\
        );

    \I__3432\ : InMux
    port map (
            O => \N__19010\,
            I => \N__18979\
        );

    \I__3431\ : InMux
    port map (
            O => \N__19009\,
            I => \N__18979\
        );

    \I__3430\ : InMux
    port map (
            O => \N__19008\,
            I => \N__18979\
        );

    \I__3429\ : InMux
    port map (
            O => \N__19007\,
            I => \N__18973\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__19006\,
            I => \N__18969\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__19005\,
            I => \N__18966\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__19004\,
            I => \N__18961\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__19001\,
            I => \N__18957\
        );

    \I__3424\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18952\
        );

    \I__3423\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18952\
        );

    \I__3422\ : InMux
    port map (
            O => \N__18996\,
            I => \N__18945\
        );

    \I__3421\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18945\
        );

    \I__3420\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18945\
        );

    \I__3419\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18942\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__18986\,
            I => \N__18937\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__18979\,
            I => \N__18937\
        );

    \I__3416\ : InMux
    port map (
            O => \N__18978\,
            I => \N__18930\
        );

    \I__3415\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18930\
        );

    \I__3414\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18930\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__18973\,
            I => \N__18927\
        );

    \I__3412\ : InMux
    port map (
            O => \N__18972\,
            I => \N__18924\
        );

    \I__3411\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18921\
        );

    \I__3410\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18914\
        );

    \I__3409\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18914\
        );

    \I__3408\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18914\
        );

    \I__3407\ : InMux
    port map (
            O => \N__18961\,
            I => \N__18910\
        );

    \I__3406\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18907\
        );

    \I__3405\ : Span4Mux_v
    port map (
            O => \N__18957\,
            I => \N__18904\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__18952\,
            I => \N__18901\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__18945\,
            I => \N__18898\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__18942\,
            I => \N__18895\
        );

    \I__3401\ : Span4Mux_v
    port map (
            O => \N__18937\,
            I => \N__18892\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__18930\,
            I => \N__18883\
        );

    \I__3399\ : Span4Mux_h
    port map (
            O => \N__18927\,
            I => \N__18883\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__18924\,
            I => \N__18883\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__18921\,
            I => \N__18883\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18880\
        );

    \I__3395\ : InMux
    port map (
            O => \N__18913\,
            I => \N__18877\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__18910\,
            I => \N__18872\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__18907\,
            I => \N__18872\
        );

    \I__3392\ : Span4Mux_h
    port map (
            O => \N__18904\,
            I => \N__18865\
        );

    \I__3391\ : Span4Mux_h
    port map (
            O => \N__18901\,
            I => \N__18865\
        );

    \I__3390\ : Span4Mux_v
    port map (
            O => \N__18898\,
            I => \N__18865\
        );

    \I__3389\ : Span4Mux_v
    port map (
            O => \N__18895\,
            I => \N__18858\
        );

    \I__3388\ : Span4Mux_h
    port map (
            O => \N__18892\,
            I => \N__18858\
        );

    \I__3387\ : Span4Mux_v
    port map (
            O => \N__18883\,
            I => \N__18858\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__18880\,
            I => \N__18855\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__18877\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__3384\ : Odrv12
    port map (
            O => \N__18872\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__18865\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__18858\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__18855\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__3380\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18839\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__18843\,
            I => \N__18836\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__18842\,
            I => \N__18831\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__18839\,
            I => \N__18827\
        );

    \I__3376\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18822\
        );

    \I__3375\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18822\
        );

    \I__3374\ : InMux
    port map (
            O => \N__18834\,
            I => \N__18817\
        );

    \I__3373\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18817\
        );

    \I__3372\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18814\
        );

    \I__3371\ : Odrv4
    port map (
            O => \N__18827\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__18822\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__18817\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__18814\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__3367\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18802\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__18802\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0\
        );

    \I__3365\ : InMux
    port map (
            O => \N__18799\,
            I => \N__18796\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__18796\,
            I => \N__18793\
        );

    \I__3363\ : Span4Mux_h
    port map (
            O => \N__18793\,
            I => \N__18790\
        );

    \I__3362\ : Span4Mux_v
    port map (
            O => \N__18790\,
            I => \N__18787\
        );

    \I__3361\ : Span4Mux_h
    port map (
            O => \N__18787\,
            I => \N__18784\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__18784\,
            I => \this_sprites_ram.mem_out_bus4_2\
        );

    \I__3359\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18778\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__18778\,
            I => \N__18775\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__18775\,
            I => \N__18772\
        );

    \I__3356\ : Span4Mux_h
    port map (
            O => \N__18772\,
            I => \N__18769\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__18769\,
            I => \N__18766\
        );

    \I__3354\ : Span4Mux_v
    port map (
            O => \N__18766\,
            I => \N__18763\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__18763\,
            I => \this_sprites_ram.mem_out_bus0_2\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__18760\,
            I => \this_ppu.un1_M_count_q_1_axb_0_cascade_\
        );

    \I__3351\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18754\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__18754\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_6\
        );

    \I__3349\ : InMux
    port map (
            O => \N__18751\,
            I => \N__18747\
        );

    \I__3348\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18744\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__18747\,
            I => \N__18741\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__18744\,
            I => \N__18738\
        );

    \I__3345\ : Span4Mux_v
    port map (
            O => \N__18741\,
            I => \N__18735\
        );

    \I__3344\ : Odrv12
    port map (
            O => \N__18738\,
            I => \this_ppu.line_clk.M_last_qZ0\
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__18735\,
            I => \this_ppu.line_clk.M_last_qZ0\
        );

    \I__3342\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18727\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__18727\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__18724\,
            I => \this_ppu.N_82_i_cascade_\
        );

    \I__3339\ : InMux
    port map (
            O => \N__18721\,
            I => \N__18718\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__18718\,
            I => \this_ppu.M_last_q_RNIMRAD5_3\
        );

    \I__3337\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18712\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__18712\,
            I => \this_reset_cond.M_stage_qZ0Z_3\
        );

    \I__3335\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18706\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18703\
        );

    \I__3333\ : Span4Mux_h
    port map (
            O => \N__18703\,
            I => \N__18700\
        );

    \I__3332\ : Span4Mux_v
    port map (
            O => \N__18700\,
            I => \N__18697\
        );

    \I__3331\ : Span4Mux_h
    port map (
            O => \N__18697\,
            I => \N__18694\
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__18694\,
            I => \this_sprites_ram.mem_out_bus4_0\
        );

    \I__3329\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18688\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__18688\,
            I => \N__18685\
        );

    \I__3327\ : Span4Mux_h
    port map (
            O => \N__18685\,
            I => \N__18682\
        );

    \I__3326\ : Span4Mux_h
    port map (
            O => \N__18682\,
            I => \N__18679\
        );

    \I__3325\ : Span4Mux_v
    port map (
            O => \N__18679\,
            I => \N__18676\
        );

    \I__3324\ : Span4Mux_v
    port map (
            O => \N__18676\,
            I => \N__18673\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__18673\,
            I => \this_sprites_ram.mem_out_bus0_0\
        );

    \I__3322\ : InMux
    port map (
            O => \N__18670\,
            I => \this_ppu.un1_M_count_q_1_cry_2\
        );

    \I__3321\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18664\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__18664\,
            I => \this_ppu.M_last_q_RNIMRAD5_4\
        );

    \I__3319\ : InMux
    port map (
            O => \N__18661\,
            I => \this_ppu.un1_M_count_q_1_cry_3\
        );

    \I__3318\ : InMux
    port map (
            O => \N__18658\,
            I => \this_ppu.un1_M_count_q_1_cry_4\
        );

    \I__3317\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18652\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__18652\,
            I => \this_ppu.M_last_q_RNIMRAD5_5\
        );

    \I__3315\ : InMux
    port map (
            O => \N__18649\,
            I => \this_ppu.un1_M_count_q_1_cry_5\
        );

    \I__3314\ : InMux
    port map (
            O => \N__18646\,
            I => \this_ppu.un1_M_count_q_1_cry_6\
        );

    \I__3313\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18640\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__18640\,
            I => \this_ppu.M_last_q_RNIMRAD5_1\
        );

    \I__3311\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18634\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__18634\,
            I => \this_ppu.M_last_q_RNIMRAD5_0\
        );

    \I__3309\ : InMux
    port map (
            O => \N__18631\,
            I => \N__18628\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__18628\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_4\
        );

    \I__3307\ : InMux
    port map (
            O => \N__18625\,
            I => \N__18622\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__18622\,
            I => \this_vga_signals.i13_mux_0_i\
        );

    \I__3305\ : InMux
    port map (
            O => \N__18619\,
            I => \N__18616\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__18616\,
            I => \N__18613\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__18613\,
            I => \this_vga_signals.if_i1_mux\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__18610\,
            I => \this_vga_signals.g1_0_0_cascade_\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__18607\,
            I => \N__18604\
        );

    \I__3300\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18601\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__18601\,
            I => \N__18598\
        );

    \I__3298\ : Span4Mux_h
    port map (
            O => \N__18598\,
            I => \N__18595\
        );

    \I__3297\ : Span4Mux_h
    port map (
            O => \N__18595\,
            I => \N__18592\
        );

    \I__3296\ : Span4Mux_h
    port map (
            O => \N__18592\,
            I => \N__18589\
        );

    \I__3295\ : Odrv4
    port map (
            O => \N__18589\,
            I => \M_this_vga_signals_address_7\
        );

    \I__3294\ : InMux
    port map (
            O => \N__18586\,
            I => \N__18583\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__18583\,
            I => \N__18580\
        );

    \I__3292\ : Span4Mux_h
    port map (
            O => \N__18580\,
            I => \N__18576\
        );

    \I__3291\ : InMux
    port map (
            O => \N__18579\,
            I => \N__18573\
        );

    \I__3290\ : Span4Mux_v
    port map (
            O => \N__18576\,
            I => \N__18567\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18567\
        );

    \I__3288\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18564\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__18567\,
            I => \N__18561\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__18564\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__18561\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__3284\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18553\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__18553\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_N_4L5_1\
        );

    \I__3282\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18545\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__18549\,
            I => \N__18541\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__18548\,
            I => \N__18538\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__18545\,
            I => \N__18535\
        );

    \I__3278\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18528\
        );

    \I__3277\ : InMux
    port map (
            O => \N__18541\,
            I => \N__18528\
        );

    \I__3276\ : InMux
    port map (
            O => \N__18538\,
            I => \N__18528\
        );

    \I__3275\ : Span4Mux_h
    port map (
            O => \N__18535\,
            I => \N__18523\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__18528\,
            I => \N__18520\
        );

    \I__3273\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18517\
        );

    \I__3272\ : InMux
    port map (
            O => \N__18526\,
            I => \N__18514\
        );

    \I__3271\ : Span4Mux_v
    port map (
            O => \N__18523\,
            I => \N__18506\
        );

    \I__3270\ : Span4Mux_v
    port map (
            O => \N__18520\,
            I => \N__18506\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__18517\,
            I => \N__18506\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__18514\,
            I => \N__18503\
        );

    \I__3267\ : InMux
    port map (
            O => \N__18513\,
            I => \N__18500\
        );

    \I__3266\ : Span4Mux_h
    port map (
            O => \N__18506\,
            I => \N__18497\
        );

    \I__3265\ : Odrv12
    port map (
            O => \N__18503\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__18500\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__3263\ : Odrv4
    port map (
            O => \N__18497\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__18490\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_N_4L5_cascade_\
        );

    \I__3261\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18484\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__18484\,
            I => \this_vga_signals.N_5_i\
        );

    \I__3259\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18478\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__18478\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_0\
        );

    \I__3257\ : InMux
    port map (
            O => \N__18475\,
            I => \N__18472\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__18472\,
            I => \N__18469\
        );

    \I__3255\ : Span12Mux_h
    port map (
            O => \N__18469\,
            I => \N__18466\
        );

    \I__3254\ : Odrv12
    port map (
            O => \N__18466\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__3253\ : InMux
    port map (
            O => \N__18463\,
            I => \N__18460\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__18460\,
            I => \this_ppu.un1_M_count_q_1_cry_0_0_c_RNOZ0\
        );

    \I__3251\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18454\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__18454\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_1\
        );

    \I__3249\ : InMux
    port map (
            O => \N__18451\,
            I => \this_ppu.un1_M_count_q_1_cry_0\
        );

    \I__3248\ : InMux
    port map (
            O => \N__18448\,
            I => \N__18445\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__18445\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_2\
        );

    \I__3246\ : InMux
    port map (
            O => \N__18442\,
            I => \this_ppu.un1_M_count_q_1_cry_1\
        );

    \I__3245\ : InMux
    port map (
            O => \N__18439\,
            I => \N__18436\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__18436\,
            I => \N__18433\
        );

    \I__3243\ : Span4Mux_h
    port map (
            O => \N__18433\,
            I => \N__18430\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__18430\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2_0\
        );

    \I__3241\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18424\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__18424\,
            I => \this_vga_signals.g0_1_1_0\
        );

    \I__3239\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18417\
        );

    \I__3238\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18414\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__18417\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__18414\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__18409\,
            I => \this_vga_signals.g0_1_2_0_cascade_\
        );

    \I__3234\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18403\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__18403\,
            I => \this_vga_signals.g1_3\
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__18400\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_2_cascade_\
        );

    \I__3231\ : InMux
    port map (
            O => \N__18397\,
            I => \N__18386\
        );

    \I__3230\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18381\
        );

    \I__3229\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18381\
        );

    \I__3228\ : InMux
    port map (
            O => \N__18394\,
            I => \N__18378\
        );

    \I__3227\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18373\
        );

    \I__3226\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18373\
        );

    \I__3225\ : InMux
    port map (
            O => \N__18391\,
            I => \N__18363\
        );

    \I__3224\ : InMux
    port map (
            O => \N__18390\,
            I => \N__18363\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__18389\,
            I => \N__18357\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__18386\,
            I => \N__18349\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__18381\,
            I => \N__18349\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__18378\,
            I => \N__18346\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__18373\,
            I => \N__18343\
        );

    \I__3218\ : InMux
    port map (
            O => \N__18372\,
            I => \N__18340\
        );

    \I__3217\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18331\
        );

    \I__3216\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18331\
        );

    \I__3215\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18331\
        );

    \I__3214\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18331\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__18363\,
            I => \N__18324\
        );

    \I__3212\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18321\
        );

    \I__3211\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18316\
        );

    \I__3210\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18316\
        );

    \I__3209\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18311\
        );

    \I__3208\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18311\
        );

    \I__3207\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18306\
        );

    \I__3206\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18306\
        );

    \I__3205\ : Span4Mux_v
    port map (
            O => \N__18349\,
            I => \N__18295\
        );

    \I__3204\ : Span4Mux_h
    port map (
            O => \N__18346\,
            I => \N__18295\
        );

    \I__3203\ : Span4Mux_v
    port map (
            O => \N__18343\,
            I => \N__18295\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__18340\,
            I => \N__18295\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__18331\,
            I => \N__18295\
        );

    \I__3200\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18288\
        );

    \I__3199\ : InMux
    port map (
            O => \N__18329\,
            I => \N__18288\
        );

    \I__3198\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18288\
        );

    \I__3197\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18285\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__18324\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__18321\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__18316\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__18311\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__18306\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__18295\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__18288\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__18285\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3188\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18259\
        );

    \I__3187\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18256\
        );

    \I__3186\ : InMux
    port map (
            O => \N__18266\,
            I => \N__18251\
        );

    \I__3185\ : InMux
    port map (
            O => \N__18265\,
            I => \N__18251\
        );

    \I__3184\ : InMux
    port map (
            O => \N__18264\,
            I => \N__18248\
        );

    \I__3183\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18243\
        );

    \I__3182\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18243\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__18259\,
            I => if_generate_plus_mult1_un68_sum_axb1_520
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__18256\,
            I => if_generate_plus_mult1_un68_sum_axb1_520
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__18251\,
            I => if_generate_plus_mult1_un68_sum_axb1_520
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__18248\,
            I => if_generate_plus_mult1_un68_sum_axb1_520
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__18243\,
            I => if_generate_plus_mult1_un68_sum_axb1_520
        );

    \I__3176\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18225\
        );

    \I__3175\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18222\
        );

    \I__3174\ : InMux
    port map (
            O => \N__18230\,
            I => \N__18214\
        );

    \I__3173\ : InMux
    port map (
            O => \N__18229\,
            I => \N__18209\
        );

    \I__3172\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18209\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__18225\,
            I => \N__18204\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__18222\,
            I => \N__18204\
        );

    \I__3169\ : InMux
    port map (
            O => \N__18221\,
            I => \N__18197\
        );

    \I__3168\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18197\
        );

    \I__3167\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18197\
        );

    \I__3166\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18194\
        );

    \I__3165\ : InMux
    port map (
            O => \N__18217\,
            I => \N__18191\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__18214\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__18209\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__18204\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__18197\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__18194\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__18191\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__18178\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\
        );

    \I__3157\ : InMux
    port map (
            O => \N__18175\,
            I => \N__18172\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__18172\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\
        );

    \I__3155\ : InMux
    port map (
            O => \N__18169\,
            I => \N__18166\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__18166\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_i\
        );

    \I__3153\ : InMux
    port map (
            O => \N__18163\,
            I => \N__18160\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__18160\,
            I => \N__18157\
        );

    \I__3151\ : Span4Mux_h
    port map (
            O => \N__18157\,
            I => \N__18153\
        );

    \I__3150\ : InMux
    port map (
            O => \N__18156\,
            I => \N__18150\
        );

    \I__3149\ : Odrv4
    port map (
            O => \N__18153\,
            I => \this_vga_signals.g2_0_0_0\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__18150\,
            I => \this_vga_signals.g2_0_0_0\
        );

    \I__3147\ : InMux
    port map (
            O => \N__18145\,
            I => \N__18142\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__18142\,
            I => \N__18138\
        );

    \I__3145\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18135\
        );

    \I__3144\ : Odrv12
    port map (
            O => \N__18138\,
            I => \this_vga_signals.g1_1\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__18135\,
            I => \this_vga_signals.g1_1\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__18130\,
            I => \N__18124\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__18129\,
            I => \N__18120\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__18128\,
            I => \N__18117\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__18127\,
            I => \N__18112\
        );

    \I__3138\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18109\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__18123\,
            I => \N__18106\
        );

    \I__3136\ : InMux
    port map (
            O => \N__18120\,
            I => \N__18097\
        );

    \I__3135\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18094\
        );

    \I__3134\ : InMux
    port map (
            O => \N__18116\,
            I => \N__18091\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__18115\,
            I => \N__18085\
        );

    \I__3132\ : InMux
    port map (
            O => \N__18112\,
            I => \N__18080\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__18109\,
            I => \N__18077\
        );

    \I__3130\ : InMux
    port map (
            O => \N__18106\,
            I => \N__18074\
        );

    \I__3129\ : InMux
    port map (
            O => \N__18105\,
            I => \N__18071\
        );

    \I__3128\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18068\
        );

    \I__3127\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18065\
        );

    \I__3126\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18060\
        );

    \I__3125\ : InMux
    port map (
            O => \N__18101\,
            I => \N__18060\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__18100\,
            I => \N__18057\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__18097\,
            I => \N__18054\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__18094\,
            I => \N__18051\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__18091\,
            I => \N__18048\
        );

    \I__3120\ : InMux
    port map (
            O => \N__18090\,
            I => \N__18043\
        );

    \I__3119\ : InMux
    port map (
            O => \N__18089\,
            I => \N__18043\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__18088\,
            I => \N__18039\
        );

    \I__3117\ : InMux
    port map (
            O => \N__18085\,
            I => \N__18035\
        );

    \I__3116\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18032\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__18083\,
            I => \N__18028\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__18080\,
            I => \N__18019\
        );

    \I__3113\ : Span4Mux_v
    port map (
            O => \N__18077\,
            I => \N__18019\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__18074\,
            I => \N__18019\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__18071\,
            I => \N__18014\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__18068\,
            I => \N__18014\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__18065\,
            I => \N__18009\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__18060\,
            I => \N__18009\
        );

    \I__3107\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18006\
        );

    \I__3106\ : Span4Mux_v
    port map (
            O => \N__18054\,
            I => \N__17997\
        );

    \I__3105\ : Span4Mux_v
    port map (
            O => \N__18051\,
            I => \N__17997\
        );

    \I__3104\ : Span4Mux_v
    port map (
            O => \N__18048\,
            I => \N__17997\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__18043\,
            I => \N__17997\
        );

    \I__3102\ : InMux
    port map (
            O => \N__18042\,
            I => \N__17994\
        );

    \I__3101\ : InMux
    port map (
            O => \N__18039\,
            I => \N__17989\
        );

    \I__3100\ : InMux
    port map (
            O => \N__18038\,
            I => \N__17989\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__18035\,
            I => \N__17984\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__18032\,
            I => \N__17984\
        );

    \I__3097\ : InMux
    port map (
            O => \N__18031\,
            I => \N__17981\
        );

    \I__3096\ : InMux
    port map (
            O => \N__18028\,
            I => \N__17978\
        );

    \I__3095\ : InMux
    port map (
            O => \N__18027\,
            I => \N__17973\
        );

    \I__3094\ : InMux
    port map (
            O => \N__18026\,
            I => \N__17973\
        );

    \I__3093\ : Span4Mux_h
    port map (
            O => \N__18019\,
            I => \N__17968\
        );

    \I__3092\ : Span4Mux_h
    port map (
            O => \N__18014\,
            I => \N__17968\
        );

    \I__3091\ : Span4Mux_v
    port map (
            O => \N__18009\,
            I => \N__17963\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__18006\,
            I => \N__17963\
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__17997\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__17994\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__17989\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__17984\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__17981\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__17978\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__17973\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__17968\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__17963\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3080\ : InMux
    port map (
            O => \N__17944\,
            I => \N__17936\
        );

    \I__3079\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17933\
        );

    \I__3078\ : InMux
    port map (
            O => \N__17942\,
            I => \N__17930\
        );

    \I__3077\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17922\
        );

    \I__3076\ : InMux
    port map (
            O => \N__17940\,
            I => \N__17922\
        );

    \I__3075\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17922\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__17936\,
            I => \N__17912\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__17933\,
            I => \N__17907\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__17930\,
            I => \N__17907\
        );

    \I__3071\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17904\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__17922\,
            I => \N__17898\
        );

    \I__3069\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17891\
        );

    \I__3068\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17891\
        );

    \I__3067\ : InMux
    port map (
            O => \N__17919\,
            I => \N__17891\
        );

    \I__3066\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17888\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__17917\,
            I => \N__17884\
        );

    \I__3064\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17880\
        );

    \I__3063\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17877\
        );

    \I__3062\ : Span4Mux_v
    port map (
            O => \N__17912\,
            I => \N__17870\
        );

    \I__3061\ : Span4Mux_v
    port map (
            O => \N__17907\,
            I => \N__17870\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__17904\,
            I => \N__17870\
        );

    \I__3059\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17863\
        );

    \I__3058\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17863\
        );

    \I__3057\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17863\
        );

    \I__3056\ : Span4Mux_h
    port map (
            O => \N__17898\,
            I => \N__17856\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__17891\,
            I => \N__17856\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__17888\,
            I => \N__17856\
        );

    \I__3053\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17849\
        );

    \I__3052\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17849\
        );

    \I__3051\ : InMux
    port map (
            O => \N__17883\,
            I => \N__17849\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__17880\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__17877\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__17870\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__17863\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__17856\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__17849\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3044\ : InMux
    port map (
            O => \N__17836\,
            I => \N__17833\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__17833\,
            I => \N__17830\
        );

    \I__3042\ : Span4Mux_h
    port map (
            O => \N__17830\,
            I => \N__17827\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__17827\,
            I => \this_vga_signals.g1_0_2\
        );

    \I__3040\ : InMux
    port map (
            O => \N__17824\,
            I => \N__17821\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__17821\,
            I => \this_vga_signals.g0_0_0\
        );

    \I__3038\ : InMux
    port map (
            O => \N__17818\,
            I => \N__17814\
        );

    \I__3037\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17808\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__17814\,
            I => \N__17798\
        );

    \I__3035\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17795\
        );

    \I__3034\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17790\
        );

    \I__3033\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17790\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__17808\,
            I => \N__17786\
        );

    \I__3031\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17781\
        );

    \I__3030\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17781\
        );

    \I__3029\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17778\
        );

    \I__3028\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17775\
        );

    \I__3027\ : InMux
    port map (
            O => \N__17803\,
            I => \N__17772\
        );

    \I__3026\ : InMux
    port map (
            O => \N__17802\,
            I => \N__17769\
        );

    \I__3025\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17766\
        );

    \I__3024\ : Span4Mux_v
    port map (
            O => \N__17798\,
            I => \N__17763\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__17795\,
            I => \N__17758\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__17790\,
            I => \N__17758\
        );

    \I__3021\ : InMux
    port map (
            O => \N__17789\,
            I => \N__17755\
        );

    \I__3020\ : Span4Mux_v
    port map (
            O => \N__17786\,
            I => \N__17748\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__17781\,
            I => \N__17748\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__17778\,
            I => \N__17748\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__17775\,
            I => \N__17739\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__17772\,
            I => \N__17739\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__17769\,
            I => \N__17739\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__17766\,
            I => \N__17739\
        );

    \I__3013\ : Span4Mux_h
    port map (
            O => \N__17763\,
            I => \N__17734\
        );

    \I__3012\ : Span4Mux_v
    port map (
            O => \N__17758\,
            I => \N__17734\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__17755\,
            I => \N__17727\
        );

    \I__3010\ : Span4Mux_v
    port map (
            O => \N__17748\,
            I => \N__17727\
        );

    \I__3009\ : Span4Mux_v
    port map (
            O => \N__17739\,
            I => \N__17727\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__17734\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__3007\ : Odrv4
    port map (
            O => \N__17727\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__3006\ : InMux
    port map (
            O => \N__17722\,
            I => \N__17719\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__17719\,
            I => \N__17716\
        );

    \I__3004\ : Odrv12
    port map (
            O => \N__17716\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_0_0_0\
        );

    \I__3003\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17710\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__17710\,
            I => \this_vga_signals.m21_0_1\
        );

    \I__3001\ : InMux
    port map (
            O => \N__17707\,
            I => \N__17704\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__17704\,
            I => \N__17701\
        );

    \I__2999\ : Span4Mux_h
    port map (
            O => \N__17701\,
            I => \N__17698\
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__17698\,
            I => \this_vga_signals.i14_mux_i\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__17695\,
            I => \this_vga_signals.N_25_0_0_cascade_\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__17692\,
            I => \this_vga_signals.M_vcounter_q_RNITP439_0Z0Z_2_cascade_\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__17689\,
            I => \N__17686\
        );

    \I__2994\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17683\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__17683\,
            I => \this_vga_signals.m16_0_1\
        );

    \I__2992\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17669\
        );

    \I__2991\ : InMux
    port map (
            O => \N__17679\,
            I => \N__17666\
        );

    \I__2990\ : InMux
    port map (
            O => \N__17678\,
            I => \N__17659\
        );

    \I__2989\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17659\
        );

    \I__2988\ : InMux
    port map (
            O => \N__17676\,
            I => \N__17659\
        );

    \I__2987\ : InMux
    port map (
            O => \N__17675\,
            I => \N__17654\
        );

    \I__2986\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17651\
        );

    \I__2985\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17641\
        );

    \I__2984\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17641\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__17669\,
            I => \N__17634\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__17666\,
            I => \N__17634\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__17659\,
            I => \N__17634\
        );

    \I__2980\ : InMux
    port map (
            O => \N__17658\,
            I => \N__17629\
        );

    \I__2979\ : InMux
    port map (
            O => \N__17657\,
            I => \N__17629\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__17654\,
            I => \N__17624\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__17651\,
            I => \N__17624\
        );

    \I__2976\ : InMux
    port map (
            O => \N__17650\,
            I => \N__17621\
        );

    \I__2975\ : InMux
    port map (
            O => \N__17649\,
            I => \N__17612\
        );

    \I__2974\ : InMux
    port map (
            O => \N__17648\,
            I => \N__17612\
        );

    \I__2973\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17612\
        );

    \I__2972\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17612\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__17641\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__17634\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__17629\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i
        );

    \I__2968\ : Odrv12
    port map (
            O => \N__17624\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__17621\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__17612\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i
        );

    \I__2965\ : InMux
    port map (
            O => \N__17599\,
            I => \N__17596\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__17596\,
            I => \N__17590\
        );

    \I__2963\ : InMux
    port map (
            O => \N__17595\,
            I => \N__17586\
        );

    \I__2962\ : InMux
    port map (
            O => \N__17594\,
            I => \N__17581\
        );

    \I__2961\ : InMux
    port map (
            O => \N__17593\,
            I => \N__17581\
        );

    \I__2960\ : Span4Mux_h
    port map (
            O => \N__17590\,
            I => \N__17578\
        );

    \I__2959\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17575\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__17586\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__17581\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__17578\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__17575\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__17566\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_cascade_\
        );

    \I__2953\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17560\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__17560\,
            I => \N__17557\
        );

    \I__2951\ : Span4Mux_h
    port map (
            O => \N__17557\,
            I => \N__17554\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__17554\,
            I => \this_vga_signals.g0_12\
        );

    \I__2949\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17548\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__17548\,
            I => \this_vga_signals.M_vcounter_q_RNITP439Z0Z_2\
        );

    \I__2947\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17542\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__17542\,
            I => \N__17539\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__17539\,
            I => \this_vga_signals.g2_1_1\
        );

    \I__2944\ : InMux
    port map (
            O => \N__17536\,
            I => \N__17533\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__17533\,
            I => \this_vga_signals.g1_1_1_0\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__17530\,
            I => \N__17527\
        );

    \I__2941\ : InMux
    port map (
            O => \N__17527\,
            I => \N__17524\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__17524\,
            I => \N__17521\
        );

    \I__2939\ : Odrv4
    port map (
            O => \N__17521\,
            I => \this_vga_signals.if_N_5_1\
        );

    \I__2938\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17515\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__17515\,
            I => \this_vga_signals.g0_5_0\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__17512\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_cascade_\
        );

    \I__2935\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17505\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__17508\,
            I => \N__17502\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__17505\,
            I => \N__17499\
        );

    \I__2932\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17496\
        );

    \I__2931\ : Span4Mux_v
    port map (
            O => \N__17499\,
            I => \N__17491\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__17496\,
            I => \N__17491\
        );

    \I__2929\ : Span4Mux_h
    port map (
            O => \N__17491\,
            I => \N__17488\
        );

    \I__2928\ : Span4Mux_h
    port map (
            O => \N__17488\,
            I => \N__17485\
        );

    \I__2927\ : Odrv4
    port map (
            O => \N__17485\,
            I => \this_vga_signals.vaddress_2_5\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__17482\,
            I => \this_vga_signals.g1_1_0_0_cascade_\
        );

    \I__2925\ : InMux
    port map (
            O => \N__17479\,
            I => \N__17476\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__17476\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_0_0\
        );

    \I__2923\ : InMux
    port map (
            O => \N__17473\,
            I => \N__17470\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__17470\,
            I => \this_vga_signals.g1_2_0_0\
        );

    \I__2921\ : InMux
    port map (
            O => \N__17467\,
            I => \N__17462\
        );

    \I__2920\ : InMux
    port map (
            O => \N__17466\,
            I => \N__17458\
        );

    \I__2919\ : InMux
    port map (
            O => \N__17465\,
            I => \N__17455\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__17462\,
            I => \N__17452\
        );

    \I__2917\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17449\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__17458\,
            I => \this_vga_signals.if_i2_mux\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__17455\,
            I => \this_vga_signals.if_i2_mux\
        );

    \I__2914\ : Odrv4
    port map (
            O => \N__17452\,
            I => \this_vga_signals.if_i2_mux\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__17449\,
            I => \this_vga_signals.if_i2_mux\
        );

    \I__2912\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17437\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__17437\,
            I => \this_vga_signals.M_vcounter_d7lt3\
        );

    \I__2910\ : InMux
    port map (
            O => \N__17434\,
            I => \N__17430\
        );

    \I__2909\ : InMux
    port map (
            O => \N__17433\,
            I => \N__17427\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__17430\,
            I => \N__17424\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__17427\,
            I => \N__17421\
        );

    \I__2906\ : Span4Mux_v
    port map (
            O => \N__17424\,
            I => \N__17416\
        );

    \I__2905\ : Span4Mux_v
    port map (
            O => \N__17421\,
            I => \N__17416\
        );

    \I__2904\ : Span4Mux_h
    port map (
            O => \N__17416\,
            I => \N__17413\
        );

    \I__2903\ : Span4Mux_h
    port map (
            O => \N__17413\,
            I => \N__17410\
        );

    \I__2902\ : Odrv4
    port map (
            O => \N__17410\,
            I => \this_vga_signals.M_vcounter_d7lt9_1\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__17407\,
            I => \this_vga_signals.M_vcounter_d7lt9_1_cascade_\
        );

    \I__2900\ : InMux
    port map (
            O => \N__17404\,
            I => \N__17400\
        );

    \I__2899\ : InMux
    port map (
            O => \N__17403\,
            I => \N__17397\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__17400\,
            I => \N__17394\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__17397\,
            I => \N__17389\
        );

    \I__2896\ : Span4Mux_v
    port map (
            O => \N__17394\,
            I => \N__17389\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__17389\,
            I => \this_vga_signals.un4_lvisibility_1\
        );

    \I__2894\ : InMux
    port map (
            O => \N__17386\,
            I => \N__17383\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__17383\,
            I => \N__17379\
        );

    \I__2892\ : InMux
    port map (
            O => \N__17382\,
            I => \N__17376\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__17379\,
            I => \N__17371\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__17376\,
            I => \N__17371\
        );

    \I__2889\ : Span4Mux_h
    port map (
            O => \N__17371\,
            I => \N__17368\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__17368\,
            I => \this_vga_signals.if_m8_0_a3_1_1_0\
        );

    \I__2887\ : InMux
    port map (
            O => \N__17365\,
            I => \N__17362\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__17362\,
            I => \N__17359\
        );

    \I__2885\ : Span4Mux_v
    port map (
            O => \N__17359\,
            I => \N__17356\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__17356\,
            I => \this_vga_signals.g0_0\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__17353\,
            I => \this_vga_signals.vaddress_1_5_cascade_\
        );

    \I__2882\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17347\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__17347\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_0_1\
        );

    \I__2880\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17332\
        );

    \I__2879\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17327\
        );

    \I__2878\ : InMux
    port map (
            O => \N__17342\,
            I => \N__17324\
        );

    \I__2877\ : InMux
    port map (
            O => \N__17341\,
            I => \N__17319\
        );

    \I__2876\ : InMux
    port map (
            O => \N__17340\,
            I => \N__17319\
        );

    \I__2875\ : InMux
    port map (
            O => \N__17339\,
            I => \N__17314\
        );

    \I__2874\ : InMux
    port map (
            O => \N__17338\,
            I => \N__17314\
        );

    \I__2873\ : InMux
    port map (
            O => \N__17337\,
            I => \N__17307\
        );

    \I__2872\ : InMux
    port map (
            O => \N__17336\,
            I => \N__17307\
        );

    \I__2871\ : InMux
    port map (
            O => \N__17335\,
            I => \N__17307\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__17332\,
            I => \N__17300\
        );

    \I__2869\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17297\
        );

    \I__2868\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17294\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__17327\,
            I => \N__17289\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__17324\,
            I => \N__17289\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17286\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__17314\,
            I => \N__17283\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__17307\,
            I => \N__17280\
        );

    \I__2862\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17275\
        );

    \I__2861\ : InMux
    port map (
            O => \N__17305\,
            I => \N__17275\
        );

    \I__2860\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17270\
        );

    \I__2859\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17270\
        );

    \I__2858\ : Span4Mux_h
    port map (
            O => \N__17300\,
            I => \N__17267\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__17297\,
            I => \N__17260\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__17294\,
            I => \N__17260\
        );

    \I__2855\ : Span4Mux_h
    port map (
            O => \N__17289\,
            I => \N__17260\
        );

    \I__2854\ : Span4Mux_h
    port map (
            O => \N__17286\,
            I => \N__17257\
        );

    \I__2853\ : Odrv12
    port map (
            O => \N__17283\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__17280\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__17275\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__17270\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__17267\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__17260\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__17257\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2846\ : InMux
    port map (
            O => \N__17242\,
            I => \N__17239\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__17239\,
            I => \this_vga_signals.vaddress_1_5\
        );

    \I__2844\ : InMux
    port map (
            O => \N__17236\,
            I => \N__17229\
        );

    \I__2843\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17226\
        );

    \I__2842\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17221\
        );

    \I__2841\ : InMux
    port map (
            O => \N__17233\,
            I => \N__17212\
        );

    \I__2840\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17212\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__17229\,
            I => \N__17208\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__17226\,
            I => \N__17205\
        );

    \I__2837\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17201\
        );

    \I__2836\ : InMux
    port map (
            O => \N__17224\,
            I => \N__17196\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__17221\,
            I => \N__17193\
        );

    \I__2834\ : InMux
    port map (
            O => \N__17220\,
            I => \N__17190\
        );

    \I__2833\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17183\
        );

    \I__2832\ : InMux
    port map (
            O => \N__17218\,
            I => \N__17183\
        );

    \I__2831\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17183\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__17212\,
            I => \N__17180\
        );

    \I__2829\ : InMux
    port map (
            O => \N__17211\,
            I => \N__17167\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__17208\,
            I => \N__17162\
        );

    \I__2827\ : Span4Mux_v
    port map (
            O => \N__17205\,
            I => \N__17162\
        );

    \I__2826\ : InMux
    port map (
            O => \N__17204\,
            I => \N__17159\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__17201\,
            I => \N__17156\
        );

    \I__2824\ : InMux
    port map (
            O => \N__17200\,
            I => \N__17151\
        );

    \I__2823\ : InMux
    port map (
            O => \N__17199\,
            I => \N__17151\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__17196\,
            I => \N__17140\
        );

    \I__2821\ : Span4Mux_h
    port map (
            O => \N__17193\,
            I => \N__17140\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__17190\,
            I => \N__17140\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__17183\,
            I => \N__17140\
        );

    \I__2818\ : Span4Mux_h
    port map (
            O => \N__17180\,
            I => \N__17140\
        );

    \I__2817\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17137\
        );

    \I__2816\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17132\
        );

    \I__2815\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17132\
        );

    \I__2814\ : InMux
    port map (
            O => \N__17176\,
            I => \N__17127\
        );

    \I__2813\ : InMux
    port map (
            O => \N__17175\,
            I => \N__17127\
        );

    \I__2812\ : InMux
    port map (
            O => \N__17174\,
            I => \N__17116\
        );

    \I__2811\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17116\
        );

    \I__2810\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17116\
        );

    \I__2809\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17116\
        );

    \I__2808\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17116\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__17167\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__17162\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__17159\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__17156\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__17151\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__17140\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__17137\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__17132\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__17127\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__17116\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__17095\,
            I => \this_vga_signals.vaddress_2_6_cascade_\
        );

    \I__2796\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17089\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__17089\,
            I => \this_vga_signals.g1_2_0\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__17086\,
            I => \M_this_vga_signals_line_clk_0_cascade_\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__17083\,
            I => \this_ppu.M_state_d_0_sqmuxa_cascade_\
        );

    \I__2792\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17077\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__17077\,
            I => \N__17074\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__17074\,
            I => \N__17071\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__17071\,
            I => \N__17068\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__17068\,
            I => \this_sprites_ram.mem_out_bus5_2\
        );

    \I__2787\ : InMux
    port map (
            O => \N__17065\,
            I => \N__17062\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__17062\,
            I => \N__17059\
        );

    \I__2785\ : Span12Mux_v
    port map (
            O => \N__17059\,
            I => \N__17056\
        );

    \I__2784\ : Odrv12
    port map (
            O => \N__17056\,
            I => \this_sprites_ram.mem_out_bus1_2\
        );

    \I__2783\ : InMux
    port map (
            O => \N__17053\,
            I => \N__17050\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__17050\,
            I => \N__17047\
        );

    \I__2781\ : Span12Mux_v
    port map (
            O => \N__17047\,
            I => \N__17044\
        );

    \I__2780\ : Odrv12
    port map (
            O => \N__17044\,
            I => \this_sprites_ram.mem_out_bus7_1\
        );

    \I__2779\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17038\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__17038\,
            I => \N__17035\
        );

    \I__2777\ : Span12Mux_v
    port map (
            O => \N__17035\,
            I => \N__17032\
        );

    \I__2776\ : Odrv12
    port map (
            O => \N__17032\,
            I => \this_sprites_ram.mem_out_bus3_1\
        );

    \I__2775\ : InMux
    port map (
            O => \N__17029\,
            I => \N__17025\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__17028\,
            I => \N__17022\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__17025\,
            I => \N__17019\
        );

    \I__2772\ : InMux
    port map (
            O => \N__17022\,
            I => \N__17015\
        );

    \I__2771\ : Span4Mux_h
    port map (
            O => \N__17019\,
            I => \N__17012\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__17018\,
            I => \N__17009\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__17015\,
            I => \N__17005\
        );

    \I__2768\ : Span4Mux_v
    port map (
            O => \N__17012\,
            I => \N__17002\
        );

    \I__2767\ : InMux
    port map (
            O => \N__17009\,
            I => \N__16999\
        );

    \I__2766\ : InMux
    port map (
            O => \N__17008\,
            I => \N__16996\
        );

    \I__2765\ : Span4Mux_v
    port map (
            O => \N__17005\,
            I => \N__16993\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__17002\,
            I => \N__16988\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__16999\,
            I => \N__16988\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__16996\,
            I => \N__16985\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__16993\,
            I => \N__16982\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__16988\,
            I => \N__16979\
        );

    \I__2759\ : Odrv12
    port map (
            O => \N__16985\,
            I => this_vga_signals_vvisibility
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__16982\,
            I => this_vga_signals_vvisibility
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__16979\,
            I => this_vga_signals_vvisibility
        );

    \I__2756\ : InMux
    port map (
            O => \N__16972\,
            I => \N__16968\
        );

    \I__2755\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16965\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__16968\,
            I => \N__16962\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__16965\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0\
        );

    \I__2752\ : Odrv4
    port map (
            O => \N__16962\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0\
        );

    \I__2751\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16954\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__16954\,
            I => \N__16951\
        );

    \I__2749\ : Span4Mux_h
    port map (
            O => \N__16951\,
            I => \N__16947\
        );

    \I__2748\ : InMux
    port map (
            O => \N__16950\,
            I => \N__16944\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__16947\,
            I => this_vga_signals_un5_vaddress_g1_1_0
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__16944\,
            I => this_vga_signals_un5_vaddress_g1_1_0
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__16939\,
            I => \N__16936\
        );

    \I__2744\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16933\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__16933\,
            I => \N__16930\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__16930\,
            I => \N__16927\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__16927\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_0\
        );

    \I__2740\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16921\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__16921\,
            I => \this_vga_signals.g1_2\
        );

    \I__2738\ : InMux
    port map (
            O => \N__16918\,
            I => \N__16915\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__16915\,
            I => \this_vga_signals.m21_0_1_1\
        );

    \I__2736\ : InMux
    port map (
            O => \N__16912\,
            I => \N__16909\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__16909\,
            I => \N__16906\
        );

    \I__2734\ : Span4Mux_h
    port map (
            O => \N__16906\,
            I => \N__16903\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__16903\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\
        );

    \I__2732\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16897\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__16897\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\
        );

    \I__2730\ : InMux
    port map (
            O => \N__16894\,
            I => \N__16891\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__16891\,
            I => \N__16888\
        );

    \I__2728\ : Span4Mux_v
    port map (
            O => \N__16888\,
            I => \N__16885\
        );

    \I__2727\ : Sp12to4
    port map (
            O => \N__16885\,
            I => \N__16882\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__16882\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__2725\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16876\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__16876\,
            I => \this_vga_ramdac.m16\
        );

    \I__2723\ : InMux
    port map (
            O => \N__16873\,
            I => \N__16870\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__16870\,
            I => \N__16865\
        );

    \I__2721\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16862\
        );

    \I__2720\ : InMux
    port map (
            O => \N__16868\,
            I => \N__16859\
        );

    \I__2719\ : Span4Mux_v
    port map (
            O => \N__16865\,
            I => \N__16856\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__16862\,
            I => \N__16851\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__16859\,
            I => \N__16848\
        );

    \I__2716\ : Sp12to4
    port map (
            O => \N__16856\,
            I => \N__16845\
        );

    \I__2715\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16840\
        );

    \I__2714\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16840\
        );

    \I__2713\ : Sp12to4
    port map (
            O => \N__16851\,
            I => \N__16837\
        );

    \I__2712\ : Span12Mux_v
    port map (
            O => \N__16848\,
            I => \N__16832\
        );

    \I__2711\ : Span12Mux_s3_h
    port map (
            O => \N__16845\,
            I => \N__16832\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__16840\,
            I => \N__16827\
        );

    \I__2709\ : Span12Mux_v
    port map (
            O => \N__16837\,
            I => \N__16827\
        );

    \I__2708\ : Span12Mux_h
    port map (
            O => \N__16832\,
            I => \N__16824\
        );

    \I__2707\ : Span12Mux_h
    port map (
            O => \N__16827\,
            I => \N__16821\
        );

    \I__2706\ : Odrv12
    port map (
            O => \N__16824\,
            I => \M_this_vram_read_data_2\
        );

    \I__2705\ : Odrv12
    port map (
            O => \N__16821\,
            I => \M_this_vram_read_data_2\
        );

    \I__2704\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16811\
        );

    \I__2703\ : InMux
    port map (
            O => \N__16815\,
            I => \N__16808\
        );

    \I__2702\ : InMux
    port map (
            O => \N__16814\,
            I => \N__16805\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__16811\,
            I => \N__16800\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__16808\,
            I => \N__16795\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__16805\,
            I => \N__16795\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__16804\,
            I => \N__16792\
        );

    \I__2697\ : InMux
    port map (
            O => \N__16803\,
            I => \N__16788\
        );

    \I__2696\ : Span4Mux_v
    port map (
            O => \N__16800\,
            I => \N__16785\
        );

    \I__2695\ : Span4Mux_v
    port map (
            O => \N__16795\,
            I => \N__16782\
        );

    \I__2694\ : InMux
    port map (
            O => \N__16792\,
            I => \N__16777\
        );

    \I__2693\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16777\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__16788\,
            I => \N__16774\
        );

    \I__2691\ : Sp12to4
    port map (
            O => \N__16785\,
            I => \N__16769\
        );

    \I__2690\ : Sp12to4
    port map (
            O => \N__16782\,
            I => \N__16769\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__16777\,
            I => \N__16764\
        );

    \I__2688\ : Span12Mux_v
    port map (
            O => \N__16774\,
            I => \N__16764\
        );

    \I__2687\ : Span12Mux_h
    port map (
            O => \N__16769\,
            I => \N__16761\
        );

    \I__2686\ : Span12Mux_h
    port map (
            O => \N__16764\,
            I => \N__16758\
        );

    \I__2685\ : Odrv12
    port map (
            O => \N__16761\,
            I => \M_this_vram_read_data_1\
        );

    \I__2684\ : Odrv12
    port map (
            O => \N__16758\,
            I => \M_this_vram_read_data_1\
        );

    \I__2683\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16748\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__16752\,
            I => \N__16744\
        );

    \I__2681\ : InMux
    port map (
            O => \N__16751\,
            I => \N__16740\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__16748\,
            I => \N__16736\
        );

    \I__2679\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16733\
        );

    \I__2678\ : InMux
    port map (
            O => \N__16744\,
            I => \N__16728\
        );

    \I__2677\ : InMux
    port map (
            O => \N__16743\,
            I => \N__16728\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__16740\,
            I => \N__16725\
        );

    \I__2675\ : InMux
    port map (
            O => \N__16739\,
            I => \N__16722\
        );

    \I__2674\ : Span4Mux_h
    port map (
            O => \N__16736\,
            I => \N__16717\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__16733\,
            I => \N__16717\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__16728\,
            I => \N__16714\
        );

    \I__2671\ : Span4Mux_h
    port map (
            O => \N__16725\,
            I => \N__16711\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__16722\,
            I => \N__16706\
        );

    \I__2669\ : Span4Mux_h
    port map (
            O => \N__16717\,
            I => \N__16706\
        );

    \I__2668\ : Span4Mux_v
    port map (
            O => \N__16714\,
            I => \N__16701\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__16711\,
            I => \N__16701\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__16706\,
            I => \N__16698\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__16701\,
            I => \N__16695\
        );

    \I__2664\ : Sp12to4
    port map (
            O => \N__16698\,
            I => \N__16692\
        );

    \I__2663\ : Span4Mux_h
    port map (
            O => \N__16695\,
            I => \N__16689\
        );

    \I__2662\ : Span12Mux_v
    port map (
            O => \N__16692\,
            I => \N__16686\
        );

    \I__2661\ : Span4Mux_h
    port map (
            O => \N__16689\,
            I => \N__16683\
        );

    \I__2660\ : Odrv12
    port map (
            O => \N__16686\,
            I => \M_this_vram_read_data_0\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__16683\,
            I => \M_this_vram_read_data_0\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__16678\,
            I => \N__16675\
        );

    \I__2657\ : InMux
    port map (
            O => \N__16675\,
            I => \N__16670\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__16674\,
            I => \N__16667\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__16673\,
            I => \N__16663\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__16670\,
            I => \N__16660\
        );

    \I__2653\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16657\
        );

    \I__2652\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16654\
        );

    \I__2651\ : InMux
    port map (
            O => \N__16663\,
            I => \N__16651\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__16660\,
            I => \N__16646\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__16657\,
            I => \N__16646\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__16654\,
            I => \N__16641\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__16651\,
            I => \N__16636\
        );

    \I__2646\ : Span4Mux_h
    port map (
            O => \N__16646\,
            I => \N__16636\
        );

    \I__2645\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16631\
        );

    \I__2644\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16631\
        );

    \I__2643\ : Span4Mux_v
    port map (
            O => \N__16641\,
            I => \N__16628\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__16636\,
            I => \N__16625\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__16631\,
            I => \N__16622\
        );

    \I__2640\ : Sp12to4
    port map (
            O => \N__16628\,
            I => \N__16619\
        );

    \I__2639\ : Span4Mux_h
    port map (
            O => \N__16625\,
            I => \N__16616\
        );

    \I__2638\ : Span4Mux_h
    port map (
            O => \N__16622\,
            I => \N__16613\
        );

    \I__2637\ : Span12Mux_s4_h
    port map (
            O => \N__16619\,
            I => \N__16610\
        );

    \I__2636\ : Span4Mux_h
    port map (
            O => \N__16616\,
            I => \N__16607\
        );

    \I__2635\ : Sp12to4
    port map (
            O => \N__16613\,
            I => \N__16602\
        );

    \I__2634\ : Span12Mux_h
    port map (
            O => \N__16610\,
            I => \N__16602\
        );

    \I__2633\ : Span4Mux_h
    port map (
            O => \N__16607\,
            I => \N__16599\
        );

    \I__2632\ : Odrv12
    port map (
            O => \N__16602\,
            I => \M_this_vram_read_data_3\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__16599\,
            I => \M_this_vram_read_data_3\
        );

    \I__2630\ : InMux
    port map (
            O => \N__16594\,
            I => \N__16591\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__16591\,
            I => \this_vga_ramdac.i2_mux\
        );

    \I__2628\ : InMux
    port map (
            O => \N__16588\,
            I => \N__16579\
        );

    \I__2627\ : InMux
    port map (
            O => \N__16587\,
            I => \N__16579\
        );

    \I__2626\ : InMux
    port map (
            O => \N__16586\,
            I => \N__16575\
        );

    \I__2625\ : InMux
    port map (
            O => \N__16585\,
            I => \N__16572\
        );

    \I__2624\ : InMux
    port map (
            O => \N__16584\,
            I => \N__16567\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__16579\,
            I => \N__16564\
        );

    \I__2622\ : InMux
    port map (
            O => \N__16578\,
            I => \N__16561\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__16575\,
            I => \N__16557\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__16572\,
            I => \N__16554\
        );

    \I__2619\ : InMux
    port map (
            O => \N__16571\,
            I => \N__16551\
        );

    \I__2618\ : InMux
    port map (
            O => \N__16570\,
            I => \N__16548\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__16567\,
            I => \N__16545\
        );

    \I__2616\ : Span4Mux_v
    port map (
            O => \N__16564\,
            I => \N__16540\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__16561\,
            I => \N__16540\
        );

    \I__2614\ : InMux
    port map (
            O => \N__16560\,
            I => \N__16535\
        );

    \I__2613\ : Span4Mux_v
    port map (
            O => \N__16557\,
            I => \N__16530\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__16554\,
            I => \N__16530\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__16551\,
            I => \N__16525\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16525\
        );

    \I__2609\ : Span4Mux_v
    port map (
            O => \N__16545\,
            I => \N__16520\
        );

    \I__2608\ : Span4Mux_h
    port map (
            O => \N__16540\,
            I => \N__16520\
        );

    \I__2607\ : InMux
    port map (
            O => \N__16539\,
            I => \N__16515\
        );

    \I__2606\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16515\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__16535\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__16530\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2603\ : Odrv12
    port map (
            O => \N__16525\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__16520\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__16515\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__16504\,
            I => \N__16495\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__16503\,
            I => \N__16491\
        );

    \I__2598\ : InMux
    port map (
            O => \N__16502\,
            I => \N__16488\
        );

    \I__2597\ : InMux
    port map (
            O => \N__16501\,
            I => \N__16485\
        );

    \I__2596\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16482\
        );

    \I__2595\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16479\
        );

    \I__2594\ : InMux
    port map (
            O => \N__16498\,
            I => \N__16476\
        );

    \I__2593\ : InMux
    port map (
            O => \N__16495\,
            I => \N__16473\
        );

    \I__2592\ : InMux
    port map (
            O => \N__16494\,
            I => \N__16470\
        );

    \I__2591\ : InMux
    port map (
            O => \N__16491\,
            I => \N__16464\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__16488\,
            I => \N__16461\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__16485\,
            I => \N__16456\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__16482\,
            I => \N__16456\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__16479\,
            I => \N__16449\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__16476\,
            I => \N__16449\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__16473\,
            I => \N__16449\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__16470\,
            I => \N__16446\
        );

    \I__2583\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16443\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__16468\,
            I => \N__16439\
        );

    \I__2581\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16436\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__16464\,
            I => \N__16433\
        );

    \I__2579\ : Span4Mux_h
    port map (
            O => \N__16461\,
            I => \N__16430\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__16456\,
            I => \N__16425\
        );

    \I__2577\ : Span4Mux_v
    port map (
            O => \N__16449\,
            I => \N__16425\
        );

    \I__2576\ : Span4Mux_v
    port map (
            O => \N__16446\,
            I => \N__16420\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__16443\,
            I => \N__16420\
        );

    \I__2574\ : InMux
    port map (
            O => \N__16442\,
            I => \N__16415\
        );

    \I__2573\ : InMux
    port map (
            O => \N__16439\,
            I => \N__16415\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__16436\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__16433\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__16430\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__16425\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2568\ : Odrv4
    port map (
            O => \N__16420\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__16415\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__16402\,
            I => \N__16399\
        );

    \I__2565\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16396\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__16396\,
            I => \N__16392\
        );

    \I__2563\ : InMux
    port map (
            O => \N__16395\,
            I => \N__16389\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__16392\,
            I => \this_vga_signals.line_clk_1\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__16389\,
            I => \this_vga_signals.line_clk_1\
        );

    \I__2560\ : InMux
    port map (
            O => \N__16384\,
            I => \N__16381\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__16381\,
            I => \N__16378\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__16378\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__2557\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16372\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__16372\,
            I => \N__16369\
        );

    \I__2555\ : Odrv4
    port map (
            O => \N__16369\,
            I => \this_vga_signals.g0_2_0_2\
        );

    \I__2554\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16363\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__16363\,
            I => \this_vga_signals.g1_0_0_0_1\
        );

    \I__2552\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16357\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__16357\,
            I => \this_vga_signals.N_51\
        );

    \I__2550\ : InMux
    port map (
            O => \N__16354\,
            I => \N__16351\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__16351\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0\
        );

    \I__2548\ : InMux
    port map (
            O => \N__16348\,
            I => \N__16344\
        );

    \I__2547\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16341\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__16344\,
            I => \N__16338\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__16341\,
            I => \N__16335\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__16338\,
            I => \N__16332\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__16335\,
            I => \this_vga_signals.g2_1\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__16332\,
            I => \this_vga_signals.g2_1\
        );

    \I__2541\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16324\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__16324\,
            I => \N__16321\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__16321\,
            I => \this_vga_signals.g1_0\
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__16318\,
            I => \this_vga_signals.g1_N_4L5_1_cascade_\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__16315\,
            I => \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5EZ0Z1_cascade_\
        );

    \I__2536\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16303\
        );

    \I__2535\ : InMux
    port map (
            O => \N__16311\,
            I => \N__16303\
        );

    \I__2534\ : InMux
    port map (
            O => \N__16310\,
            I => \N__16298\
        );

    \I__2533\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16298\
        );

    \I__2532\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16295\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__16303\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__16298\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__16295\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__2528\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16285\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__16285\,
            I => \this_vga_signals.g0_1_1\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__16282\,
            I => \N__16277\
        );

    \I__2525\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16274\
        );

    \I__2524\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16271\
        );

    \I__2523\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16268\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__16274\,
            I => \this_vga_signals.d_N_3_0_i\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__16271\,
            I => \this_vga_signals.d_N_3_0_i\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__16268\,
            I => \this_vga_signals.d_N_3_0_i\
        );

    \I__2519\ : InMux
    port map (
            O => \N__16261\,
            I => \N__16258\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__16258\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_x0\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__16255\,
            I => \this_vga_signals.mult1_un61_sum_c3_cascade_\
        );

    \I__2516\ : InMux
    port map (
            O => \N__16252\,
            I => \N__16249\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__16249\,
            I => \this_vga_signals.g0_7\
        );

    \I__2514\ : InMux
    port map (
            O => \N__16246\,
            I => \N__16243\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__16243\,
            I => \this_vga_signals.g2_2\
        );

    \I__2512\ : InMux
    port map (
            O => \N__16240\,
            I => \N__16237\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__16237\,
            I => \m18x_N_3LZ0Z3\
        );

    \I__2510\ : InMux
    port map (
            O => \N__16234\,
            I => \N__16231\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__16231\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI5BS7NZ0Z_5\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__16228\,
            I => \N__16225\
        );

    \I__2507\ : InMux
    port map (
            O => \N__16225\,
            I => \N__16221\
        );

    \I__2506\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16218\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__16221\,
            I => \N__16213\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__16218\,
            I => \N__16213\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__16213\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_0_0\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__16210\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0_x0_cascade_\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__16207\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0_cascade_\
        );

    \I__2500\ : InMux
    port map (
            O => \N__16204\,
            I => \N__16201\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__16201\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0_x1\
        );

    \I__2498\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16195\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__16195\,
            I => \N__16192\
        );

    \I__2496\ : Span4Mux_h
    port map (
            O => \N__16192\,
            I => \N__16189\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__16189\,
            I => \N__16186\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__16186\,
            I => \this_vga_signals.vaddress_4_5\
        );

    \I__2493\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16180\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__16180\,
            I => \N__16175\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__16179\,
            I => \N__16172\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__16178\,
            I => \N__16169\
        );

    \I__2489\ : Span4Mux_h
    port map (
            O => \N__16175\,
            I => \N__16163\
        );

    \I__2488\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16158\
        );

    \I__2487\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16158\
        );

    \I__2486\ : InMux
    port map (
            O => \N__16168\,
            I => \N__16155\
        );

    \I__2485\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16150\
        );

    \I__2484\ : InMux
    port map (
            O => \N__16166\,
            I => \N__16150\
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__16163\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__16158\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__16155\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__16150\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__16141\,
            I => \N__16131\
        );

    \I__2478\ : InMux
    port map (
            O => \N__16140\,
            I => \N__16128\
        );

    \I__2477\ : InMux
    port map (
            O => \N__16139\,
            I => \N__16123\
        );

    \I__2476\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16123\
        );

    \I__2475\ : InMux
    port map (
            O => \N__16137\,
            I => \N__16118\
        );

    \I__2474\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16118\
        );

    \I__2473\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16113\
        );

    \I__2472\ : InMux
    port map (
            O => \N__16134\,
            I => \N__16113\
        );

    \I__2471\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16110\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__16128\,
            I => \N__16107\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__16123\,
            I => \N__16104\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__16118\,
            I => \N__16099\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__16113\,
            I => \N__16099\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__16110\,
            I => \N__16092\
        );

    \I__2465\ : Span4Mux_h
    port map (
            O => \N__16107\,
            I => \N__16092\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__16104\,
            I => \N__16092\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__16099\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__16092\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2461\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16084\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__16084\,
            I => \N__16081\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__16081\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_0\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__16078\,
            I => \this_vga_signals.mult1_un47_sum_c3_cascade_\
        );

    \I__2457\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16072\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__16072\,
            I => \this_vga_signals.N_5_i_0_0\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__16069\,
            I => \N__16066\
        );

    \I__2454\ : InMux
    port map (
            O => \N__16066\,
            I => \N__16063\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__16063\,
            I => \this_vga_signals.i2_mux\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__16060\,
            I => \this_vga_signals.i2_mux_cascade_\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__16057\,
            I => \this_vga_signals.if_i2_mux_cascade_\
        );

    \I__2450\ : InMux
    port map (
            O => \N__16054\,
            I => \N__16051\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__16051\,
            I => \N__16047\
        );

    \I__2448\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16044\
        );

    \I__2447\ : Span4Mux_v
    port map (
            O => \N__16047\,
            I => \N__16041\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__16044\,
            I => \N__16036\
        );

    \I__2445\ : Span4Mux_h
    port map (
            O => \N__16041\,
            I => \N__16036\
        );

    \I__2444\ : Odrv4
    port map (
            O => \N__16036\,
            I => \this_vga_signals.vaddress_0_6\
        );

    \I__2443\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16026\
        );

    \I__2442\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16026\
        );

    \I__2441\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16023\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__16026\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__16023\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__2438\ : InMux
    port map (
            O => \N__16018\,
            I => \N__16013\
        );

    \I__2437\ : InMux
    port map (
            O => \N__16017\,
            I => \N__16010\
        );

    \I__2436\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16007\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__16013\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__16010\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__16007\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2432\ : InMux
    port map (
            O => \N__16000\,
            I => \N__15991\
        );

    \I__2431\ : InMux
    port map (
            O => \N__15999\,
            I => \N__15987\
        );

    \I__2430\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15984\
        );

    \I__2429\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15981\
        );

    \I__2428\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15976\
        );

    \I__2427\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15976\
        );

    \I__2426\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15972\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__15991\,
            I => \N__15969\
        );

    \I__2424\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15966\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__15987\,
            I => \N__15961\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__15984\,
            I => \N__15955\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__15981\,
            I => \N__15955\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__15976\,
            I => \N__15952\
        );

    \I__2419\ : InMux
    port map (
            O => \N__15975\,
            I => \N__15949\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__15972\,
            I => \N__15942\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__15969\,
            I => \N__15942\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__15966\,
            I => \N__15942\
        );

    \I__2415\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15939\
        );

    \I__2414\ : InMux
    port map (
            O => \N__15964\,
            I => \N__15932\
        );

    \I__2413\ : Span12Mux_v
    port map (
            O => \N__15961\,
            I => \N__15929\
        );

    \I__2412\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15926\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__15955\,
            I => \N__15921\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__15952\,
            I => \N__15921\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__15949\,
            I => \N__15914\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__15942\,
            I => \N__15914\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__15939\,
            I => \N__15914\
        );

    \I__2406\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15911\
        );

    \I__2405\ : InMux
    port map (
            O => \N__15937\,
            I => \N__15908\
        );

    \I__2404\ : InMux
    port map (
            O => \N__15936\,
            I => \N__15903\
        );

    \I__2403\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15903\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__15932\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2401\ : Odrv12
    port map (
            O => \N__15929\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__15926\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__15921\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__15914\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__15911\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__15908\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__15903\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2394\ : InMux
    port map (
            O => \N__15886\,
            I => \N__15882\
        );

    \I__2393\ : InMux
    port map (
            O => \N__15885\,
            I => \N__15879\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__15882\,
            I => \N__15876\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__15879\,
            I => \N__15871\
        );

    \I__2390\ : Span4Mux_v
    port map (
            O => \N__15876\,
            I => \N__15868\
        );

    \I__2389\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15863\
        );

    \I__2388\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15863\
        );

    \I__2387\ : Span12Mux_s5_h
    port map (
            O => \N__15871\,
            I => \N__15858\
        );

    \I__2386\ : Span4Mux_h
    port map (
            O => \N__15868\,
            I => \N__15853\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__15863\,
            I => \N__15853\
        );

    \I__2384\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15848\
        );

    \I__2383\ : InMux
    port map (
            O => \N__15861\,
            I => \N__15848\
        );

    \I__2382\ : Odrv12
    port map (
            O => \N__15858\,
            I => \G_384\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__15853\,
            I => \G_384\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__15848\,
            I => \G_384\
        );

    \I__2379\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15838\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__15838\,
            I => \N__15835\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__15835\,
            I => \N__15831\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__15834\,
            I => \N__15828\
        );

    \I__2375\ : Span4Mux_h
    port map (
            O => \N__15831\,
            I => \N__15825\
        );

    \I__2374\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15822\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__15825\,
            I => \this_vga_ramdac.N_2873_reto\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__15822\,
            I => \this_vga_ramdac.N_2873_reto\
        );

    \I__2371\ : InMux
    port map (
            O => \N__15817\,
            I => \N__15811\
        );

    \I__2370\ : InMux
    port map (
            O => \N__15816\,
            I => \N__15811\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__15811\,
            I => \N_3_0\
        );

    \I__2368\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15802\
        );

    \I__2367\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15802\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__15802\,
            I => \N_2_0\
        );

    \I__2365\ : InMux
    port map (
            O => \N__15799\,
            I => \N__15796\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__15796\,
            I => \M_this_vga_signals_pixel_clk_0_0\
        );

    \I__2363\ : CEMux
    port map (
            O => \N__15793\,
            I => \N__15789\
        );

    \I__2362\ : CEMux
    port map (
            O => \N__15792\,
            I => \N__15786\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__15789\,
            I => \N__15783\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__15786\,
            I => \N__15780\
        );

    \I__2359\ : Span4Mux_v
    port map (
            O => \N__15783\,
            I => \N__15777\
        );

    \I__2358\ : Span4Mux_h
    port map (
            O => \N__15780\,
            I => \N__15774\
        );

    \I__2357\ : Span4Mux_v
    port map (
            O => \N__15777\,
            I => \N__15771\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__15774\,
            I => \N__15768\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__15771\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__15768\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__15763\,
            I => \N__15760\
        );

    \I__2352\ : CascadeBuf
    port map (
            O => \N__15760\,
            I => \N__15757\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__15757\,
            I => \N__15754\
        );

    \I__2350\ : CascadeBuf
    port map (
            O => \N__15754\,
            I => \N__15751\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__15751\,
            I => \N__15748\
        );

    \I__2348\ : CascadeBuf
    port map (
            O => \N__15748\,
            I => \N__15745\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__15745\,
            I => \N__15742\
        );

    \I__2346\ : CascadeBuf
    port map (
            O => \N__15742\,
            I => \N__15739\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__15739\,
            I => \N__15736\
        );

    \I__2344\ : CascadeBuf
    port map (
            O => \N__15736\,
            I => \N__15733\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__15733\,
            I => \N__15730\
        );

    \I__2342\ : CascadeBuf
    port map (
            O => \N__15730\,
            I => \N__15727\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__15727\,
            I => \N__15724\
        );

    \I__2340\ : CascadeBuf
    port map (
            O => \N__15724\,
            I => \N__15721\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__15721\,
            I => \N__15718\
        );

    \I__2338\ : CascadeBuf
    port map (
            O => \N__15718\,
            I => \N__15715\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__15715\,
            I => \N__15712\
        );

    \I__2336\ : CascadeBuf
    port map (
            O => \N__15712\,
            I => \N__15709\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__15709\,
            I => \N__15706\
        );

    \I__2334\ : CascadeBuf
    port map (
            O => \N__15706\,
            I => \N__15703\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__15703\,
            I => \N__15700\
        );

    \I__2332\ : CascadeBuf
    port map (
            O => \N__15700\,
            I => \N__15697\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__15697\,
            I => \N__15694\
        );

    \I__2330\ : CascadeBuf
    port map (
            O => \N__15694\,
            I => \N__15691\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__15691\,
            I => \N__15688\
        );

    \I__2328\ : CascadeBuf
    port map (
            O => \N__15688\,
            I => \N__15685\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__15685\,
            I => \N__15682\
        );

    \I__2326\ : CascadeBuf
    port map (
            O => \N__15682\,
            I => \N__15678\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__15681\,
            I => \N__15675\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__15678\,
            I => \N__15672\
        );

    \I__2323\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15669\
        );

    \I__2322\ : CascadeBuf
    port map (
            O => \N__15672\,
            I => \N__15666\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__15669\,
            I => \N__15663\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__15666\,
            I => \N__15660\
        );

    \I__2319\ : Span4Mux_v
    port map (
            O => \N__15663\,
            I => \N__15656\
        );

    \I__2318\ : InMux
    port map (
            O => \N__15660\,
            I => \N__15652\
        );

    \I__2317\ : InMux
    port map (
            O => \N__15659\,
            I => \N__15649\
        );

    \I__2316\ : Sp12to4
    port map (
            O => \N__15656\,
            I => \N__15644\
        );

    \I__2315\ : InMux
    port map (
            O => \N__15655\,
            I => \N__15641\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__15652\,
            I => \N__15638\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__15649\,
            I => \N__15635\
        );

    \I__2312\ : InMux
    port map (
            O => \N__15648\,
            I => \N__15630\
        );

    \I__2311\ : InMux
    port map (
            O => \N__15647\,
            I => \N__15630\
        );

    \I__2310\ : Span12Mux_h
    port map (
            O => \N__15644\,
            I => \N__15627\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__15641\,
            I => \N__15622\
        );

    \I__2308\ : Span12Mux_s10_h
    port map (
            O => \N__15638\,
            I => \N__15622\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__15635\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__15630\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__2305\ : Odrv12
    port map (
            O => \N__15627\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__2304\ : Odrv12
    port map (
            O => \N__15622\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__15613\,
            I => \N__15610\
        );

    \I__2302\ : CascadeBuf
    port map (
            O => \N__15610\,
            I => \N__15607\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__15607\,
            I => \N__15604\
        );

    \I__2300\ : CascadeBuf
    port map (
            O => \N__15604\,
            I => \N__15601\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__15601\,
            I => \N__15598\
        );

    \I__2298\ : CascadeBuf
    port map (
            O => \N__15598\,
            I => \N__15595\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__15595\,
            I => \N__15592\
        );

    \I__2296\ : CascadeBuf
    port map (
            O => \N__15592\,
            I => \N__15589\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__15589\,
            I => \N__15586\
        );

    \I__2294\ : CascadeBuf
    port map (
            O => \N__15586\,
            I => \N__15583\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__15583\,
            I => \N__15580\
        );

    \I__2292\ : CascadeBuf
    port map (
            O => \N__15580\,
            I => \N__15577\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__15577\,
            I => \N__15574\
        );

    \I__2290\ : CascadeBuf
    port map (
            O => \N__15574\,
            I => \N__15571\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__15571\,
            I => \N__15568\
        );

    \I__2288\ : CascadeBuf
    port map (
            O => \N__15568\,
            I => \N__15565\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__15565\,
            I => \N__15562\
        );

    \I__2286\ : CascadeBuf
    port map (
            O => \N__15562\,
            I => \N__15559\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__15559\,
            I => \N__15556\
        );

    \I__2284\ : CascadeBuf
    port map (
            O => \N__15556\,
            I => \N__15553\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__15553\,
            I => \N__15550\
        );

    \I__2282\ : CascadeBuf
    port map (
            O => \N__15550\,
            I => \N__15547\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__15547\,
            I => \N__15544\
        );

    \I__2280\ : CascadeBuf
    port map (
            O => \N__15544\,
            I => \N__15541\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__15541\,
            I => \N__15538\
        );

    \I__2278\ : CascadeBuf
    port map (
            O => \N__15538\,
            I => \N__15535\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__15535\,
            I => \N__15532\
        );

    \I__2276\ : CascadeBuf
    port map (
            O => \N__15532\,
            I => \N__15529\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__15529\,
            I => \N__15526\
        );

    \I__2274\ : CascadeBuf
    port map (
            O => \N__15526\,
            I => \N__15523\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__15523\,
            I => \N__15520\
        );

    \I__2272\ : InMux
    port map (
            O => \N__15520\,
            I => \N__15517\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__15517\,
            I => \N__15514\
        );

    \I__2270\ : Span4Mux_h
    port map (
            O => \N__15514\,
            I => \N__15509\
        );

    \I__2269\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15506\
        );

    \I__2268\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15502\
        );

    \I__2267\ : Span4Mux_v
    port map (
            O => \N__15509\,
            I => \N__15499\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__15506\,
            I => \N__15496\
        );

    \I__2265\ : InMux
    port map (
            O => \N__15505\,
            I => \N__15493\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__15502\,
            I => \N__15488\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__15499\,
            I => \N__15488\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__15496\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__15493\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__15488\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__2259\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15478\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__15478\,
            I => \this_vga_signals.g0_2_0_2_x1\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__15475\,
            I => \this_vga_signals.g0_2_0_2_x0_cascade_\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__15472\,
            I => \this_vga_signals.g0_2_0_2_cascade_\
        );

    \I__2255\ : InMux
    port map (
            O => \N__15469\,
            I => \N__15466\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__15466\,
            I => \N__15463\
        );

    \I__2253\ : Span4Mux_v
    port map (
            O => \N__15463\,
            I => \N__15460\
        );

    \I__2252\ : Sp12to4
    port map (
            O => \N__15460\,
            I => \N__15457\
        );

    \I__2251\ : Span12Mux_v
    port map (
            O => \N__15457\,
            I => \N__15454\
        );

    \I__2250\ : Odrv12
    port map (
            O => \N__15454\,
            I => \this_sprites_ram.mem_out_bus7_2\
        );

    \I__2249\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15448\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__15448\,
            I => \N__15445\
        );

    \I__2247\ : Span4Mux_v
    port map (
            O => \N__15445\,
            I => \N__15442\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__15442\,
            I => \N__15439\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__15439\,
            I => \this_sprites_ram.mem_out_bus3_2\
        );

    \I__2244\ : InMux
    port map (
            O => \N__15436\,
            I => \N__15433\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__15433\,
            I => \N__15430\
        );

    \I__2242\ : Span4Mux_h
    port map (
            O => \N__15430\,
            I => \N__15427\
        );

    \I__2241\ : Span4Mux_v
    port map (
            O => \N__15427\,
            I => \N__15424\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__15424\,
            I => \this_sprites_ram.mem_out_bus5_0\
        );

    \I__2239\ : InMux
    port map (
            O => \N__15421\,
            I => \N__15418\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__15418\,
            I => \N__15415\
        );

    \I__2237\ : Span4Mux_h
    port map (
            O => \N__15415\,
            I => \N__15412\
        );

    \I__2236\ : Span4Mux_v
    port map (
            O => \N__15412\,
            I => \N__15409\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__15409\,
            I => \N__15406\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__15406\,
            I => \this_sprites_ram.mem_out_bus1_0\
        );

    \I__2233\ : CEMux
    port map (
            O => \N__15403\,
            I => \N__15399\
        );

    \I__2232\ : CEMux
    port map (
            O => \N__15402\,
            I => \N__15396\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__15399\,
            I => \N__15393\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__15396\,
            I => \N__15390\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__15393\,
            I => \N__15387\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__15390\,
            I => \N__15384\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__15387\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__15384\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__2225\ : InMux
    port map (
            O => \N__15379\,
            I => \N__15376\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__15376\,
            I => \this_vga_ramdac.m6\
        );

    \I__2223\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15370\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__15370\,
            I => \N__15366\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__15369\,
            I => \N__15363\
        );

    \I__2220\ : Span12Mux_s6_h
    port map (
            O => \N__15366\,
            I => \N__15360\
        );

    \I__2219\ : InMux
    port map (
            O => \N__15363\,
            I => \N__15357\
        );

    \I__2218\ : Odrv12
    port map (
            O => \N__15360\,
            I => \this_vga_ramdac.N_2871_reto\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__15357\,
            I => \this_vga_ramdac.N_2871_reto\
        );

    \I__2216\ : CascadeMux
    port map (
            O => \N__15352\,
            I => \G_384_cascade_\
        );

    \I__2215\ : InMux
    port map (
            O => \N__15349\,
            I => \N__15346\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__15346\,
            I => \N__15343\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__15343\,
            I => \N__15340\
        );

    \I__2212\ : Span4Mux_h
    port map (
            O => \N__15340\,
            I => \N__15336\
        );

    \I__2211\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15333\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__15336\,
            I => \this_vga_ramdac.N_2872_reto\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__15333\,
            I => \this_vga_ramdac.N_2872_reto\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__15328\,
            I => \this_vga_signals.if_N_5_cascade_\
        );

    \I__2207\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15319\
        );

    \I__2206\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15314\
        );

    \I__2205\ : InMux
    port map (
            O => \N__15323\,
            I => \N__15314\
        );

    \I__2204\ : InMux
    port map (
            O => \N__15322\,
            I => \N__15311\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__15319\,
            I => \N__15305\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__15314\,
            I => \N__15300\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__15311\,
            I => \N__15300\
        );

    \I__2200\ : InMux
    port map (
            O => \N__15310\,
            I => \N__15297\
        );

    \I__2199\ : InMux
    port map (
            O => \N__15309\,
            I => \N__15292\
        );

    \I__2198\ : InMux
    port map (
            O => \N__15308\,
            I => \N__15292\
        );

    \I__2197\ : Span4Mux_h
    port map (
            O => \N__15305\,
            I => \N__15285\
        );

    \I__2196\ : Span4Mux_v
    port map (
            O => \N__15300\,
            I => \N__15285\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__15297\,
            I => \N__15280\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__15292\,
            I => \N__15280\
        );

    \I__2193\ : InMux
    port map (
            O => \N__15291\,
            I => \N__15275\
        );

    \I__2192\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15275\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__15285\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__15280\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__15275\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__15268\,
            I => \this_vga_signals.vaddress_5_cascade_\
        );

    \I__2187\ : InMux
    port map (
            O => \N__15265\,
            I => \N__15261\
        );

    \I__2186\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15258\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__15261\,
            I => \this_vga_signals.g1_0_0_0\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__15258\,
            I => \this_vga_signals.g1_0_0_0\
        );

    \I__2183\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15250\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__15250\,
            I => \this_vga_signals.g0_1_2_0_1\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__15247\,
            I => \this_vga_signals.g0_1_2_cascade_\
        );

    \I__2180\ : InMux
    port map (
            O => \N__15244\,
            I => \N__15241\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__15241\,
            I => \this_vga_signals.g1_0_1_0_0\
        );

    \I__2178\ : InMux
    port map (
            O => \N__15238\,
            I => \N__15235\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__15235\,
            I => \N__15232\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__15232\,
            I => \this_vga_signals.g2_0\
        );

    \I__2175\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15226\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__15226\,
            I => \N__15223\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__15223\,
            I => \N__15220\
        );

    \I__2172\ : Span4Mux_h
    port map (
            O => \N__15220\,
            I => \N__15217\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__15217\,
            I => \this_vga_signals.g1_1_1\
        );

    \I__2170\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15211\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__15211\,
            I => \this_vga_signals.N_5_i_0\
        );

    \I__2168\ : InMux
    port map (
            O => \N__15208\,
            I => \N__15205\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__15205\,
            I => \this_vga_signals.N_50\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__15202\,
            I => \this_vga_signals.vaddress_1_6_cascade_\
        );

    \I__2165\ : InMux
    port map (
            O => \N__15199\,
            I => \N__15196\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__15196\,
            I => \N__15193\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__15193\,
            I => \N__15190\
        );

    \I__2162\ : Odrv4
    port map (
            O => \N__15190\,
            I => \this_vga_signals.if_m8_0_a3_1_1_3\
        );

    \I__2161\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15184\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__15184\,
            I => \N__15179\
        );

    \I__2159\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15174\
        );

    \I__2158\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15174\
        );

    \I__2157\ : Span4Mux_v
    port map (
            O => \N__15179\,
            I => \N__15169\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__15174\,
            I => \N__15169\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__15169\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__2154\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15163\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__15163\,
            I => \N__15160\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__15160\,
            I => \N__15155\
        );

    \I__2151\ : InMux
    port map (
            O => \N__15159\,
            I => \N__15150\
        );

    \I__2150\ : InMux
    port map (
            O => \N__15158\,
            I => \N__15150\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__15155\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__15150\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__2147\ : CEMux
    port map (
            O => \N__15145\,
            I => \N__15121\
        );

    \I__2146\ : CEMux
    port map (
            O => \N__15144\,
            I => \N__15121\
        );

    \I__2145\ : CEMux
    port map (
            O => \N__15143\,
            I => \N__15121\
        );

    \I__2144\ : CEMux
    port map (
            O => \N__15142\,
            I => \N__15121\
        );

    \I__2143\ : CEMux
    port map (
            O => \N__15141\,
            I => \N__15121\
        );

    \I__2142\ : CEMux
    port map (
            O => \N__15140\,
            I => \N__15121\
        );

    \I__2141\ : CEMux
    port map (
            O => \N__15139\,
            I => \N__15121\
        );

    \I__2140\ : CEMux
    port map (
            O => \N__15138\,
            I => \N__15121\
        );

    \I__2139\ : GlobalMux
    port map (
            O => \N__15121\,
            I => \N__15118\
        );

    \I__2138\ : gio2CtrlBuf
    port map (
            O => \N__15118\,
            I => \this_vga_signals.N_614_1_g\
        );

    \I__2137\ : SRMux
    port map (
            O => \N__15115\,
            I => \N__15088\
        );

    \I__2136\ : SRMux
    port map (
            O => \N__15114\,
            I => \N__15088\
        );

    \I__2135\ : SRMux
    port map (
            O => \N__15113\,
            I => \N__15088\
        );

    \I__2134\ : SRMux
    port map (
            O => \N__15112\,
            I => \N__15088\
        );

    \I__2133\ : SRMux
    port map (
            O => \N__15111\,
            I => \N__15088\
        );

    \I__2132\ : SRMux
    port map (
            O => \N__15110\,
            I => \N__15088\
        );

    \I__2131\ : SRMux
    port map (
            O => \N__15109\,
            I => \N__15088\
        );

    \I__2130\ : SRMux
    port map (
            O => \N__15108\,
            I => \N__15088\
        );

    \I__2129\ : SRMux
    port map (
            O => \N__15107\,
            I => \N__15088\
        );

    \I__2128\ : GlobalMux
    port map (
            O => \N__15088\,
            I => \N__15085\
        );

    \I__2127\ : gio2CtrlBuf
    port map (
            O => \N__15085\,
            I => \this_vga_signals.N_931_g\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__15082\,
            I => \N__15078\
        );

    \I__2125\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15073\
        );

    \I__2124\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15067\
        );

    \I__2123\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15067\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__15076\,
            I => \N__15061\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__15073\,
            I => \N__15057\
        );

    \I__2120\ : InMux
    port map (
            O => \N__15072\,
            I => \N__15054\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__15067\,
            I => \N__15051\
        );

    \I__2118\ : InMux
    port map (
            O => \N__15066\,
            I => \N__15048\
        );

    \I__2117\ : InMux
    port map (
            O => \N__15065\,
            I => \N__15045\
        );

    \I__2116\ : InMux
    port map (
            O => \N__15064\,
            I => \N__15040\
        );

    \I__2115\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15040\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__15060\,
            I => \N__15036\
        );

    \I__2113\ : Span4Mux_v
    port map (
            O => \N__15057\,
            I => \N__15031\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__15054\,
            I => \N__15031\
        );

    \I__2111\ : Span4Mux_v
    port map (
            O => \N__15051\,
            I => \N__15022\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__15048\,
            I => \N__15022\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__15045\,
            I => \N__15022\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__15040\,
            I => \N__15022\
        );

    \I__2107\ : InMux
    port map (
            O => \N__15039\,
            I => \N__15017\
        );

    \I__2106\ : InMux
    port map (
            O => \N__15036\,
            I => \N__15017\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__15031\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__15022\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__15017\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__15010\,
            I => \this_vga_signals.if_m8_0_a3_1_1_1_cascade_\
        );

    \I__2101\ : InMux
    port map (
            O => \N__15007\,
            I => \N__15004\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__15004\,
            I => \this_vga_signals.mult1_un40_sum_axb1_0\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__15001\,
            I => \this_vga_signals.SUM_2_i_1_2_3_cascade_\
        );

    \I__2098\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14995\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__14995\,
            I => \N__14988\
        );

    \I__2096\ : InMux
    port map (
            O => \N__14994\,
            I => \N__14983\
        );

    \I__2095\ : InMux
    port map (
            O => \N__14993\,
            I => \N__14983\
        );

    \I__2094\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14978\
        );

    \I__2093\ : InMux
    port map (
            O => \N__14991\,
            I => \N__14978\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__14988\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__14983\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__14978\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__14971\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_\
        );

    \I__2088\ : InMux
    port map (
            O => \N__14968\,
            I => \N__14962\
        );

    \I__2087\ : InMux
    port map (
            O => \N__14967\,
            I => \N__14959\
        );

    \I__2086\ : InMux
    port map (
            O => \N__14966\,
            I => \N__14954\
        );

    \I__2085\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14954\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__14962\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__14959\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__14954\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__2081\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14944\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__14944\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__14941\,
            I => \N__14934\
        );

    \I__2078\ : InMux
    port map (
            O => \N__14940\,
            I => \N__14931\
        );

    \I__2077\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14928\
        );

    \I__2076\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14923\
        );

    \I__2075\ : InMux
    port map (
            O => \N__14937\,
            I => \N__14923\
        );

    \I__2074\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14920\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__14931\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__14928\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__14923\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__14920\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__2069\ : InMux
    port map (
            O => \N__14911\,
            I => \N__14904\
        );

    \I__2068\ : InMux
    port map (
            O => \N__14910\,
            I => \N__14904\
        );

    \I__2067\ : InMux
    port map (
            O => \N__14909\,
            I => \N__14901\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__14904\,
            I => \N__14898\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__14901\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__14898\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__14893\,
            I => \N__14887\
        );

    \I__2062\ : InMux
    port map (
            O => \N__14892\,
            I => \N__14883\
        );

    \I__2061\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14880\
        );

    \I__2060\ : InMux
    port map (
            O => \N__14890\,
            I => \N__14877\
        );

    \I__2059\ : InMux
    port map (
            O => \N__14887\,
            I => \N__14872\
        );

    \I__2058\ : InMux
    port map (
            O => \N__14886\,
            I => \N__14872\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__14883\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__14880\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__14877\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__14872\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__2053\ : InMux
    port map (
            O => \N__14863\,
            I => \N__14860\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__14860\,
            I => \this_vga_signals.SUM_2_i_1_0_3\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__14857\,
            I => \N__14854\
        );

    \I__2050\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14851\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__14851\,
            I => \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5Z0Z_0\
        );

    \I__2048\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14845\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__14845\,
            I => \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJHZ0Z5\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__14842\,
            I => \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i_cascade_\
        );

    \I__2045\ : InMux
    port map (
            O => \N__14839\,
            I => \N__14836\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__14836\,
            I => \N__14830\
        );

    \I__2043\ : InMux
    port map (
            O => \N__14835\,
            I => \N__14825\
        );

    \I__2042\ : InMux
    port map (
            O => \N__14834\,
            I => \N__14825\
        );

    \I__2041\ : InMux
    port map (
            O => \N__14833\,
            I => \N__14822\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__14830\,
            I => \N__14817\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__14825\,
            I => \N__14817\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__14822\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__14817\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2036\ : InMux
    port map (
            O => \N__14812\,
            I => \N__14809\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__14809\,
            I => \N__14806\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__14806\,
            I => \N__14801\
        );

    \I__2033\ : InMux
    port map (
            O => \N__14805\,
            I => \N__14798\
        );

    \I__2032\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14795\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__14801\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__14798\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__14795\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__2028\ : InMux
    port map (
            O => \N__14788\,
            I => \N__14782\
        );

    \I__2027\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14782\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__14782\,
            I => \N__14779\
        );

    \I__2025\ : Span4Mux_h
    port map (
            O => \N__14779\,
            I => \N__14775\
        );

    \I__2024\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14772\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__14775\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__14772\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__14767\,
            I => \N__14764\
        );

    \I__2020\ : InMux
    port map (
            O => \N__14764\,
            I => \N__14761\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__14761\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__14758\,
            I => \N__14755\
        );

    \I__2017\ : InMux
    port map (
            O => \N__14755\,
            I => \N__14752\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__14752\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1\
        );

    \I__2015\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14746\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__14746\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__14743\,
            I => \this_vga_signals.N_1_4_1_cascade_\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__14740\,
            I => \N_2_0_cascade_\
        );

    \I__2011\ : InMux
    port map (
            O => \N__14737\,
            I => \N__14732\
        );

    \I__2010\ : InMux
    port map (
            O => \N__14736\,
            I => \N__14729\
        );

    \I__2009\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14726\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__14732\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__14729\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__14726\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__14719\,
            I => \N__14711\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__14718\,
            I => \N__14707\
        );

    \I__2003\ : CEMux
    port map (
            O => \N__14717\,
            I => \N__14703\
        );

    \I__2002\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14700\
        );

    \I__2001\ : InMux
    port map (
            O => \N__14715\,
            I => \N__14695\
        );

    \I__2000\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14695\
        );

    \I__1999\ : InMux
    port map (
            O => \N__14711\,
            I => \N__14684\
        );

    \I__1998\ : InMux
    port map (
            O => \N__14710\,
            I => \N__14684\
        );

    \I__1997\ : InMux
    port map (
            O => \N__14707\,
            I => \N__14679\
        );

    \I__1996\ : InMux
    port map (
            O => \N__14706\,
            I => \N__14679\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__14703\,
            I => \N__14676\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__14700\,
            I => \N__14673\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__14695\,
            I => \N__14670\
        );

    \I__1992\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14665\
        );

    \I__1991\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14665\
        );

    \I__1990\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14659\
        );

    \I__1989\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14659\
        );

    \I__1988\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14654\
        );

    \I__1987\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14654\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14651\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__14679\,
            I => \N__14645\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__14676\,
            I => \N__14645\
        );

    \I__1983\ : Span4Mux_h
    port map (
            O => \N__14673\,
            I => \N__14642\
        );

    \I__1982\ : Sp12to4
    port map (
            O => \N__14670\,
            I => \N__14637\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__14665\,
            I => \N__14637\
        );

    \I__1980\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14633\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__14659\,
            I => \N__14626\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__14654\,
            I => \N__14626\
        );

    \I__1977\ : Span4Mux_h
    port map (
            O => \N__14651\,
            I => \N__14626\
        );

    \I__1976\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14623\
        );

    \I__1975\ : Span4Mux_h
    port map (
            O => \N__14645\,
            I => \N__14620\
        );

    \I__1974\ : Span4Mux_h
    port map (
            O => \N__14642\,
            I => \N__14617\
        );

    \I__1973\ : Span12Mux_h
    port map (
            O => \N__14637\,
            I => \N__14614\
        );

    \I__1972\ : InMux
    port map (
            O => \N__14636\,
            I => \N__14611\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__14633\,
            I => \N__14604\
        );

    \I__1970\ : Span4Mux_h
    port map (
            O => \N__14626\,
            I => \N__14604\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__14623\,
            I => \N__14604\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__14620\,
            I => \M_counter_q_RNILQS8_1\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__14617\,
            I => \M_counter_q_RNILQS8_1\
        );

    \I__1966\ : Odrv12
    port map (
            O => \N__14614\,
            I => \M_counter_q_RNILQS8_1\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__14611\,
            I => \M_counter_q_RNILQS8_1\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__14604\,
            I => \M_counter_q_RNILQS8_1\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__14593\,
            I => \this_vga_signals.M_pcounter_q_3_1_cascade_\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__14590\,
            I => \N__14586\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__14589\,
            I => \N__14582\
        );

    \I__1960\ : InMux
    port map (
            O => \N__14586\,
            I => \N__14579\
        );

    \I__1959\ : InMux
    port map (
            O => \N__14585\,
            I => \N__14574\
        );

    \I__1958\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14574\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__14579\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__14574\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__14569\,
            I => \N_3_0_cascade_\
        );

    \I__1954\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14558\
        );

    \I__1953\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14558\
        );

    \I__1952\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14553\
        );

    \I__1951\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14553\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__14558\,
            I => \this_vga_signals.M_pcounter_q_i_5_1\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__14553\,
            I => \this_vga_signals.M_pcounter_q_i_5_1\
        );

    \I__1948\ : InMux
    port map (
            O => \N__14548\,
            I => \N__14544\
        );

    \I__1947\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14541\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__14544\,
            I => \this_vga_signals.M_pcounter_q_i_5_0\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__14541\,
            I => \this_vga_signals.M_pcounter_q_i_5_0\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__14536\,
            I => \N__14532\
        );

    \I__1943\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14525\
        );

    \I__1942\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14522\
        );

    \I__1941\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14519\
        );

    \I__1940\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14512\
        );

    \I__1939\ : InMux
    port map (
            O => \N__14529\,
            I => \N__14512\
        );

    \I__1938\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14512\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__14525\,
            I => \N__14509\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__14522\,
            I => \N__14506\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__14519\,
            I => \N__14501\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__14512\,
            I => \N__14498\
        );

    \I__1933\ : Span4Mux_h
    port map (
            O => \N__14509\,
            I => \N__14493\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__14506\,
            I => \N__14493\
        );

    \I__1931\ : InMux
    port map (
            O => \N__14505\,
            I => \N__14488\
        );

    \I__1930\ : InMux
    port map (
            O => \N__14504\,
            I => \N__14488\
        );

    \I__1929\ : Span4Mux_h
    port map (
            O => \N__14501\,
            I => \N__14485\
        );

    \I__1928\ : Span4Mux_h
    port map (
            O => \N__14498\,
            I => \N__14482\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__14493\,
            I => \N__14479\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14476\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__14485\,
            I => \N__14472\
        );

    \I__1924\ : Span4Mux_h
    port map (
            O => \N__14482\,
            I => \N__14469\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__14479\,
            I => \N__14464\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__14476\,
            I => \N__14464\
        );

    \I__1921\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14461\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__14472\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__14469\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__14464\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__14461\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__1916\ : InMux
    port map (
            O => \N__14452\,
            I => \N__14449\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__14449\,
            I => \this_vga_signals.M_pcounter_q_3_0\
        );

    \I__1914\ : CEMux
    port map (
            O => \N__14446\,
            I => \N__14442\
        );

    \I__1913\ : CEMux
    port map (
            O => \N__14445\,
            I => \N__14439\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__14442\,
            I => \N__14436\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__14439\,
            I => \N__14433\
        );

    \I__1910\ : Span4Mux_v
    port map (
            O => \N__14436\,
            I => \N__14430\
        );

    \I__1909\ : Span4Mux_h
    port map (
            O => \N__14433\,
            I => \N__14427\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__14430\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__14427\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__1906\ : InMux
    port map (
            O => \N__14422\,
            I => \N__14419\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__14419\,
            I => \N__14416\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__14416\,
            I => \N__14412\
        );

    \I__1903\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14409\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__14412\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__14409\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1900\ : InMux
    port map (
            O => \N__14404\,
            I => \N__14401\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__14401\,
            I => \N__14397\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__14400\,
            I => \N__14393\
        );

    \I__1897\ : Span4Mux_h
    port map (
            O => \N__14397\,
            I => \N__14389\
        );

    \I__1896\ : InMux
    port map (
            O => \N__14396\,
            I => \N__14386\
        );

    \I__1895\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14381\
        );

    \I__1894\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14381\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__14389\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__14386\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__14381\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1890\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14371\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__14371\,
            I => \N__14368\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__14368\,
            I => \N__14363\
        );

    \I__1887\ : InMux
    port map (
            O => \N__14367\,
            I => \N__14358\
        );

    \I__1886\ : InMux
    port map (
            O => \N__14366\,
            I => \N__14358\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__14363\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_2\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__14358\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_2\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__14353\,
            I => \N__14350\
        );

    \I__1882\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14347\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__14347\,
            I => \N__14344\
        );

    \I__1880\ : Span12Mux_h
    port map (
            O => \N__14344\,
            I => \N__14341\
        );

    \I__1879\ : Odrv12
    port map (
            O => \N__14341\,
            I => \M_this_vga_signals_address_3\
        );

    \I__1878\ : CEMux
    port map (
            O => \N__14338\,
            I => \N__14335\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__14335\,
            I => \N__14331\
        );

    \I__1876\ : CEMux
    port map (
            O => \N__14334\,
            I => \N__14328\
        );

    \I__1875\ : Span4Mux_h
    port map (
            O => \N__14331\,
            I => \N__14325\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__14328\,
            I => \N__14322\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__14325\,
            I => \N__14319\
        );

    \I__1872\ : Span4Mux_h
    port map (
            O => \N__14322\,
            I => \N__14316\
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__14319\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__14316\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__1869\ : InMux
    port map (
            O => \N__14311\,
            I => \N__14308\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__14308\,
            I => \N__14305\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__14305\,
            I => \N__14298\
        );

    \I__1866\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14295\
        );

    \I__1865\ : InMux
    port map (
            O => \N__14303\,
            I => \N__14290\
        );

    \I__1864\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14290\
        );

    \I__1863\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14287\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__14298\,
            I => \this_vga_signals.N_3_2_1\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__14295\,
            I => \this_vga_signals.N_3_2_1\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__14290\,
            I => \this_vga_signals.N_3_2_1\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__14287\,
            I => \this_vga_signals.N_3_2_1\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__14278\,
            I => \N__14275\
        );

    \I__1857\ : InMux
    port map (
            O => \N__14275\,
            I => \N__14272\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__14272\,
            I => \N__14269\
        );

    \I__1855\ : Span12Mux_h
    port map (
            O => \N__14269\,
            I => \N__14266\
        );

    \I__1854\ : Odrv12
    port map (
            O => \N__14266\,
            I => \M_this_vga_signals_address_6\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__14263\,
            I => \N__14260\
        );

    \I__1852\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14256\
        );

    \I__1851\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14253\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__14256\,
            I => \N__14250\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__14253\,
            I => \N__14247\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__14250\,
            I => \N__14242\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__14247\,
            I => \N__14242\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__14242\,
            I => \this_vga_signals.M_vcounter_d7lto8_1\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__14239\,
            I => \N__14236\
        );

    \I__1844\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14233\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__14233\,
            I => \this_vga_signals.M_lcounter_d_0_sqmuxa\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__14230\,
            I => \this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_\
        );

    \I__1841\ : InMux
    port map (
            O => \N__14227\,
            I => \N__14224\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__14224\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_1_0\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__14221\,
            I => \this_vga_signals.g1_0_0_1_cascade_\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__14218\,
            I => \this_vga_signals.g2_0_1_cascade_\
        );

    \I__1837\ : InMux
    port map (
            O => \N__14215\,
            I => \N__14212\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__14212\,
            I => \this_vga_signals.vaddress_6_6\
        );

    \I__1835\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14206\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__14206\,
            I => \this_vga_signals.N_4_1_0\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__14203\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_\
        );

    \I__1832\ : InMux
    port map (
            O => \N__14200\,
            I => \N__14197\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__14197\,
            I => \this_vga_signals.g0_i_x4_0_0\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__14194\,
            I => \this_vga_signals.g1_4_cascade_\
        );

    \I__1829\ : InMux
    port map (
            O => \N__14191\,
            I => \N__14188\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__14188\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_1_0_0_1\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__14185\,
            I => \this_vga_signals.g0_2_0_0_1_cascade_\
        );

    \I__1826\ : InMux
    port map (
            O => \N__14182\,
            I => \N__14179\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__14179\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_0_0_0\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__14176\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\
        );

    \I__1823\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14170\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__14170\,
            I => \N__14167\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__14167\,
            I => \this_vga_signals.g1_0_1\
        );

    \I__1820\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14161\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__14161\,
            I => \this_vga_signals.g0_31_N_5L8\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__14158\,
            I => \N__14155\
        );

    \I__1817\ : InMux
    port map (
            O => \N__14155\,
            I => \N__14152\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__14152\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_0\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__14149\,
            I => \this_vga_signals.m9_1_cascade_\
        );

    \I__1814\ : InMux
    port map (
            O => \N__14146\,
            I => \N__14143\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__14143\,
            I => \this_vga_signals.g2_1_0\
        );

    \I__1812\ : InMux
    port map (
            O => \N__14140\,
            I => \N__14137\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__14137\,
            I => \N__14133\
        );

    \I__1810\ : InMux
    port map (
            O => \N__14136\,
            I => \N__14130\
        );

    \I__1809\ : Span4Mux_h
    port map (
            O => \N__14133\,
            I => \N__14125\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__14130\,
            I => \N__14125\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__14125\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__14122\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_\
        );

    \I__1805\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14116\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__14116\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__1803\ : InMux
    port map (
            O => \N__14113\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__1802\ : InMux
    port map (
            O => \N__14110\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__1801\ : InMux
    port map (
            O => \N__14107\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__1800\ : InMux
    port map (
            O => \N__14104\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__1799\ : InMux
    port map (
            O => \N__14101\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__1798\ : InMux
    port map (
            O => \N__14098\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__1797\ : InMux
    port map (
            O => \N__14095\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__1796\ : InMux
    port map (
            O => \N__14092\,
            I => \bfn_10_12_0_\
        );

    \I__1795\ : InMux
    port map (
            O => \N__14089\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__1794\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14083\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__14083\,
            I => \N__14080\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__14080\,
            I => \this_sprites_ram.mem_out_bus4_3\
        );

    \I__1791\ : InMux
    port map (
            O => \N__14077\,
            I => \N__14074\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__14074\,
            I => \N__14071\
        );

    \I__1789\ : Span4Mux_v
    port map (
            O => \N__14071\,
            I => \N__14068\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__14068\,
            I => \N__14065\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__14065\,
            I => \N__14062\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__14062\,
            I => \this_sprites_ram.mem_out_bus0_3\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__14059\,
            I => \N__14056\
        );

    \I__1784\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14053\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__14053\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\
        );

    \I__1782\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14047\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__14047\,
            I => \N__14044\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__14044\,
            I => \N__14041\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__14041\,
            I => \this_sprites_ram.mem_out_bus5_3\
        );

    \I__1778\ : InMux
    port map (
            O => \N__14038\,
            I => \N__14035\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__14035\,
            I => \N__14032\
        );

    \I__1776\ : Span4Mux_v
    port map (
            O => \N__14032\,
            I => \N__14029\
        );

    \I__1775\ : Span4Mux_v
    port map (
            O => \N__14029\,
            I => \N__14026\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__14026\,
            I => \this_sprites_ram.mem_out_bus1_3\
        );

    \I__1773\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14020\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__14020\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\
        );

    \I__1771\ : InMux
    port map (
            O => \N__14017\,
            I => \N__14014\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__14014\,
            I => \N__14007\
        );

    \I__1769\ : InMux
    port map (
            O => \N__14013\,
            I => \N__14004\
        );

    \I__1768\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14001\
        );

    \I__1767\ : InMux
    port map (
            O => \N__14011\,
            I => \N__13998\
        );

    \I__1766\ : InMux
    port map (
            O => \N__14010\,
            I => \N__13995\
        );

    \I__1765\ : Span4Mux_h
    port map (
            O => \N__14007\,
            I => \N__13990\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__14004\,
            I => \N__13985\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__14001\,
            I => \N__13985\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__13998\,
            I => \N__13980\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__13995\,
            I => \N__13980\
        );

    \I__1760\ : InMux
    port map (
            O => \N__13994\,
            I => \N__13977\
        );

    \I__1759\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13974\
        );

    \I__1758\ : Odrv4
    port map (
            O => \N__13990\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__13985\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__13980\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__13977\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__13974\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__13963\,
            I => \N__13960\
        );

    \I__1752\ : InMux
    port map (
            O => \N__13960\,
            I => \N__13957\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__13957\,
            I => \N__13954\
        );

    \I__1750\ : Span12Mux_h
    port map (
            O => \N__13954\,
            I => \N__13951\
        );

    \I__1749\ : Odrv12
    port map (
            O => \N__13951\,
            I => \M_this_vga_signals_address_4\
        );

    \I__1748\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13945\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__13945\,
            I => \N__13942\
        );

    \I__1746\ : Span4Mux_v
    port map (
            O => \N__13942\,
            I => \N__13939\
        );

    \I__1745\ : Span4Mux_v
    port map (
            O => \N__13939\,
            I => \N__13936\
        );

    \I__1744\ : Span4Mux_v
    port map (
            O => \N__13936\,
            I => \N__13933\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__13933\,
            I => \this_sprites_ram.mem_out_bus7_0\
        );

    \I__1742\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13927\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__13927\,
            I => \N__13924\
        );

    \I__1740\ : Span4Mux_h
    port map (
            O => \N__13924\,
            I => \N__13921\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__13921\,
            I => \this_sprites_ram.mem_out_bus3_0\
        );

    \I__1738\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13915\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__13915\,
            I => \N__13910\
        );

    \I__1736\ : InMux
    port map (
            O => \N__13914\,
            I => \N__13905\
        );

    \I__1735\ : InMux
    port map (
            O => \N__13913\,
            I => \N__13905\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__13910\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__13905\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__13900\,
            I => \N__13897\
        );

    \I__1731\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13894\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__13894\,
            I => \N__13891\
        );

    \I__1729\ : Span12Mux_h
    port map (
            O => \N__13891\,
            I => \N__13888\
        );

    \I__1728\ : Odrv12
    port map (
            O => \N__13888\,
            I => \M_this_vga_signals_address_2\
        );

    \I__1727\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13882\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__13882\,
            I => \N__13879\
        );

    \I__1725\ : Span4Mux_h
    port map (
            O => \N__13879\,
            I => \N__13876\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__13876\,
            I => \this_vga_ramdac.m19\
        );

    \I__1723\ : InMux
    port map (
            O => \N__13873\,
            I => \N__13870\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__13870\,
            I => \N__13867\
        );

    \I__1721\ : Span4Mux_v
    port map (
            O => \N__13867\,
            I => \N__13863\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__13866\,
            I => \N__13860\
        );

    \I__1719\ : Span4Mux_h
    port map (
            O => \N__13863\,
            I => \N__13857\
        );

    \I__1718\ : InMux
    port map (
            O => \N__13860\,
            I => \N__13854\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__13857\,
            I => \this_vga_ramdac.N_2874_reto\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__13854\,
            I => \this_vga_ramdac.N_2874_reto\
        );

    \I__1715\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13841\
        );

    \I__1714\ : InMux
    port map (
            O => \N__13848\,
            I => \N__13841\
        );

    \I__1713\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13838\
        );

    \I__1712\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13835\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__13841\,
            I => \N__13831\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__13838\,
            I => \N__13826\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__13835\,
            I => \N__13826\
        );

    \I__1708\ : InMux
    port map (
            O => \N__13834\,
            I => \N__13822\
        );

    \I__1707\ : Span4Mux_v
    port map (
            O => \N__13831\,
            I => \N__13817\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__13826\,
            I => \N__13817\
        );

    \I__1705\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13814\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__13822\,
            I => \N__13806\
        );

    \I__1703\ : Sp12to4
    port map (
            O => \N__13817\,
            I => \N__13806\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__13814\,
            I => \N__13806\
        );

    \I__1701\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13803\
        );

    \I__1700\ : Odrv12
    port map (
            O => \N__13806\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__13803\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__1698\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13795\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__13795\,
            I => \N__13792\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__13792\,
            I => \N__13789\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__13789\,
            I => \N__13786\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__13786\,
            I => \N__13783\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__13783\,
            I => \this_sprites_ram.mem_out_bus7_3\
        );

    \I__1692\ : InMux
    port map (
            O => \N__13780\,
            I => \N__13777\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__13777\,
            I => \N__13774\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__13774\,
            I => \this_sprites_ram.mem_out_bus3_3\
        );

    \I__1689\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13768\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__13768\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\
        );

    \I__1687\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13762\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__13762\,
            I => \N__13758\
        );

    \I__1685\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13755\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__13758\,
            I => \this_vga_signals.vaddress_6_5\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__13755\,
            I => \this_vga_signals.vaddress_6_5\
        );

    \I__1682\ : InMux
    port map (
            O => \N__13750\,
            I => \N__13747\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__13747\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_1_0_0\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__13744\,
            I => \N__13740\
        );

    \I__1679\ : InMux
    port map (
            O => \N__13743\,
            I => \N__13735\
        );

    \I__1678\ : InMux
    port map (
            O => \N__13740\,
            I => \N__13735\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__13735\,
            I => \N__13732\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__13732\,
            I => \this_vga_signals.vaddress_3_0_6\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__13729\,
            I => \this_vga_signals.vaddress_3_5_cascade_\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__13726\,
            I => \this_vga_signals.vaddress_3_6_cascade_\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__13723\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\
        );

    \I__1672\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13717\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__13717\,
            I => \N__13714\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__13714\,
            I => \N__13711\
        );

    \I__1669\ : Sp12to4
    port map (
            O => \N__13711\,
            I => \N__13708\
        );

    \I__1668\ : Span12Mux_h
    port map (
            O => \N__13708\,
            I => \N__13705\
        );

    \I__1667\ : Odrv12
    port map (
            O => \N__13705\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__1666\ : InMux
    port map (
            O => \N__13702\,
            I => \N__13699\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__13699\,
            I => \N__13696\
        );

    \I__1664\ : Span4Mux_v
    port map (
            O => \N__13696\,
            I => \N__13693\
        );

    \I__1663\ : Span4Mux_v
    port map (
            O => \N__13693\,
            I => \N__13690\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__13690\,
            I => \this_sprites_ram.mem_out_bus6_3\
        );

    \I__1661\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13684\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__13684\,
            I => \N__13681\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__13681\,
            I => \N__13678\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__13678\,
            I => \this_sprites_ram.mem_out_bus2_3\
        );

    \I__1657\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13672\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__13672\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__13669\,
            I => \this_vga_signals.vaddress_3_0_6_cascade_\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__13666\,
            I => \this_vga_signals.g2_3_cascade_\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__13663\,
            I => \this_vga_signals.g1_1_1_cascade_\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__13660\,
            I => \this_vga_signals.g0_i_x4_0_2_cascade_\
        );

    \I__1651\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13654\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__13654\,
            I => \this_vga_signals.g0_31_N_4L6\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__13651\,
            I => \this_vga_signals.if_m8_0_a3_1_1_4_cascade_\
        );

    \I__1648\ : InMux
    port map (
            O => \N__13648\,
            I => \N__13645\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__13645\,
            I => \this_vga_signals.g0_31_N_3L3\
        );

    \I__1646\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13639\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__13639\,
            I => \this_vga_signals.g3_3_0\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__13636\,
            I => \this_vga_signals.if_m8_0_a3_1_1_2_cascade_\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__13633\,
            I => \this_vga_signals.g0_8_0_cascade_\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__13630\,
            I => \this_vga_signals.vaddress_2_5_cascade_\
        );

    \I__1641\ : InMux
    port map (
            O => \N__13627\,
            I => \N__13622\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__13626\,
            I => \N__13619\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__13625\,
            I => \N__13615\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__13622\,
            I => \N__13609\
        );

    \I__1637\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13605\
        );

    \I__1636\ : InMux
    port map (
            O => \N__13618\,
            I => \N__13600\
        );

    \I__1635\ : InMux
    port map (
            O => \N__13615\,
            I => \N__13600\
        );

    \I__1634\ : InMux
    port map (
            O => \N__13614\,
            I => \N__13595\
        );

    \I__1633\ : InMux
    port map (
            O => \N__13613\,
            I => \N__13595\
        );

    \I__1632\ : InMux
    port map (
            O => \N__13612\,
            I => \N__13592\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__13609\,
            I => \N__13589\
        );

    \I__1630\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13586\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__13605\,
            I => \N__13581\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__13600\,
            I => \N__13581\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__13595\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__13592\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__13589\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__13586\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__13581\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1622\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13567\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__13567\,
            I => \N__13564\
        );

    \I__1620\ : Span4Mux_h
    port map (
            O => \N__13564\,
            I => \N__13560\
        );

    \I__1619\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13557\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__13560\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__13557\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0\
        );

    \I__1616\ : InMux
    port map (
            O => \N__13552\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__1615\ : InMux
    port map (
            O => \N__13549\,
            I => \bfn_7_20_0_\
        );

    \I__1614\ : InMux
    port map (
            O => \N__13546\,
            I => \N__13542\
        );

    \I__1613\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13539\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__13542\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__13539\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0\
        );

    \I__1610\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13529\
        );

    \I__1609\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13526\
        );

    \I__1608\ : InMux
    port map (
            O => \N__13532\,
            I => \N__13522\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__13529\,
            I => \N__13519\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__13526\,
            I => \N__13516\
        );

    \I__1605\ : InMux
    port map (
            O => \N__13525\,
            I => \N__13513\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__13522\,
            I => \N__13510\
        );

    \I__1603\ : Span4Mux_v
    port map (
            O => \N__13519\,
            I => \N__13503\
        );

    \I__1602\ : Span4Mux_h
    port map (
            O => \N__13516\,
            I => \N__13496\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__13513\,
            I => \N__13496\
        );

    \I__1600\ : Span4Mux_v
    port map (
            O => \N__13510\,
            I => \N__13496\
        );

    \I__1599\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13493\
        );

    \I__1598\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13486\
        );

    \I__1597\ : InMux
    port map (
            O => \N__13507\,
            I => \N__13486\
        );

    \I__1596\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13486\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__13503\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__13496\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__13493\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__13486\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1591\ : CEMux
    port map (
            O => \N__13477\,
            I => \N__13473\
        );

    \I__1590\ : CEMux
    port map (
            O => \N__13476\,
            I => \N__13469\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__13473\,
            I => \N__13466\
        );

    \I__1588\ : CEMux
    port map (
            O => \N__13472\,
            I => \N__13463\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__13469\,
            I => \N__13460\
        );

    \I__1586\ : Span4Mux_h
    port map (
            O => \N__13466\,
            I => \N__13455\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__13463\,
            I => \N__13455\
        );

    \I__1584\ : Span4Mux_v
    port map (
            O => \N__13460\,
            I => \N__13452\
        );

    \I__1583\ : Span4Mux_h
    port map (
            O => \N__13455\,
            I => \N__13449\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__13452\,
            I => \this_vga_signals.N_614_0\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__13449\,
            I => \this_vga_signals.N_614_0\
        );

    \I__1580\ : SRMux
    port map (
            O => \N__13444\,
            I => \N__13440\
        );

    \I__1579\ : SRMux
    port map (
            O => \N__13443\,
            I => \N__13437\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__13440\,
            I => \N__13433\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__13437\,
            I => \N__13428\
        );

    \I__1576\ : SRMux
    port map (
            O => \N__13436\,
            I => \N__13425\
        );

    \I__1575\ : Span4Mux_v
    port map (
            O => \N__13433\,
            I => \N__13422\
        );

    \I__1574\ : SRMux
    port map (
            O => \N__13432\,
            I => \N__13419\
        );

    \I__1573\ : SRMux
    port map (
            O => \N__13431\,
            I => \N__13416\
        );

    \I__1572\ : Span4Mux_h
    port map (
            O => \N__13428\,
            I => \N__13412\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__13425\,
            I => \N__13409\
        );

    \I__1570\ : Span4Mux_h
    port map (
            O => \N__13422\,
            I => \N__13404\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__13419\,
            I => \N__13404\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__13416\,
            I => \N__13401\
        );

    \I__1567\ : InMux
    port map (
            O => \N__13415\,
            I => \N__13398\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__13412\,
            I => \this_vga_signals.N_931_1\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__13409\,
            I => \this_vga_signals.N_931_1\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__13404\,
            I => \this_vga_signals.N_931_1\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__13401\,
            I => \this_vga_signals.N_931_1\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__13398\,
            I => \this_vga_signals.N_931_1\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__13387\,
            I => \this_vga_signals.vaddress_0_5_cascade_\
        );

    \I__1560\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13381\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__13381\,
            I => \N__13375\
        );

    \I__1558\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13370\
        );

    \I__1557\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13370\
        );

    \I__1556\ : InMux
    port map (
            O => \N__13378\,
            I => \N__13367\
        );

    \I__1555\ : Odrv12
    port map (
            O => \N__13375\,
            I => \this_vga_signals.mult1_un75_sum_axb2\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__13370\,
            I => \this_vga_signals.mult1_un75_sum_axb2\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__13367\,
            I => \this_vga_signals.mult1_un75_sum_axb2\
        );

    \I__1552\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13356\
        );

    \I__1551\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13353\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__13356\,
            I => \this_vga_signals.mult1_un75_sum_axb1\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__13353\,
            I => \this_vga_signals.mult1_un75_sum_axb1\
        );

    \I__1548\ : InMux
    port map (
            O => \N__13348\,
            I => \N__13345\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__13345\,
            I => \N__13342\
        );

    \I__1546\ : Span4Mux_h
    port map (
            O => \N__13342\,
            I => \N__13338\
        );

    \I__1545\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13335\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__13338\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_d\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__13335\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_d\
        );

    \I__1542\ : InMux
    port map (
            O => \N__13330\,
            I => \N__13325\
        );

    \I__1541\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13320\
        );

    \I__1540\ : InMux
    port map (
            O => \N__13328\,
            I => \N__13320\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__13325\,
            I => \N__13311\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__13320\,
            I => \N__13307\
        );

    \I__1537\ : InMux
    port map (
            O => \N__13319\,
            I => \N__13304\
        );

    \I__1536\ : InMux
    port map (
            O => \N__13318\,
            I => \N__13299\
        );

    \I__1535\ : InMux
    port map (
            O => \N__13317\,
            I => \N__13299\
        );

    \I__1534\ : InMux
    port map (
            O => \N__13316\,
            I => \N__13292\
        );

    \I__1533\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13292\
        );

    \I__1532\ : InMux
    port map (
            O => \N__13314\,
            I => \N__13292\
        );

    \I__1531\ : Span4Mux_h
    port map (
            O => \N__13311\,
            I => \N__13289\
        );

    \I__1530\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13286\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__13307\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__13304\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__13299\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__13292\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__13289\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__13286\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__13273\,
            I => \N__13270\
        );

    \I__1522\ : InMux
    port map (
            O => \N__13270\,
            I => \N__13266\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__13269\,
            I => \N__13260\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__13266\,
            I => \N__13256\
        );

    \I__1519\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13251\
        );

    \I__1518\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13251\
        );

    \I__1517\ : InMux
    port map (
            O => \N__13263\,
            I => \N__13248\
        );

    \I__1516\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13243\
        );

    \I__1515\ : InMux
    port map (
            O => \N__13259\,
            I => \N__13243\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__13256\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__13251\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__13248\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__13243\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1510\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__13231\,
            I => \N__13228\
        );

    \I__1508\ : Odrv12
    port map (
            O => \N__13228\,
            I => \this_vga_signals.M_hcounter_d7lt4\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__13225\,
            I => \N__13219\
        );

    \I__1506\ : InMux
    port map (
            O => \N__13224\,
            I => \N__13214\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__13223\,
            I => \N__13210\
        );

    \I__1504\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13204\
        );

    \I__1503\ : InMux
    port map (
            O => \N__13219\,
            I => \N__13201\
        );

    \I__1502\ : InMux
    port map (
            O => \N__13218\,
            I => \N__13196\
        );

    \I__1501\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13196\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__13214\,
            I => \N__13191\
        );

    \I__1499\ : InMux
    port map (
            O => \N__13213\,
            I => \N__13188\
        );

    \I__1498\ : InMux
    port map (
            O => \N__13210\,
            I => \N__13181\
        );

    \I__1497\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13181\
        );

    \I__1496\ : InMux
    port map (
            O => \N__13208\,
            I => \N__13181\
        );

    \I__1495\ : InMux
    port map (
            O => \N__13207\,
            I => \N__13178\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__13204\,
            I => \N__13170\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__13201\,
            I => \N__13170\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__13196\,
            I => \N__13170\
        );

    \I__1491\ : InMux
    port map (
            O => \N__13195\,
            I => \N__13167\
        );

    \I__1490\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13164\
        );

    \I__1489\ : Span4Mux_h
    port map (
            O => \N__13191\,
            I => \N__13161\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__13188\,
            I => \N__13154\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__13181\,
            I => \N__13154\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__13178\,
            I => \N__13154\
        );

    \I__1485\ : InMux
    port map (
            O => \N__13177\,
            I => \N__13151\
        );

    \I__1484\ : Span4Mux_v
    port map (
            O => \N__13170\,
            I => \N__13146\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__13167\,
            I => \N__13146\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__13164\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__13161\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__13154\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__13151\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__13146\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1477\ : InMux
    port map (
            O => \N__13135\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__13132\,
            I => \N__13123\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__13131\,
            I => \N__13120\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__13130\,
            I => \N__13115\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__13129\,
            I => \N__13112\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__13128\,
            I => \N__13107\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__13127\,
            I => \N__13101\
        );

    \I__1470\ : InMux
    port map (
            O => \N__13126\,
            I => \N__13094\
        );

    \I__1469\ : InMux
    port map (
            O => \N__13123\,
            I => \N__13094\
        );

    \I__1468\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13094\
        );

    \I__1467\ : InMux
    port map (
            O => \N__13119\,
            I => \N__13087\
        );

    \I__1466\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13087\
        );

    \I__1465\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13087\
        );

    \I__1464\ : InMux
    port map (
            O => \N__13112\,
            I => \N__13084\
        );

    \I__1463\ : InMux
    port map (
            O => \N__13111\,
            I => \N__13081\
        );

    \I__1462\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13078\
        );

    \I__1461\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13075\
        );

    \I__1460\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13068\
        );

    \I__1459\ : InMux
    port map (
            O => \N__13105\,
            I => \N__13068\
        );

    \I__1458\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13068\
        );

    \I__1457\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13063\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__13094\,
            I => \N__13052\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__13087\,
            I => \N__13052\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__13084\,
            I => \N__13052\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__13081\,
            I => \N__13052\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__13078\,
            I => \N__13052\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__13075\,
            I => \N__13049\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__13068\,
            I => \N__13046\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__13067\,
            I => \N__13043\
        );

    \I__1448\ : InMux
    port map (
            O => \N__13066\,
            I => \N__13039\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__13063\,
            I => \N__13036\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__13052\,
            I => \N__13031\
        );

    \I__1445\ : Span4Mux_h
    port map (
            O => \N__13049\,
            I => \N__13031\
        );

    \I__1444\ : Span4Mux_h
    port map (
            O => \N__13046\,
            I => \N__13028\
        );

    \I__1443\ : InMux
    port map (
            O => \N__13043\,
            I => \N__13023\
        );

    \I__1442\ : InMux
    port map (
            O => \N__13042\,
            I => \N__13023\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__13039\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__13036\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1439\ : Odrv4
    port map (
            O => \N__13031\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__13028\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__13023\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1436\ : InMux
    port map (
            O => \N__13012\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__13009\,
            I => \N__13006\
        );

    \I__1434\ : InMux
    port map (
            O => \N__13006\,
            I => \N__12992\
        );

    \I__1433\ : InMux
    port map (
            O => \N__13005\,
            I => \N__12992\
        );

    \I__1432\ : InMux
    port map (
            O => \N__13004\,
            I => \N__12989\
        );

    \I__1431\ : InMux
    port map (
            O => \N__13003\,
            I => \N__12986\
        );

    \I__1430\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12981\
        );

    \I__1429\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12981\
        );

    \I__1428\ : InMux
    port map (
            O => \N__13000\,
            I => \N__12978\
        );

    \I__1427\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12973\
        );

    \I__1426\ : InMux
    port map (
            O => \N__12998\,
            I => \N__12973\
        );

    \I__1425\ : InMux
    port map (
            O => \N__12997\,
            I => \N__12967\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__12992\,
            I => \N__12962\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__12989\,
            I => \N__12962\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__12986\,
            I => \N__12953\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__12981\,
            I => \N__12953\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__12978\,
            I => \N__12953\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__12973\,
            I => \N__12953\
        );

    \I__1418\ : InMux
    port map (
            O => \N__12972\,
            I => \N__12943\
        );

    \I__1417\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12943\
        );

    \I__1416\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12943\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__12967\,
            I => \N__12936\
        );

    \I__1414\ : Span4Mux_h
    port map (
            O => \N__12962\,
            I => \N__12936\
        );

    \I__1413\ : Span4Mux_v
    port map (
            O => \N__12953\,
            I => \N__12936\
        );

    \I__1412\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12933\
        );

    \I__1411\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12928\
        );

    \I__1410\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12928\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__12943\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__12936\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__12933\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__12928\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1405\ : InMux
    port map (
            O => \N__12919\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__1404\ : InMux
    port map (
            O => \N__12916\,
            I => \N__12907\
        );

    \I__1403\ : InMux
    port map (
            O => \N__12915\,
            I => \N__12907\
        );

    \I__1402\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12904\
        );

    \I__1401\ : InMux
    port map (
            O => \N__12913\,
            I => \N__12899\
        );

    \I__1400\ : InMux
    port map (
            O => \N__12912\,
            I => \N__12899\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__12907\,
            I => \N__12890\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__12904\,
            I => \N__12890\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__12899\,
            I => \N__12890\
        );

    \I__1396\ : InMux
    port map (
            O => \N__12898\,
            I => \N__12887\
        );

    \I__1395\ : InMux
    port map (
            O => \N__12897\,
            I => \N__12875\
        );

    \I__1394\ : Span4Mux_v
    port map (
            O => \N__12890\,
            I => \N__12870\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__12887\,
            I => \N__12870\
        );

    \I__1392\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12861\
        );

    \I__1391\ : InMux
    port map (
            O => \N__12885\,
            I => \N__12861\
        );

    \I__1390\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12861\
        );

    \I__1389\ : InMux
    port map (
            O => \N__12883\,
            I => \N__12861\
        );

    \I__1388\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12856\
        );

    \I__1387\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12856\
        );

    \I__1386\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12849\
        );

    \I__1385\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12849\
        );

    \I__1384\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12849\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__12875\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__12870\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__12861\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__12856\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__12849\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1378\ : InMux
    port map (
            O => \N__12838\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__1377\ : InMux
    port map (
            O => \N__12835\,
            I => \N__12827\
        );

    \I__1376\ : InMux
    port map (
            O => \N__12834\,
            I => \N__12827\
        );

    \I__1375\ : InMux
    port map (
            O => \N__12833\,
            I => \N__12818\
        );

    \I__1374\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12818\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__12827\,
            I => \N__12814\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__12826\,
            I => \N__12810\
        );

    \I__1371\ : InMux
    port map (
            O => \N__12825\,
            I => \N__12805\
        );

    \I__1370\ : InMux
    port map (
            O => \N__12824\,
            I => \N__12805\
        );

    \I__1369\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12802\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__12818\,
            I => \N__12799\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__12817\,
            I => \N__12794\
        );

    \I__1366\ : Span4Mux_v
    port map (
            O => \N__12814\,
            I => \N__12788\
        );

    \I__1365\ : InMux
    port map (
            O => \N__12813\,
            I => \N__12785\
        );

    \I__1364\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12782\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__12805\,
            I => \N__12779\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__12802\,
            I => \N__12774\
        );

    \I__1361\ : Span4Mux_h
    port map (
            O => \N__12799\,
            I => \N__12774\
        );

    \I__1360\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12771\
        );

    \I__1359\ : InMux
    port map (
            O => \N__12797\,
            I => \N__12766\
        );

    \I__1358\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12766\
        );

    \I__1357\ : InMux
    port map (
            O => \N__12793\,
            I => \N__12759\
        );

    \I__1356\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12759\
        );

    \I__1355\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12759\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__12788\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__12785\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__12782\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__12779\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__12774\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__12771\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__12766\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__12759\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1346\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12736\
        );

    \I__1345\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12736\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__12736\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0\
        );

    \I__1343\ : InMux
    port map (
            O => \N__12733\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__1342\ : InMux
    port map (
            O => \N__12730\,
            I => \N__12727\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__12727\,
            I => \N__12722\
        );

    \I__1340\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12714\
        );

    \I__1339\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12711\
        );

    \I__1338\ : Span4Mux_v
    port map (
            O => \N__12722\,
            I => \N__12708\
        );

    \I__1337\ : InMux
    port map (
            O => \N__12721\,
            I => \N__12705\
        );

    \I__1336\ : InMux
    port map (
            O => \N__12720\,
            I => \N__12696\
        );

    \I__1335\ : InMux
    port map (
            O => \N__12719\,
            I => \N__12696\
        );

    \I__1334\ : InMux
    port map (
            O => \N__12718\,
            I => \N__12696\
        );

    \I__1333\ : InMux
    port map (
            O => \N__12717\,
            I => \N__12696\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__12714\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__12711\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__12708\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__12705\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__12696\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1327\ : InMux
    port map (
            O => \N__12685\,
            I => \N__12682\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__12682\,
            I => \N__12679\
        );

    \I__1325\ : Span4Mux_h
    port map (
            O => \N__12679\,
            I => \N__12675\
        );

    \I__1324\ : InMux
    port map (
            O => \N__12678\,
            I => \N__12672\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__12675\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__12672\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0\
        );

    \I__1321\ : InMux
    port map (
            O => \N__12667\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__12664\,
            I => \this_vga_signals.if_m7_0_x4_0_cascade_\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__12661\,
            I => \this_vga_signals.if_N_9_1_cascade_\
        );

    \I__1318\ : InMux
    port map (
            O => \N__12658\,
            I => \N__12653\
        );

    \I__1317\ : InMux
    port map (
            O => \N__12657\,
            I => \N__12648\
        );

    \I__1316\ : InMux
    port map (
            O => \N__12656\,
            I => \N__12648\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__12653\,
            I => \this_vga_signals.mult1_un75_sum_c2_0\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__12648\,
            I => \this_vga_signals.mult1_un75_sum_c2_0\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__12643\,
            I => \N__12640\
        );

    \I__1312\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12637\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__12637\,
            I => \this_vga_signals.mult1_un82_sum_c3\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__12634\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_cascade_\
        );

    \I__1309\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12628\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__12628\,
            I => \this_vga_signals.mult1_un89_sum_c3\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__12625\,
            I => \N__12622\
        );

    \I__1306\ : InMux
    port map (
            O => \N__12622\,
            I => \N__12619\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__12619\,
            I => \N__12616\
        );

    \I__1304\ : Span12Mux_h
    port map (
            O => \N__12616\,
            I => \N__12613\
        );

    \I__1303\ : Odrv12
    port map (
            O => \N__12613\,
            I => \M_this_vga_signals_address_0\
        );

    \I__1302\ : InMux
    port map (
            O => \N__12610\,
            I => \N__12607\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__12607\,
            I => \this_vga_signals.d_N_12\
        );

    \I__1300\ : InMux
    port map (
            O => \N__12604\,
            I => \N__12601\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__12601\,
            I => \this_vga_signals.d_N_11\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__12598\,
            I => \N__12595\
        );

    \I__1297\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12592\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__12592\,
            I => \N__12589\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__12589\,
            I => \this_vga_signals.M_hcounter_q_RNIUAKU9Z0Z_4\
        );

    \I__1294\ : InMux
    port map (
            O => \N__12586\,
            I => \N__12583\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__12583\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_0\
        );

    \I__1292\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12576\
        );

    \I__1291\ : InMux
    port map (
            O => \N__12579\,
            I => \N__12569\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__12576\,
            I => \N__12566\
        );

    \I__1289\ : InMux
    port map (
            O => \N__12575\,
            I => \N__12557\
        );

    \I__1288\ : InMux
    port map (
            O => \N__12574\,
            I => \N__12557\
        );

    \I__1287\ : InMux
    port map (
            O => \N__12573\,
            I => \N__12557\
        );

    \I__1286\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12557\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__12569\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1284\ : Odrv4
    port map (
            O => \N__12566\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__12557\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1282\ : InMux
    port map (
            O => \N__12550\,
            I => \N__12547\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__12547\,
            I => \this_vga_signals.N_2_7_0\
        );

    \I__1280\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12540\
        );

    \I__1279\ : InMux
    port map (
            O => \N__12543\,
            I => \N__12537\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__12540\,
            I => \this_vga_signals.N_236\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__12537\,
            I => \this_vga_signals.N_236\
        );

    \I__1276\ : InMux
    port map (
            O => \N__12532\,
            I => \N__12529\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__12529\,
            I => \N__12525\
        );

    \I__1274\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12520\
        );

    \I__1273\ : Span4Mux_v
    port map (
            O => \N__12525\,
            I => \N__12517\
        );

    \I__1272\ : InMux
    port map (
            O => \N__12524\,
            I => \N__12514\
        );

    \I__1271\ : InMux
    port map (
            O => \N__12523\,
            I => \N__12511\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__12520\,
            I => \this_vga_signals.SUM_3_i_0_0_3\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__12517\,
            I => \this_vga_signals.SUM_3_i_0_0_3\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__12514\,
            I => \this_vga_signals.SUM_3_i_0_0_3\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__12511\,
            I => \this_vga_signals.SUM_3_i_0_0_3\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__12502\,
            I => \N__12499\
        );

    \I__1265\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12496\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__12496\,
            I => \N__12493\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__12493\,
            I => \N__12490\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__12490\,
            I => \this_vga_signals.g0_1\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__12487\,
            I => \this_vga_signals.un6_vvisibilitylt8_cascade_\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__12484\,
            I => \this_vga_signals.vvisibility_1_cascade_\
        );

    \I__1259\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12478\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__12478\,
            I => \N__12475\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__12475\,
            I => \this_vga_signals.vsync_1_3\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__12472\,
            I => \this_vga_signals.vsync_1_2_cascade_\
        );

    \I__1255\ : IoInMux
    port map (
            O => \N__12469\,
            I => \N__12466\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__12466\,
            I => \N__12463\
        );

    \I__1253\ : IoSpan4Mux
    port map (
            O => \N__12463\,
            I => \N__12460\
        );

    \I__1252\ : Span4Mux_s2_v
    port map (
            O => \N__12460\,
            I => \N__12457\
        );

    \I__1251\ : Sp12to4
    port map (
            O => \N__12457\,
            I => \N__12454\
        );

    \I__1250\ : Span12Mux_s10_v
    port map (
            O => \N__12454\,
            I => \N__12451\
        );

    \I__1249\ : Odrv12
    port map (
            O => \N__12451\,
            I => this_vga_signals_vsync_1_i
        );

    \I__1248\ : InMux
    port map (
            O => \N__12448\,
            I => \N__12440\
        );

    \I__1247\ : InMux
    port map (
            O => \N__12447\,
            I => \N__12437\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__12446\,
            I => \N__12434\
        );

    \I__1245\ : InMux
    port map (
            O => \N__12445\,
            I => \N__12431\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__12444\,
            I => \N__12428\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__12443\,
            I => \N__12425\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__12440\,
            I => \N__12420\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__12437\,
            I => \N__12420\
        );

    \I__1240\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12417\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__12431\,
            I => \N__12414\
        );

    \I__1238\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12409\
        );

    \I__1237\ : InMux
    port map (
            O => \N__12425\,
            I => \N__12409\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__12420\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__12417\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__12414\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__12409\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9\
        );

    \I__1232\ : InMux
    port map (
            O => \N__12400\,
            I => \N__12397\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__12397\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1\
        );

    \I__1230\ : InMux
    port map (
            O => \N__12394\,
            I => \N__12391\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__12391\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_7\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__12388\,
            I => \N__12384\
        );

    \I__1227\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12381\
        );

    \I__1226\ : InMux
    port map (
            O => \N__12384\,
            I => \N__12378\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__12381\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_8\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__12378\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_8\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__12373\,
            I => \N__12370\
        );

    \I__1222\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12367\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__12367\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_9\
        );

    \I__1220\ : InMux
    port map (
            O => \N__12364\,
            I => \N__12360\
        );

    \I__1219\ : InMux
    port map (
            O => \N__12363\,
            I => \N__12357\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__12360\,
            I => \N__12354\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__12357\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_6\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__12354\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_6\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__12349\,
            I => \this_vga_signals.SUM_3_i_0_0_3_cascade_\
        );

    \I__1214\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12342\
        );

    \I__1213\ : InMux
    port map (
            O => \N__12345\,
            I => \N__12339\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__12342\,
            I => \N__12333\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__12339\,
            I => \N__12333\
        );

    \I__1210\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12330\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__12333\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__12330\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__12325\,
            I => \N__12321\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__12324\,
            I => \N__12317\
        );

    \I__1205\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12314\
        );

    \I__1204\ : InMux
    port map (
            O => \N__12320\,
            I => \N__12310\
        );

    \I__1203\ : InMux
    port map (
            O => \N__12317\,
            I => \N__12307\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__12314\,
            I => \N__12304\
        );

    \I__1201\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12301\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__12310\,
            I => \N__12296\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__12307\,
            I => \N__12296\
        );

    \I__1198\ : Odrv12
    port map (
            O => \N__12304\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__12301\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__12296\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__12289\,
            I => \this_vga_signals.mult1_un61_sum_axb1_cascade_\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__12286\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_cascade_\
        );

    \I__1193\ : InMux
    port map (
            O => \N__12283\,
            I => \N__12280\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__12280\,
            I => \this_vga_signals.mult1_un75_sum_axb2_1\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__12277\,
            I => \this_vga_signals.N_236_cascade_\
        );

    \I__1190\ : InMux
    port map (
            O => \N__12274\,
            I => \N__12271\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__12271\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_0\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__12268\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__12265\,
            I => \this_vga_signals.N_3_2_1_cascade_\
        );

    \I__1186\ : InMux
    port map (
            O => \N__12262\,
            I => \N__12259\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__12259\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__12256\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_0_0_cascade_\
        );

    \I__1183\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12250\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__12250\,
            I => \this_vga_signals.g2_0_0\
        );

    \I__1181\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12244\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__12244\,
            I => \this_vga_signals.if_N_9_0_0\
        );

    \I__1179\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12237\
        );

    \I__1178\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12234\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__12237\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__12234\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__12229\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__12226\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_cascade_\
        );

    \I__1173\ : IoInMux
    port map (
            O => \N__12223\,
            I => \N__12220\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__12220\,
            I => \N__12217\
        );

    \I__1171\ : Odrv12
    port map (
            O => \N__12217\,
            I => this_vga_signals_vvisibility_i
        );

    \I__1170\ : InMux
    port map (
            O => \N__12214\,
            I => \N__12210\
        );

    \I__1169\ : InMux
    port map (
            O => \N__12213\,
            I => \N__12207\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__12210\,
            I => \N__12204\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__12207\,
            I => \this_vga_signals.N_5_i_5\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__12204\,
            I => \this_vga_signals.N_5_i_5\
        );

    \I__1165\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12196\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__12196\,
            I => \N__12193\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__12193\,
            I => \this_vga_signals.mult1_un82_sum_c3_0\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__12190\,
            I => \this_vga_signals.g0_4_cascade_\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__12187\,
            I => \this_vga_signals.g0_7_0_cascade_\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__12184\,
            I => \N__12181\
        );

    \I__1159\ : InMux
    port map (
            O => \N__12181\,
            I => \N__12178\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__12178\,
            I => \N__12175\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__12175\,
            I => \N__12172\
        );

    \I__1156\ : Sp12to4
    port map (
            O => \N__12172\,
            I => \N__12169\
        );

    \I__1155\ : Span12Mux_h
    port map (
            O => \N__12169\,
            I => \N__12166\
        );

    \I__1154\ : Odrv12
    port map (
            O => \N__12166\,
            I => \M_this_vga_signals_address_1\
        );

    \I__1153\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12160\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__12160\,
            I => \N__12157\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__12157\,
            I => \this_vga_ramdac.N_24_mux\
        );

    \I__1150\ : InMux
    port map (
            O => \N__12154\,
            I => \N__12150\
        );

    \I__1149\ : InMux
    port map (
            O => \N__12153\,
            I => \N__12147\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__12150\,
            I => \N__12144\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__12147\,
            I => \N__12141\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__12144\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__12141\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\
        );

    \I__1144\ : InMux
    port map (
            O => \N__12136\,
            I => \N__12133\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__12133\,
            I => \this_vga_signals.g1\
        );

    \I__1142\ : InMux
    port map (
            O => \N__12130\,
            I => \N__12127\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__12127\,
            I => \N__12124\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__12124\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_0_0\
        );

    \I__1139\ : InMux
    port map (
            O => \N__12121\,
            I => \N__12118\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__12118\,
            I => \this_vga_signals.un2_hsynclt6_0\
        );

    \I__1137\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12109\
        );

    \I__1136\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12109\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__12109\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_1\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__12106\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__12103\,
            I => \this_vga_signals.M_hcounter_d7lt7_0_cascade_\
        );

    \I__1132\ : InMux
    port map (
            O => \N__12100\,
            I => \N__12097\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__12097\,
            I => \this_vga_signals.M_hcounter_d7lto7_1\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__12094\,
            I => \this_vga_signals.mult1_un61_sum_0_3_cascade_\
        );

    \I__1129\ : IoInMux
    port map (
            O => \N__12091\,
            I => \N__12088\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__12088\,
            I => \N__12085\
        );

    \I__1127\ : Odrv12
    port map (
            O => \N__12085\,
            I => \this_vga_signals.N_614_1\
        );

    \I__1126\ : InMux
    port map (
            O => \N__12082\,
            I => \N__12079\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__12079\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_0\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__12076\,
            I => \this_vga_signals.g0_i_x4_0_cascade_\
        );

    \I__1123\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12070\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__12070\,
            I => \N__12067\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__12067\,
            I => \this_vga_signals.g0_i_x4_2\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__12064\,
            I => \this_vga_signals.N_931_1_cascade_\
        );

    \I__1119\ : IoInMux
    port map (
            O => \N__12061\,
            I => \N__12058\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__12058\,
            I => \N__12055\
        );

    \I__1117\ : Span12Mux_s8_v
    port map (
            O => \N__12055\,
            I => \N__12052\
        );

    \I__1116\ : Span12Mux_h
    port map (
            O => \N__12052\,
            I => \N__12048\
        );

    \I__1115\ : InMux
    port map (
            O => \N__12051\,
            I => \N__12045\
        );

    \I__1114\ : Odrv12
    port map (
            O => \N__12048\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI0JBR6Z0Z_9\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__12045\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI0JBR6Z0Z_9\
        );

    \I__1112\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12037\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__12037\,
            I => \this_vga_signals.un4_hsynclto3_0\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__12034\,
            I => \this_vga_signals.un2_hsynclt7_cascade_\
        );

    \I__1109\ : InMux
    port map (
            O => \N__12031\,
            I => \N__12028\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__12028\,
            I => \this_vga_signals.hsync_1_0\
        );

    \I__1107\ : IoInMux
    port map (
            O => \N__12025\,
            I => \N__12022\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__12022\,
            I => \N__12019\
        );

    \I__1105\ : Span4Mux_s0_v
    port map (
            O => \N__12019\,
            I => \N__12016\
        );

    \I__1104\ : Span4Mux_v
    port map (
            O => \N__12016\,
            I => \N__12013\
        );

    \I__1103\ : Span4Mux_v
    port map (
            O => \N__12013\,
            I => \N__12010\
        );

    \I__1102\ : Span4Mux_v
    port map (
            O => \N__12010\,
            I => \N__12007\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__12007\,
            I => this_vga_signals_hvisibility_i
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__12004\,
            I => \this_vga_signals.if_N_8_i_0_cascade_\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__12001\,
            I => \this_vga_signals.if_N_9_0_0_cascade_\
        );

    \I__1098\ : InMux
    port map (
            O => \N__11998\,
            I => \N__11994\
        );

    \I__1097\ : InMux
    port map (
            O => \N__11997\,
            I => \N__11991\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__11994\,
            I => \N__11988\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__11991\,
            I => \this_pixel_clk.M_counter_q_i_1\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__11988\,
            I => \this_pixel_clk.M_counter_q_i_1\
        );

    \I__1093\ : InMux
    port map (
            O => \N__11983\,
            I => \N__11978\
        );

    \I__1092\ : InMux
    port map (
            O => \N__11982\,
            I => \N__11975\
        );

    \I__1091\ : InMux
    port map (
            O => \N__11981\,
            I => \N__11972\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__11978\,
            I => \this_pixel_clk.M_counter_qZ0Z_0\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__11975\,
            I => \this_pixel_clk.M_counter_qZ0Z_0\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__11972\,
            I => \this_pixel_clk.M_counter_qZ0Z_0\
        );

    \I__1087\ : IoInMux
    port map (
            O => \N__11965\,
            I => \N__11962\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__11962\,
            I => \N__11959\
        );

    \I__1085\ : Span4Mux_s2_h
    port map (
            O => \N__11959\,
            I => \N__11956\
        );

    \I__1084\ : Sp12to4
    port map (
            O => \N__11956\,
            I => \N__11953\
        );

    \I__1083\ : Odrv12
    port map (
            O => \N__11953\,
            I => rgb_c_3
        );

    \I__1082\ : IoInMux
    port map (
            O => \N__11950\,
            I => \N__11947\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__11947\,
            I => \N__11944\
        );

    \I__1080\ : Span4Mux_s2_h
    port map (
            O => \N__11944\,
            I => \N__11941\
        );

    \I__1079\ : Span4Mux_v
    port map (
            O => \N__11941\,
            I => \N__11938\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__11938\,
            I => \N__11935\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__11935\,
            I => rgb_c_4
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__11932\,
            I => \N__11928\
        );

    \I__1075\ : InMux
    port map (
            O => \N__11931\,
            I => \N__11925\
        );

    \I__1074\ : InMux
    port map (
            O => \N__11928\,
            I => \N__11922\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__11925\,
            I => \this_vga_ramdac.N_2870_reto\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__11922\,
            I => \this_vga_ramdac.N_2870_reto\
        );

    \I__1071\ : IoInMux
    port map (
            O => \N__11917\,
            I => \N__11914\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__11914\,
            I => \N__11911\
        );

    \I__1069\ : Odrv12
    port map (
            O => \N__11911\,
            I => rgb_c_2
        );

    \I__1068\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11905\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__11905\,
            I => \this_vga_ramdac.i2_mux_0\
        );

    \I__1066\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11898\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__11901\,
            I => \N__11895\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__11898\,
            I => \N__11892\
        );

    \I__1063\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11889\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__11892\,
            I => \this_vga_ramdac.N_2875_reto\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__11889\,
            I => \this_vga_ramdac.N_2875_reto\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__11884\,
            I => \this_vga_signals.un4_hsynclto7_0_cascade_\
        );

    \I__1059\ : IoInMux
    port map (
            O => \N__11881\,
            I => \N__11878\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__11878\,
            I => \N__11875\
        );

    \I__1057\ : IoSpan4Mux
    port map (
            O => \N__11875\,
            I => \N__11872\
        );

    \I__1056\ : Span4Mux_s3_v
    port map (
            O => \N__11872\,
            I => \N__11869\
        );

    \I__1055\ : Sp12to4
    port map (
            O => \N__11869\,
            I => \N__11866\
        );

    \I__1054\ : Odrv12
    port map (
            O => \N__11866\,
            I => this_vga_signals_hsync_1_i
        );

    \I__1053\ : IoInMux
    port map (
            O => \N__11863\,
            I => \N__11860\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__11860\,
            I => \N__11857\
        );

    \I__1051\ : Span4Mux_s0_h
    port map (
            O => \N__11857\,
            I => \N__11854\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__11854\,
            I => \N__11851\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__11851\,
            I => port_nmib_0_i
        );

    \I__1048\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11845\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__11845\,
            I => \N__11842\
        );

    \I__1046\ : Span4Mux_v
    port map (
            O => \N__11842\,
            I => \N__11839\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__11839\,
            I => port_clk_c
        );

    \I__1044\ : InMux
    port map (
            O => \N__11836\,
            I => \N__11833\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__11833\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__1042\ : IoInMux
    port map (
            O => \N__11830\,
            I => \N__11827\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__11827\,
            I => \N__11824\
        );

    \I__1040\ : IoSpan4Mux
    port map (
            O => \N__11824\,
            I => \N__11821\
        );

    \I__1039\ : Span4Mux_s1_h
    port map (
            O => \N__11821\,
            I => \N__11818\
        );

    \I__1038\ : Span4Mux_v
    port map (
            O => \N__11818\,
            I => \N__11815\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__11815\,
            I => rgb_c_5
        );

    \I__1036\ : IoInMux
    port map (
            O => \N__11812\,
            I => \N__11809\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__11809\,
            I => \N__11806\
        );

    \I__1034\ : IoSpan4Mux
    port map (
            O => \N__11806\,
            I => \N__11803\
        );

    \I__1033\ : Span4Mux_s1_h
    port map (
            O => \N__11803\,
            I => \N__11800\
        );

    \I__1032\ : Odrv4
    port map (
            O => \N__11800\,
            I => port_data_rw_0_i
        );

    \I__1031\ : IoInMux
    port map (
            O => \N__11797\,
            I => \N__11794\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__11794\,
            I => \N__11791\
        );

    \I__1029\ : Span4Mux_s2_h
    port map (
            O => \N__11791\,
            I => \N__11788\
        );

    \I__1028\ : Sp12to4
    port map (
            O => \N__11788\,
            I => \N__11785\
        );

    \I__1027\ : Odrv12
    port map (
            O => \N__11785\,
            I => rgb_c_0
        );

    \I__1026\ : IoInMux
    port map (
            O => \N__11782\,
            I => \N__11779\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__11779\,
            I => \N__11776\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__11776\,
            I => rgb_c_1
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__11773\,
            I => \N__11770\
        );

    \I__1022\ : CascadeBuf
    port map (
            O => \N__11770\,
            I => \N__11767\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__11767\,
            I => \N__11764\
        );

    \I__1020\ : CascadeBuf
    port map (
            O => \N__11764\,
            I => \N__11761\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__11761\,
            I => \N__11758\
        );

    \I__1018\ : CascadeBuf
    port map (
            O => \N__11758\,
            I => \N__11755\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__11755\,
            I => \N__11752\
        );

    \I__1016\ : CascadeBuf
    port map (
            O => \N__11752\,
            I => \N__11749\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__11749\,
            I => \N__11746\
        );

    \I__1014\ : CascadeBuf
    port map (
            O => \N__11746\,
            I => \N__11743\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__11743\,
            I => \N__11740\
        );

    \I__1012\ : CascadeBuf
    port map (
            O => \N__11740\,
            I => \N__11737\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__11737\,
            I => \N__11734\
        );

    \I__1010\ : CascadeBuf
    port map (
            O => \N__11734\,
            I => \N__11731\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__11731\,
            I => \N__11728\
        );

    \I__1008\ : CascadeBuf
    port map (
            O => \N__11728\,
            I => \N__11725\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__11725\,
            I => \N__11722\
        );

    \I__1006\ : CascadeBuf
    port map (
            O => \N__11722\,
            I => \N__11719\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__11719\,
            I => \N__11716\
        );

    \I__1004\ : CascadeBuf
    port map (
            O => \N__11716\,
            I => \N__11713\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__11713\,
            I => \N__11710\
        );

    \I__1002\ : CascadeBuf
    port map (
            O => \N__11710\,
            I => \N__11707\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__11707\,
            I => \N__11704\
        );

    \I__1000\ : CascadeBuf
    port map (
            O => \N__11704\,
            I => \N__11701\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__11701\,
            I => \N__11698\
        );

    \I__998\ : CascadeBuf
    port map (
            O => \N__11698\,
            I => \N__11695\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__11695\,
            I => \N__11692\
        );

    \I__996\ : CascadeBuf
    port map (
            O => \N__11692\,
            I => \N__11689\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__11689\,
            I => \N__11686\
        );

    \I__994\ : CascadeBuf
    port map (
            O => \N__11686\,
            I => \N__11683\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__11683\,
            I => \N__11680\
        );

    \I__992\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11677\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__11677\,
            I => \N__11674\
        );

    \I__990\ : Span12Mux_h
    port map (
            O => \N__11674\,
            I => \N__11671\
        );

    \I__989\ : Span12Mux_h
    port map (
            O => \N__11671\,
            I => \N__11668\
        );

    \I__988\ : Odrv12
    port map (
            O => \N__11668\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__11665\,
            I => \N__11662\
        );

    \I__986\ : CascadeBuf
    port map (
            O => \N__11662\,
            I => \N__11659\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__11659\,
            I => \N__11656\
        );

    \I__984\ : CascadeBuf
    port map (
            O => \N__11656\,
            I => \N__11653\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__11653\,
            I => \N__11650\
        );

    \I__982\ : CascadeBuf
    port map (
            O => \N__11650\,
            I => \N__11647\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__11647\,
            I => \N__11644\
        );

    \I__980\ : CascadeBuf
    port map (
            O => \N__11644\,
            I => \N__11641\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__11641\,
            I => \N__11638\
        );

    \I__978\ : CascadeBuf
    port map (
            O => \N__11638\,
            I => \N__11635\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__11635\,
            I => \N__11632\
        );

    \I__976\ : CascadeBuf
    port map (
            O => \N__11632\,
            I => \N__11629\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__11629\,
            I => \N__11626\
        );

    \I__974\ : CascadeBuf
    port map (
            O => \N__11626\,
            I => \N__11623\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__11623\,
            I => \N__11620\
        );

    \I__972\ : CascadeBuf
    port map (
            O => \N__11620\,
            I => \N__11617\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__11617\,
            I => \N__11614\
        );

    \I__970\ : CascadeBuf
    port map (
            O => \N__11614\,
            I => \N__11611\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__11611\,
            I => \N__11608\
        );

    \I__968\ : CascadeBuf
    port map (
            O => \N__11608\,
            I => \N__11605\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__11605\,
            I => \N__11602\
        );

    \I__966\ : CascadeBuf
    port map (
            O => \N__11602\,
            I => \N__11599\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__11599\,
            I => \N__11596\
        );

    \I__964\ : CascadeBuf
    port map (
            O => \N__11596\,
            I => \N__11593\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__11593\,
            I => \N__11590\
        );

    \I__962\ : CascadeBuf
    port map (
            O => \N__11590\,
            I => \N__11587\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__11587\,
            I => \N__11584\
        );

    \I__960\ : CascadeBuf
    port map (
            O => \N__11584\,
            I => \N__11581\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__11581\,
            I => \N__11578\
        );

    \I__958\ : CascadeBuf
    port map (
            O => \N__11578\,
            I => \N__11575\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__11575\,
            I => \N__11572\
        );

    \I__956\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11569\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__954\ : Span4Mux_h
    port map (
            O => \N__11566\,
            I => \N__11563\
        );

    \I__953\ : Sp12to4
    port map (
            O => \N__11563\,
            I => \N__11560\
        );

    \I__952\ : Span12Mux_s3_v
    port map (
            O => \N__11560\,
            I => \N__11557\
        );

    \I__951\ : Span12Mux_h
    port map (
            O => \N__11557\,
            I => \N__11554\
        );

    \I__950\ : Odrv12
    port map (
            O => \N__11554\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__11551\,
            I => \N__11548\
        );

    \I__948\ : CascadeBuf
    port map (
            O => \N__11548\,
            I => \N__11545\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__11545\,
            I => \N__11542\
        );

    \I__946\ : CascadeBuf
    port map (
            O => \N__11542\,
            I => \N__11539\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__11539\,
            I => \N__11536\
        );

    \I__944\ : CascadeBuf
    port map (
            O => \N__11536\,
            I => \N__11533\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__11533\,
            I => \N__11530\
        );

    \I__942\ : CascadeBuf
    port map (
            O => \N__11530\,
            I => \N__11527\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__11527\,
            I => \N__11524\
        );

    \I__940\ : CascadeBuf
    port map (
            O => \N__11524\,
            I => \N__11521\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__11521\,
            I => \N__11518\
        );

    \I__938\ : CascadeBuf
    port map (
            O => \N__11518\,
            I => \N__11515\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__11515\,
            I => \N__11512\
        );

    \I__936\ : CascadeBuf
    port map (
            O => \N__11512\,
            I => \N__11509\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__11509\,
            I => \N__11506\
        );

    \I__934\ : CascadeBuf
    port map (
            O => \N__11506\,
            I => \N__11503\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__11503\,
            I => \N__11500\
        );

    \I__932\ : CascadeBuf
    port map (
            O => \N__11500\,
            I => \N__11497\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__11497\,
            I => \N__11494\
        );

    \I__930\ : CascadeBuf
    port map (
            O => \N__11494\,
            I => \N__11491\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__11491\,
            I => \N__11488\
        );

    \I__928\ : CascadeBuf
    port map (
            O => \N__11488\,
            I => \N__11485\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__11485\,
            I => \N__11482\
        );

    \I__926\ : CascadeBuf
    port map (
            O => \N__11482\,
            I => \N__11479\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__11479\,
            I => \N__11476\
        );

    \I__924\ : CascadeBuf
    port map (
            O => \N__11476\,
            I => \N__11473\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__11473\,
            I => \N__11470\
        );

    \I__922\ : CascadeBuf
    port map (
            O => \N__11470\,
            I => \N__11467\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__11467\,
            I => \N__11464\
        );

    \I__920\ : CascadeBuf
    port map (
            O => \N__11464\,
            I => \N__11461\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__11461\,
            I => \N__11458\
        );

    \I__918\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11455\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__11455\,
            I => \N__11452\
        );

    \I__916\ : Span4Mux_s2_v
    port map (
            O => \N__11452\,
            I => \N__11449\
        );

    \I__915\ : Sp12to4
    port map (
            O => \N__11449\,
            I => \N__11446\
        );

    \I__914\ : Span12Mux_s6_h
    port map (
            O => \N__11446\,
            I => \N__11443\
        );

    \I__913\ : Span12Mux_h
    port map (
            O => \N__11443\,
            I => \N__11440\
        );

    \I__912\ : Odrv12
    port map (
            O => \N__11440\,
            I => \M_this_ppu_sprites_addr_7\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__11437\,
            I => \N__11434\
        );

    \I__910\ : CascadeBuf
    port map (
            O => \N__11434\,
            I => \N__11431\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__11431\,
            I => \N__11428\
        );

    \I__908\ : CascadeBuf
    port map (
            O => \N__11428\,
            I => \N__11425\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__11425\,
            I => \N__11422\
        );

    \I__906\ : CascadeBuf
    port map (
            O => \N__11422\,
            I => \N__11419\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__11419\,
            I => \N__11416\
        );

    \I__904\ : CascadeBuf
    port map (
            O => \N__11416\,
            I => \N__11413\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__11413\,
            I => \N__11410\
        );

    \I__902\ : CascadeBuf
    port map (
            O => \N__11410\,
            I => \N__11407\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__11407\,
            I => \N__11404\
        );

    \I__900\ : CascadeBuf
    port map (
            O => \N__11404\,
            I => \N__11401\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__11401\,
            I => \N__11398\
        );

    \I__898\ : CascadeBuf
    port map (
            O => \N__11398\,
            I => \N__11395\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__11395\,
            I => \N__11392\
        );

    \I__896\ : CascadeBuf
    port map (
            O => \N__11392\,
            I => \N__11389\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__11389\,
            I => \N__11386\
        );

    \I__894\ : CascadeBuf
    port map (
            O => \N__11386\,
            I => \N__11383\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__11383\,
            I => \N__11380\
        );

    \I__892\ : CascadeBuf
    port map (
            O => \N__11380\,
            I => \N__11377\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__11377\,
            I => \N__11374\
        );

    \I__890\ : CascadeBuf
    port map (
            O => \N__11374\,
            I => \N__11371\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__11371\,
            I => \N__11368\
        );

    \I__888\ : CascadeBuf
    port map (
            O => \N__11368\,
            I => \N__11365\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__11365\,
            I => \N__11362\
        );

    \I__886\ : CascadeBuf
    port map (
            O => \N__11362\,
            I => \N__11359\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__11359\,
            I => \N__11356\
        );

    \I__884\ : CascadeBuf
    port map (
            O => \N__11356\,
            I => \N__11353\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__11353\,
            I => \N__11350\
        );

    \I__882\ : CascadeBuf
    port map (
            O => \N__11350\,
            I => \N__11347\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__11347\,
            I => \N__11344\
        );

    \I__880\ : InMux
    port map (
            O => \N__11344\,
            I => \N__11341\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__11341\,
            I => \N__11338\
        );

    \I__878\ : Span4Mux_s2_v
    port map (
            O => \N__11338\,
            I => \N__11335\
        );

    \I__877\ : Sp12to4
    port map (
            O => \N__11335\,
            I => \N__11332\
        );

    \I__876\ : Span12Mux_h
    port map (
            O => \N__11332\,
            I => \N__11329\
        );

    \I__875\ : Odrv12
    port map (
            O => \N__11329\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__11326\,
            I => \N__11323\
        );

    \I__873\ : CascadeBuf
    port map (
            O => \N__11323\,
            I => \N__11320\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__11320\,
            I => \N__11317\
        );

    \I__871\ : CascadeBuf
    port map (
            O => \N__11317\,
            I => \N__11314\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__11314\,
            I => \N__11311\
        );

    \I__869\ : CascadeBuf
    port map (
            O => \N__11311\,
            I => \N__11308\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__11308\,
            I => \N__11305\
        );

    \I__867\ : CascadeBuf
    port map (
            O => \N__11305\,
            I => \N__11302\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__11302\,
            I => \N__11299\
        );

    \I__865\ : CascadeBuf
    port map (
            O => \N__11299\,
            I => \N__11296\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__11296\,
            I => \N__11293\
        );

    \I__863\ : CascadeBuf
    port map (
            O => \N__11293\,
            I => \N__11290\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__11290\,
            I => \N__11287\
        );

    \I__861\ : CascadeBuf
    port map (
            O => \N__11287\,
            I => \N__11284\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__11284\,
            I => \N__11281\
        );

    \I__859\ : CascadeBuf
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__11278\,
            I => \N__11275\
        );

    \I__857\ : CascadeBuf
    port map (
            O => \N__11275\,
            I => \N__11272\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__11272\,
            I => \N__11269\
        );

    \I__855\ : CascadeBuf
    port map (
            O => \N__11269\,
            I => \N__11266\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__11266\,
            I => \N__11263\
        );

    \I__853\ : CascadeBuf
    port map (
            O => \N__11263\,
            I => \N__11260\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__11260\,
            I => \N__11257\
        );

    \I__851\ : CascadeBuf
    port map (
            O => \N__11257\,
            I => \N__11254\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__11254\,
            I => \N__11251\
        );

    \I__849\ : CascadeBuf
    port map (
            O => \N__11251\,
            I => \N__11248\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__11248\,
            I => \N__11245\
        );

    \I__847\ : CascadeBuf
    port map (
            O => \N__11245\,
            I => \N__11242\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__11242\,
            I => \N__11239\
        );

    \I__845\ : CascadeBuf
    port map (
            O => \N__11239\,
            I => \N__11236\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__11236\,
            I => \N__11233\
        );

    \I__843\ : InMux
    port map (
            O => \N__11233\,
            I => \N__11230\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__11230\,
            I => \N__11227\
        );

    \I__841\ : Span4Mux_v
    port map (
            O => \N__11227\,
            I => \N__11224\
        );

    \I__840\ : Span4Mux_h
    port map (
            O => \N__11224\,
            I => \N__11221\
        );

    \I__839\ : Sp12to4
    port map (
            O => \N__11221\,
            I => \N__11218\
        );

    \I__838\ : Span12Mux_h
    port map (
            O => \N__11218\,
            I => \N__11215\
        );

    \I__837\ : Odrv12
    port map (
            O => \N__11215\,
            I => \M_this_map_ram_read_data_4\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_23_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_17_0_\
        );

    \IN_MUX_bfv_23_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_data_count_q_cry_7\,
            carryinitout => \bfn_23_18_0_\
        );

    \IN_MUX_bfv_10_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_11_0_\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_10_12_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_sprites_address_q_cry_7\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_19_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_22_0_\
        );

    \IN_MUX_bfv_19_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_map_address_q_cry_7\,
            carryinitout => \bfn_19_23_0_\
        );

    \IN_MUX_bfv_22_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_20_0_\
        );

    \IN_MUX_bfv_22_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_external_address_q_cry_7\,
            carryinitout => \bfn_22_21_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILD847_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12091\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_614_1_g\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI0JBR6_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12061\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_931_g\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__27493\,
            GLOBALBUFFEROUTPUT => \M_this_reset_cond_out_g_0\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21412\,
            GLOBALBUFFEROUTPUT => \N_989_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIOJ6UA_8_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17008\,
            in2 => \_gnd_net_\,
            in3 => \N__21642\,
            lcout => port_nmib_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11848\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11836\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11902\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.port_data_rw_0_i_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__25287\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21652\,
            lcout => port_data_rw_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11931\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15373\,
            in2 => \_gnd_net_\,
            in3 => \N__13825\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13848\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15841\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13873\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13849\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_0_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11982\,
            lcout => \this_pixel_clk.M_counter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32028\,
            ce => 'H',
            sr => \N__32393\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__12163\,
            in1 => \N__27502\,
            in2 => \N__11932\,
            in3 => \N__15886\,
            lcout => \this_vga_ramdac.N_2870_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100100101"
        )
    port map (
            in0 => \N__16868\,
            in1 => \N__16816\,
            in2 => \N__16678\,
            in3 => \N__16753\,
            lcout => \this_vga_ramdac.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13846\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__11908\,
            in1 => \N__27497\,
            in2 => \N__11901\,
            in3 => \N__15885\,
            lcout => \this_vga_ramdac.N_2875_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIADGD1_2_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__12040\,
            in1 => \N__13005\,
            in2 => \N__13225\,
            in3 => \N__12915\,
            lcout => OPEN,
            ltout => \this_vga_signals.un4_hsynclto7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIF7AC4_8_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__13614\,
            in1 => \N__12031\,
            in2 => \N__11884\,
            in3 => \N__12834\,
            lcout => this_vga_signals_hsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNINT9T1_6_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12916\,
            in1 => \N__12121\,
            in2 => \N__13009\,
            in3 => \N__12835\,
            lcout => OPEN,
            ltout => \this_vga_signals.un2_hsynclt7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI73DH2_9_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__13534\,
            in1 => \N__13613\,
            in2 => \N__12034\,
            in3 => \N__12726\,
            lcout => \this_vga_signals.hsync_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__13533\,
            in1 => \N__13612\,
            in2 => \_gnd_net_\,
            in3 => \N__12725\,
            lcout => this_vga_signals_hvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__11997\,
            in1 => \N__11983\,
            in2 => \_gnd_net_\,
            in3 => \N__32437\,
            lcout => \this_pixel_clk.M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32025\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110110110100"
        )
    port map (
            in0 => \N__13000\,
            in1 => \N__13111\,
            in2 => \N__12324\,
            in3 => \N__14010\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_8_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13217\,
            in2 => \N__12004\,
            in3 => \N__13330\,
            lcout => \this_vga_signals.if_N_9_0_0\,
            ltout => \this_vga_signals.if_N_9_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_m2_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100011101"
        )
    port map (
            in0 => \N__13218\,
            in1 => \N__12213\,
            in2 => \N__12001\,
            in3 => \N__12073\,
            lcout => \this_vga_signals.mult1_un82_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_RNILQS8_1_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__11998\,
            in1 => \N__11981\,
            in2 => \_gnd_net_\,
            in3 => \N__32427\,
            lcout => \M_counter_q_RNILQS8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_3_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__12345\,
            in1 => \N__12448\,
            in2 => \_gnd_net_\,
            in3 => \N__12153\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_8_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12115\,
            in1 => \N__12082\,
            in2 => \N__12094\,
            in3 => \N__14396\,
            lcout => \this_vga_signals.N_5_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILD847_9_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__14636\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12051\,
            lcout => \this_vga_signals.N_614_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_5_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011011101"
        )
    port map (
            in0 => \N__12114\,
            in1 => \N__12914\,
            in2 => \_gnd_net_\,
            in3 => \N__12998\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001111001001"
        )
    port map (
            in0 => \N__12999\,
            in1 => \N__12313\,
            in2 => \N__13129\,
            in3 => \N__14011\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_x4_0_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12913\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13104\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_x4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_x4_2_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__12833\,
            in1 => \N__12543\,
            in2 => \N__12076\,
            in3 => \N__12532\,
            lcout => \this_vga_signals.g0_i_x4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIST9Q2_9_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14650\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14475\,
            lcout => \this_vga_signals.N_931_1\,
            ltout => \this_vga_signals.N_931_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI0JBR6_9_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__14259\,
            in1 => \N__17433\,
            in2 => \N__12064\,
            in3 => \N__15999\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNI0JBR6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m5_i_a4_0_1_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13106\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13329\,
            lcout => \this_vga_signals.un4_hsynclto3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13328\,
            in1 => \N__13222\,
            in2 => \N__13273\,
            in3 => \N__13105\,
            lcout => \this_vga_signals.un2_hsynclt6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001010110000"
        )
    port map (
            in0 => \N__12832\,
            in1 => \N__12912\,
            in2 => \N__12446\,
            in3 => \N__14304\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIHO633_9_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13415\,
            in2 => \_gnd_net_\,
            in3 => \N__14664\,
            lcout => \this_vga_signals.N_614_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12523\,
            in1 => \N__12262\,
            in2 => \_gnd_net_\,
            in3 => \N__12400\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__12338\,
            in1 => \_gnd_net_\,
            in2 => \N__12106\,
            in3 => \N__12445\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__13195\,
            in1 => \N__13234\,
            in2 => \N__13128\,
            in3 => \N__13004\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_d7lt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI73DH2_0_9_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__12100\,
            in1 => \N__13608\,
            in2 => \N__12103\,
            in3 => \N__13532\,
            lcout => \this_vga_signals.M_hcounter_d7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI11GM_7_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12898\,
            in1 => \N__12721\,
            in2 => \_gnd_net_\,
            in3 => \N__12823\,
            lcout => \this_vga_signals.M_hcounter_d7lto7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_7_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12685\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32048\,
            ce => \N__13472\,
            sr => \N__13431\
        );

    \this_vga_signals.M_hcounter_q_esr_8_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13570\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32048\,
            ce => \N__13472\,
            sr => \N__13431\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_8_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17029\,
            lcout => this_vga_signals_vvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_4_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12136\,
            in1 => \N__12320\,
            in2 => \N__12502\,
            in3 => \N__12214\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_7_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12199\,
            in1 => \N__12658\,
            in2 => \N__12190\,
            in3 => \N__13384\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIQFEIV5_9_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010000010"
        )
    port map (
            in0 => \N__20963\,
            in1 => \N__12130\,
            in2 => \N__12187\,
            in3 => \N__13348\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010111011"
        )
    port map (
            in0 => \N__13119\,
            in1 => \N__13207\,
            in2 => \_gnd_net_\,
            in3 => \N__12580\,
            lcout => \this_vga_signals.mult1_un75_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__16815\,
            in1 => \N__16666\,
            in2 => \_gnd_net_\,
            in3 => \N__16751\,
            lcout => \this_vga_ramdac.N_24_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000101111"
        )
    port map (
            in0 => \N__12253\,
            in1 => \N__12154\,
            in2 => \N__13130\,
            in3 => \N__13001\,
            lcout => \this_vga_signals.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIUAKU9_4_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001001001011"
        )
    port map (
            in0 => \N__13002\,
            in1 => \N__13118\,
            in2 => \N__12325\,
            in3 => \N__14013\,
            lcout => \this_vga_signals.M_hcounter_q_RNIUAKU9Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_0_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111011010"
        )
    port map (
            in0 => \N__13003\,
            in1 => \N__12572\,
            in2 => \N__13131\,
            in3 => \N__14012\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_3_0_0\,
            ltout => \this_vga_signals.mult1_un75_sum_ac0_3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010010110"
        )
    port map (
            in0 => \N__12573\,
            in1 => \N__12241\,
            in2 => \N__12256\,
            in3 => \N__13341\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g2_0_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12447\,
            in2 => \_gnd_net_\,
            in3 => \N__12346\,
            lcout => \this_vga_signals.g2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100101101111"
        )
    port map (
            in0 => \N__12575\,
            in1 => \N__13126\,
            in2 => \N__13223\,
            in3 => \N__12247\,
            lcout => \this_vga_signals.mult1_un82_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIB3UCP_1_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011100"
        )
    port map (
            in0 => \N__13317\,
            in1 => \N__13209\,
            in2 => \N__13132\,
            in3 => \N__12574\,
            lcout => \this_vga_signals.d_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIVPQGA_1_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__13318\,
            in1 => \N__13208\,
            in2 => \_gnd_net_\,
            in3 => \N__12240\,
            lcout => \this_vga_signals.d_N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010100101011"
        )
    port map (
            in0 => \N__16873\,
            in1 => \N__16814\,
            in2 => \N__16674\,
            in3 => \N__16747\,
            lcout => \this_vga_ramdac.m19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_1_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001010110100"
        )
    port map (
            in0 => \N__12886\,
            in1 => \N__20912\,
            in2 => \N__13067\,
            in3 => \N__12971\,
            lcout => \this_vga_signals.mult1_un75_sum_axb2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001010110000"
        )
    port map (
            in0 => \N__12824\,
            in1 => \N__12883\,
            in2 => \N__12443\,
            in3 => \N__14302\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010101111"
        )
    port map (
            in0 => \N__12885\,
            in1 => \_gnd_net_\,
            in2 => \N__12229\,
            in3 => \N__12972\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un61_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13110\,
            in1 => \N__14392\,
            in2 => \N__12226\,
            in3 => \N__14366\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__14367\,
            in1 => \_gnd_net_\,
            in2 => \N__14400\,
            in3 => \N__14415\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000110000011"
        )
    port map (
            in0 => \N__12825\,
            in1 => \N__12884\,
            in2 => \N__12444\,
            in3 => \N__14303\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1\,
            ltout => \this_vga_signals.mult1_un61_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011111000001"
        )
    port map (
            in0 => \N__13042\,
            in1 => \N__12970\,
            in2 => \N__12289\,
            in3 => \N__13994\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20913\,
            in1 => \N__12274\,
            in2 => \N__12286\,
            in3 => \N__12283\,
            lcout => \this_vga_signals.mult1_un75_sum_axb2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__12719\,
            in1 => \N__12793\,
            in2 => \N__13626\,
            in3 => \N__13509\,
            lcout => \this_vga_signals.N_236\,
            ltout => \this_vga_signals.N_236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__12880\,
            in1 => \N__12797\,
            in2 => \N__12277\,
            in3 => \N__12524\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_3_0\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20911\,
            in2 => \N__12268\,
            in3 => \N__13993\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNIOIVT_6_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011100011111"
        )
    port map (
            in0 => \N__12364\,
            in1 => \N__13506\,
            in2 => \N__12388\,
            in3 => \N__12717\,
            lcout => \this_vga_signals.N_3_2_1\,
            ltout => \this_vga_signals.N_3_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100011000000"
        )
    port map (
            in0 => \N__12950\,
            in1 => \N__12792\,
            in2 => \N__12265\,
            in3 => \N__12878\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100101100101"
        )
    port map (
            in0 => \N__12791\,
            in1 => \N__13507\,
            in2 => \N__13625\,
            in3 => \N__12718\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101110000011"
        )
    port map (
            in0 => \N__12951\,
            in1 => \N__12879\,
            in2 => \N__12817\,
            in3 => \N__14301\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI43BG3_9_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__13618\,
            in1 => \N__13508\,
            in2 => \N__17018\,
            in3 => \N__12720\,
            lcout => \M_this_vga_ramdac_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_8_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13563\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32046\,
            ce => \N__13476\,
            sr => \N__13436\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_7_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12678\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32046\,
            ce => \N__13476\,
            sr => \N__13436\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_9_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13546\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32046\,
            ce => \N__13476\,
            sr => \N__13436\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_6_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12742\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32046\,
            ce => \N__13476\,
            sr => \N__13436\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNIIL511_7_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001001000"
        )
    port map (
            in0 => \N__12394\,
            in1 => \N__12387\,
            in2 => \N__12373\,
            in3 => \N__12363\,
            lcout => \this_vga_signals.SUM_3_i_0_0_3\,
            ltout => \this_vga_signals.SUM_3_i_0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001011101"
        )
    port map (
            in0 => \N__12881\,
            in1 => \N__12798\,
            in2 => \N__12349\,
            in3 => \N__12952\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_6_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12741\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32046\,
            ce => \N__13476\,
            sr => \N__13436\
        );

    \this_vga_signals.un4_haddress_g0_1_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__12882\,
            in1 => \N__12544\,
            in2 => \N__12826\,
            in3 => \N__12528\,
            lcout => \this_vga_signals.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIJELD1_8_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15998\,
            in1 => \N__19230\,
            in2 => \N__18129\,
            in3 => \N__16494\,
            lcout => \this_vga_signals.vsync_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__19233\,
            in1 => \N__18089\,
            in2 => \_gnd_net_\,
            in3 => \N__19701\,
            lcout => OPEN,
            ltout => \this_vga_signals.un6_vvisibilitylt8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI81G42_7_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000010001"
        )
    port map (
            in0 => \N__18090\,
            in1 => \N__16500\,
            in2 => \N__12487\,
            in3 => \N__16571\,
            lcout => OPEN,
            ltout => \this_vga_signals.vvisibility_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_8_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000101"
        )
    port map (
            in0 => \N__15997\,
            in1 => \N__16501\,
            in2 => \N__12484\,
            in3 => \N__14140\,
            lcout => this_vga_signals_vvisibility,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19708\,
            in1 => \N__16502\,
            in2 => \N__18128\,
            in3 => \N__16587\,
            lcout => \this_vga_signals.M_vcounter_d7lto8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__17818\,
            in1 => \N__19246\,
            in2 => \N__19018\,
            in3 => \N__18550\,
            lcout => OPEN,
            ltout => \this_vga_signals.vsync_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIUAQ3_7_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__19709\,
            in1 => \N__12481\,
            in2 => \N__12472\,
            in3 => \N__16588\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13379\,
            in2 => \_gnd_net_\,
            in3 => \N__13360\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m7_0_x4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100010111"
        )
    port map (
            in0 => \N__13315\,
            in1 => \N__13263\,
            in2 => \N__12664\,
            in3 => \N__12656\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100011011"
        )
    port map (
            in0 => \N__13914\,
            in1 => \N__13316\,
            in2 => \N__12661\,
            in3 => \N__13224\,
            lcout => \this_vga_signals.mult1_un89_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13380\,
            in1 => \N__12657\,
            in2 => \N__12643\,
            in3 => \N__13913\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI32C8PD_9_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20962\,
            in1 => \N__12586\,
            in2 => \N__12634\,
            in3 => \N__12631\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101000100"
        )
    port map (
            in0 => \N__12610\,
            in1 => \N__12604\,
            in2 => \N__12598\,
            in3 => \N__12550\,
            lcout => \this_vga_signals.mult1_un89_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m5_i_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001100010"
        )
    port map (
            in0 => \N__13314\,
            in1 => \N__13213\,
            in2 => \N__13127\,
            in3 => \N__12579\,
            lcout => \this_vga_signals.N_2_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13264\,
            in2 => \N__14718\,
            in3 => \N__13319\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32029\,
            ce => 'H',
            sr => \N__13432\
        );

    \this_vga_signals.M_hcounter_q_0_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__13265\,
            in1 => \N__14706\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32029\,
            ce => 'H',
            sr => \N__13432\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_d_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13177\,
            in1 => \N__13378\,
            in2 => \_gnd_net_\,
            in3 => \N__13359\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_3_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__13259\,
            in1 => \N__13310\,
            in2 => \N__13269\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_d7lt4\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14691\,
            in1 => \N__13194\,
            in2 => \_gnd_net_\,
            in3 => \N__13135\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__32038\,
            ce => 'H',
            sr => \N__13443\
        );

    \this_vga_signals.M_hcounter_q_3_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14689\,
            in1 => \N__13066\,
            in2 => \_gnd_net_\,
            in3 => \N__13012\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__32038\,
            ce => 'H',
            sr => \N__13443\
        );

    \this_vga_signals.M_hcounter_q_4_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14692\,
            in1 => \N__12997\,
            in2 => \_gnd_net_\,
            in3 => \N__12919\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__32038\,
            ce => 'H',
            sr => \N__13443\
        );

    \this_vga_signals.M_hcounter_q_5_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14690\,
            in1 => \N__12897\,
            in2 => \_gnd_net_\,
            in3 => \N__12838\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__32038\,
            ce => 'H',
            sr => \N__13443\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12813\,
            in2 => \_gnd_net_\,
            in3 => \N__12733\,
            lcout => \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12730\,
            in2 => \_gnd_net_\,
            in3 => \N__12667\,
            lcout => \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13627\,
            in2 => \_gnd_net_\,
            in3 => \N__13552\,
            lcout => \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13525\,
            in2 => \_gnd_net_\,
            in3 => \N__13549\,
            lcout => \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13545\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32041\,
            ce => \N__13477\,
            sr => \N__13444\
        );

    \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__17305\,
            in1 => \N__15072\,
            in2 => \_gnd_net_\,
            in3 => \N__15325\,
            lcout => \this_vga_signals.g0_31_N_4L6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19475\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17306\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_11_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19750\,
            in1 => \N__16140\,
            in2 => \N__13387\,
            in3 => \N__17225\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14998\,
            in2 => \_gnd_net_\,
            in3 => \N__14968\,
            lcout => \this_vga_signals.vaddress_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14788\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31980\,
            ce => \N__15140\,
            sr => \N__15114\
        );

    \this_vga_signals.un5_vaddress_g0_34_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__16578\,
            in1 => \N__15081\,
            in2 => \N__16504\,
            in3 => \N__15960\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m8_0_a3_1_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000011101"
        )
    port map (
            in0 => \N__13657\,
            in1 => \N__13648\,
            in2 => \N__13651\,
            in3 => \N__17179\,
            lcout => \this_vga_signals.g0_31_N_5L8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_31_N_3L3_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19615\,
            in2 => \_gnd_net_\,
            in3 => \N__19474\,
            lcout => \this_vga_signals.g0_31_N_3L3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14787\,
            lcout => \this_vga_signals.M_vcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31980\,
            ce => \N__15140\,
            sr => \N__15114\
        );

    \this_vga_signals.un5_vaddress_g3_3_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__18042\,
            in1 => \N__19617\,
            in2 => \_gnd_net_\,
            in3 => \N__19458\,
            lcout => \this_vga_signals.g3_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_32_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110110110111"
        )
    port map (
            in0 => \N__16498\,
            in1 => \N__16585\,
            in2 => \N__18115\,
            in3 => \N__15975\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m8_0_a3_1_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_8_0_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__13761\,
            in1 => \N__13642\,
            in2 => \N__13636\,
            in3 => \N__17211\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_27_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__19131\,
            in1 => \N__17675\,
            in2 => \N__13633\,
            in3 => \N__18394\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19616\,
            in2 => \_gnd_net_\,
            in3 => \N__19462\,
            lcout => \this_vga_signals.vaddress_2_5\,
            ltout => \this_vga_signals.vaddress_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000101001001"
        )
    port map (
            in0 => \N__17943\,
            in1 => \N__17224\,
            in2 => \N__13630\,
            in3 => \N__16054\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17303\,
            in2 => \_gnd_net_\,
            in3 => \N__15322\,
            lcout => \this_vga_signals.g1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__17304\,
            in1 => \_gnd_net_\,
            in2 => \N__19508\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.vaddress_6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_19_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__15990\,
            in1 => \N__16469\,
            in2 => \N__18083\,
            in3 => \N__16570\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14812\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31992\,
            ce => \N__15138\,
            sr => \N__15115\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14839\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31992\,
            ce => \N__15138\,
            sr => \N__15115\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__18031\,
            in1 => \N__19463\,
            in2 => \_gnd_net_\,
            in3 => \N__17331\,
            lcout => \this_vga_signals.vaddress_3_0_6\,
            ltout => \this_vga_signals.vaddress_3_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_33_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17204\,
            in2 => \N__13669\,
            in3 => \N__17942\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_1_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111001101"
        )
    port map (
            in0 => \N__18395\,
            in1 => \N__19228\,
            in2 => \N__13666\,
            in3 => \N__19643\,
            lcout => \this_vga_signals.g1_1_1\,
            ltout => \this_vga_signals.g1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_2_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13750\,
            in1 => \N__18231\,
            in2 => \N__13663\,
            in3 => \N__18396\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_x4_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100101101"
        )
    port map (
            in0 => \N__19229\,
            in1 => \N__18991\,
            in2 => \N__13660\,
            in3 => \N__14182\,
            lcout => \this_vga_signals.g0_i_x4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__18026\,
            in1 => \N__19641\,
            in2 => \_gnd_net_\,
            in3 => \N__19455\,
            lcout => \this_vga_signals.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_28_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010010011001"
        )
    port map (
            in0 => \N__13765\,
            in1 => \N__17219\,
            in2 => \N__13744\,
            in3 => \N__17940\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19642\,
            in2 => \_gnd_net_\,
            in3 => \N__19457\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_36_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010011000011"
        )
    port map (
            in0 => \N__13743\,
            in1 => \N__17218\,
            in2 => \N__13729\,
            in3 => \N__17941\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i_1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_1_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__18027\,
            in1 => \N__19456\,
            in2 => \_gnd_net_\,
            in3 => \N__17330\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_3_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_22_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010000"
        )
    port map (
            in0 => \N__16198\,
            in1 => \N__17217\,
            in2 => \N__13726\,
            in3 => \N__17939\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__23196\,
            in1 => \N__13675\,
            in2 => \N__14059\,
            in3 => \N__29674\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__14023\,
            in1 => \N__23197\,
            in2 => \N__13723\,
            in3 => \N__13771\,
            lcout => \M_this_ppu_vram_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27804\,
            in1 => \N__13702\,
            in2 => \_gnd_net_\,
            in3 => \N__13687\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27801\,
            in1 => \N__14086\,
            in2 => \_gnd_net_\,
            in3 => \N__14077\,
            lcout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14050\,
            in1 => \N__14038\,
            in2 => \_gnd_net_\,
            in3 => \N__27802\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIL26KA_9_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20982\,
            in2 => \_gnd_net_\,
            in3 => \N__14017\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13948\,
            in1 => \N__13930\,
            in2 => \_gnd_net_\,
            in3 => \N__27803\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIC813H3_9_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20981\,
            in2 => \_gnd_net_\,
            in3 => \N__13918\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__13885\,
            in1 => \N__27489\,
            in2 => \N__13866\,
            in3 => \N__15874\,
            lcout => \this_vga_ramdac.N_2874_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_ret_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__20999\,
            in1 => \N__13813\,
            in2 => \N__27501\,
            in3 => \N__15875\,
            lcout => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13798\,
            in1 => \N__13780\,
            in2 => \_gnd_net_\,
            in3 => \N__27805\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14693\,
            in1 => \N__18572\,
            in2 => \N__14536\,
            in3 => \N__14535\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_11_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__31954\,
            ce => 'H',
            sr => \N__15108\
        );

    \this_vga_signals.M_vcounter_q_1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14714\,
            in1 => \N__18513\,
            in2 => \_gnd_net_\,
            in3 => \N__14113\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__31954\,
            ce => 'H',
            sr => \N__15108\
        );

    \this_vga_signals.M_vcounter_q_2_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14694\,
            in1 => \N__17789\,
            in2 => \_gnd_net_\,
            in3 => \N__14110\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__31954\,
            ce => 'H',
            sr => \N__15108\
        );

    \this_vga_signals.M_vcounter_q_3_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14715\,
            in1 => \N__18913\,
            in2 => \_gnd_net_\,
            in3 => \N__14107\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__31954\,
            ce => 'H',
            sr => \N__15108\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19203\,
            in2 => \_gnd_net_\,
            in3 => \N__14104\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19700\,
            in2 => \_gnd_net_\,
            in3 => \N__14101\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18105\,
            in2 => \_gnd_net_\,
            in3 => \N__14098\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16584\,
            in2 => \_gnd_net_\,
            in3 => \N__14095\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16499\,
            in2 => \_gnd_net_\,
            in3 => \N__14092\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15964\,
            in2 => \_gnd_net_\,
            in3 => \N__14089\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31962\,
            ce => \N__15142\,
            sr => \N__15110\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100011101"
        )
    port map (
            in0 => \N__14939\,
            in1 => \N__15938\,
            in2 => \N__14758\,
            in3 => \N__14891\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15158\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31967\,
            ce => \N__15141\,
            sr => \N__15112\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15159\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31967\,
            ce => \N__15141\,
            sr => \N__15112\
        );

    \this_vga_signals.un5_vaddress_g1_1_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19130\,
            in2 => \_gnd_net_\,
            in3 => \N__18362\,
            lcout => this_vga_signals_un5_vaddress_g1_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14834\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31967\,
            ce => \N__15141\,
            sr => \N__15112\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31967\,
            ce => \N__15141\,
            sr => \N__15112\
        );

    \this_vga_signals.un5_vaddress_g2_3_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111111001"
        )
    port map (
            in0 => \N__17199\,
            in1 => \N__18038\,
            in2 => \N__19231\,
            in3 => \N__19663\,
            lcout => \this_vga_signals.g2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__14940\,
            in1 => \N__14892\,
            in2 => \N__15076\,
            in3 => \N__15965\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011100000000"
        )
    port map (
            in0 => \N__14136\,
            in1 => \N__15064\,
            in2 => \N__14122\,
            in3 => \N__14119\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100111100110"
        )
    port map (
            in0 => \N__17887\,
            in1 => \N__18084\,
            in2 => \N__14176\,
            in3 => \N__14173\,
            lcout => \this_vga_signals.g2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110110010110"
        )
    port map (
            in0 => \N__16138\,
            in1 => \N__16166\,
            in2 => \N__19512\,
            in3 => \N__17883\,
            lcout => \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJHZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_0_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100110010110"
        )
    port map (
            in0 => \N__16167\,
            in1 => \N__19470\,
            in2 => \N__17917\,
            in3 => \N__16139\,
            lcout => \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_31_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110011"
        )
    port map (
            in0 => \N__17679\,
            in1 => \N__14164\,
            in2 => \N__19232\,
            in3 => \N__18372\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_0_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111011100111"
        )
    port map (
            in0 => \N__19664\,
            in1 => \N__19471\,
            in2 => \N__18088\,
            in3 => \N__17200\,
            lcout => \this_vga_signals.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_20_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17673\,
            in1 => \N__15265\,
            in2 => \N__14158\,
            in3 => \N__18232\,
            lcout => \this_vga_signals.N_4_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101001101"
        )
    port map (
            in0 => \N__17177\,
            in1 => \N__19644\,
            in2 => \N__18100\,
            in3 => \N__19507\,
            lcout => \this_vga_signals.g2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICU8TI_6_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011001100011"
        )
    port map (
            in0 => \N__17920\,
            in1 => \N__16280\,
            in2 => \N__18127\,
            in3 => \N__18141\,
            lcout => OPEN,
            ltout => \this_vga_signals.m9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIVKPDR_5_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010100101"
        )
    port map (
            in0 => \N__19703\,
            in1 => \N__18156\,
            in2 => \N__14149\,
            in3 => \N__17921\,
            lcout => \this_vga_signals.N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_3_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110011011101"
        )
    port map (
            in0 => \N__18361\,
            in1 => \N__19202\,
            in2 => \N__19692\,
            in3 => \N__14146\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_30_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18960\,
            in1 => \N__14227\,
            in2 => \N__14221\,
            in3 => \N__17672\,
            lcout => \this_vga_signals.g0_1_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_2_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001100110"
        )
    port map (
            in0 => \N__17919\,
            in1 => \N__14215\,
            in2 => \_gnd_net_\,
            in3 => \N__17178\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_0_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110101011"
        )
    port map (
            in0 => \N__19201\,
            in1 => \N__18360\,
            in2 => \N__14218\,
            in3 => \N__19648\,
            lcout => \this_vga_signals.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__17335\,
            in1 => \N__15077\,
            in2 => \_gnd_net_\,
            in3 => \N__15323\,
            lcout => \this_vga_signals.vaddress_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100010"
        )
    port map (
            in0 => \N__15244\,
            in1 => \N__14209\,
            in2 => \N__19004\,
            in3 => \N__15214\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010001001101"
        )
    port map (
            in0 => \N__18526\,
            in1 => \N__17813\,
            in2 => \N__14203\,
            in3 => \N__14200\,
            lcout => \this_vga_signals.if_i1_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_5_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010000111"
        )
    port map (
            in0 => \N__15324\,
            in1 => \N__17337\,
            in2 => \N__15082\,
            in3 => \N__17220\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_29_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010111000"
        )
    port map (
            in0 => \N__15199\,
            in1 => \N__19241\,
            in2 => \N__14194\,
            in3 => \N__19702\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_2_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_35_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__19242\,
            in1 => \N__14191\,
            in2 => \N__14185\,
            in3 => \N__18397\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__17336\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19472\,
            lcout => \this_vga_signals.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIT8RA8_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__19473\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17680\,
            lcout => \this_vga_signals.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNICEV1S_9_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__14422\,
            in1 => \N__14404\,
            in2 => \N__21001\,
            in3 => \N__14374\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_4_0_wclke_3_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20801\,
            in1 => \N__25732\,
            in2 => \N__23348\,
            in3 => \N__24577\,
            lcout => \this_sprites_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNISLAE4_6_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20998\,
            in2 => \_gnd_net_\,
            in3 => \N__14311\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_0_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110010011001100"
        )
    port map (
            in0 => \N__14716\,
            in1 => \N__16018\,
            in2 => \N__14239\,
            in3 => \N__14531\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31994\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_e_0_RNIR1JA4_1_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110011"
        )
    port map (
            in0 => \N__17434\,
            in1 => \N__16032\,
            in2 => \N__14263\,
            in3 => \N__15994\,
            lcout => \this_vga_signals.M_lcounter_d_0_sqmuxa\,
            ltout => \this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_e_0_1_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000010101010"
        )
    port map (
            in0 => \N__16033\,
            in1 => \N__16017\,
            in2 => \N__14230\,
            in3 => \N__14528\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32002\,
            ce => \N__14717\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_1_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__14566\,
            in1 => \N__14737\,
            in2 => \N__14590\,
            in3 => \N__14530\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32002\,
            ce => \N__14717\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_0_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14529\,
            in1 => \N__14548\,
            in2 => \_gnd_net_\,
            in3 => \N__14565\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32002\,
            ce => \N__14717\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNIOB8H3_0_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14736\,
            in1 => \_gnd_net_\,
            in2 => \N__14719\,
            in3 => \N__14452\,
            lcout => \N_2_0\,
            ltout => \N_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14740\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_pcounter_q_i_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32007\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_RNI5JMN3_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__14505\,
            in1 => \N__14735\,
            in2 => \N__14589\,
            in3 => \N__14564\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_pcounter_q_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNILGGG4_1_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14710\,
            in2 => \N__14593\,
            in3 => \N__14585\,
            lcout => \N_3_0\,
            ltout => \N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14569\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_pcounter_q_i_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32007\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_RNI9FEO2_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__14563\,
            in1 => \N__14547\,
            in2 => \_gnd_net_\,
            in3 => \N__14504\,
            lcout => \this_vga_signals.M_pcounter_q_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_5_0_wclke_3_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__25728\,
            in1 => \N__24568\,
            in2 => \N__23347\,
            in3 => \N__20809\,
            lcout => \this_sprites_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14804\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31950\,
            ce => \N__15145\,
            sr => \N__15107\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__15039\,
            in1 => \N__17342\,
            in2 => \_gnd_net_\,
            in3 => \N__15291\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14833\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31955\,
            ce => \N__15144\,
            sr => \N__15109\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000111"
        )
    port map (
            in0 => \N__14993\,
            in1 => \N__15290\,
            in2 => \N__15060\,
            in3 => \N__14890\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14805\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31955\,
            ce => \N__15144\,
            sr => \N__15109\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14778\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31955\,
            ce => \N__15144\,
            sr => \N__15109\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14909\,
            in1 => \N__14994\,
            in2 => \N__14767\,
            in3 => \N__14967\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15183\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31963\,
            ce => \N__15143\,
            sr => \N__15111\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__14992\,
            in1 => \N__14966\,
            in2 => \_gnd_net_\,
            in3 => \N__14749\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_1_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111101111"
        )
    port map (
            in0 => \N__14911\,
            in1 => \N__14938\,
            in2 => \N__14743\,
            in3 => \N__15937\,
            lcout => OPEN,
            ltout => \this_vga_signals.SUM_2_i_1_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__15007\,
            in1 => \N__14863\,
            in2 => \N__15001\,
            in3 => \N__14947\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__15935\,
            in1 => \N__14991\,
            in2 => \N__14941\,
            in3 => \N__14886\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14971\,
            in3 => \N__14965\,
            lcout => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15182\,
            lcout => \this_vga_signals.M_vcounter_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31963\,
            ce => \N__15143\,
            sr => \N__15111\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001111111"
        )
    port map (
            in0 => \N__14937\,
            in1 => \N__14910\,
            in2 => \N__14893\,
            in3 => \N__15936\,
            lcout => \this_vga_signals.SUM_2_i_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m2_1_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010011000011"
        )
    port map (
            in0 => \N__17171\,
            in1 => \N__16136\,
            in2 => \N__16178\,
            in3 => \N__17901\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI87FSD_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17170\,
            in2 => \N__14857\,
            in3 => \N__14848\,
            lcout => \this_vga_signals.d_N_3_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010100101"
        )
    port map (
            in0 => \N__17172\,
            in1 => \N__16137\,
            in2 => \N__16179\,
            in3 => \N__17902\,
            lcout => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i,
            ltout => \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \m18x_N_3L3_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111001000"
        )
    port map (
            in0 => \N__16950\,
            in1 => \N__17593\,
            in2 => \N__14842\,
            in3 => \N__18267\,
            lcout => \m18x_N_3LZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_15_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17174\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18116\,
            lcout => \this_vga_signals.N_5_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIM43JE1_5_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__15208\,
            in1 => \N__17467\,
            in2 => \N__16069\,
            in3 => \N__17594\,
            lcout => \this_vga_signals.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_1_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__17344\,
            in1 => \N__15066\,
            in2 => \_gnd_net_\,
            in3 => \N__15310\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_1_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001011010"
        )
    port map (
            in0 => \N__17903\,
            in1 => \_gnd_net_\,
            in2 => \N__15202\,
            in3 => \N__17173\,
            lcout => \this_vga_signals.g2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_37_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__15996\,
            in1 => \N__16442\,
            in2 => \N__18123\,
            in3 => \N__16539\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15187\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31972\,
            ce => \N__15139\,
            sr => \N__15113\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15166\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31972\,
            ce => \N__15139\,
            sr => \N__15113\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__16538\,
            in1 => \N__15065\,
            in2 => \N__16468\,
            in3 => \N__15995\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_1\,
            ltout => \this_vga_signals.if_m8_0_a3_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17341\,
            in2 => \N__15010\,
            in3 => \N__15309\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001110"
        )
    port map (
            in0 => \N__16134\,
            in1 => \N__16168\,
            in2 => \N__15328\,
            in3 => \N__17175\,
            lcout => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17340\,
            in2 => \_gnd_net_\,
            in3 => \N__15308\,
            lcout => \this_vga_signals.vaddress_5\,
            ltout => \this_vga_signals.vaddress_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001010"
        )
    port map (
            in0 => \N__16135\,
            in1 => \N__17176\,
            in2 => \N__15268\,
            in3 => \N__17918\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_2_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18996\,
            in1 => \N__15264\,
            in2 => \N__19257\,
            in3 => \N__17678\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_26_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101111111"
        )
    port map (
            in0 => \N__17812\,
            in1 => \N__15253\,
            in2 => \N__15247\,
            in3 => \N__18228\,
            lcout => \this_vga_signals.g1_0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIB3A8M_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__15238\,
            in1 => \N__16347\,
            in2 => \N__19360\,
            in3 => \N__18391\,
            lcout => \this_vga_signals.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x2_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15229\,
            in1 => \N__16288\,
            in2 => \_gnd_net_\,
            in3 => \N__18229\,
            lcout => \this_vga_signals.N_5_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_2_x1_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__16310\,
            in1 => \N__19237\,
            in2 => \N__19013\,
            in3 => \N__17676\,
            lcout => \this_vga_signals.g0_2_0_2_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_2_x0_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17677\,
            in1 => \N__18995\,
            in2 => \N__19255\,
            in3 => \N__16309\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_2_0_2_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_2_ns_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15481\,
            in2 => \N__15475\,
            in3 => \N__18390\,
            lcout => \this_vga_signals.g0_2_0_2\,
            ltout => \this_vga_signals.g0_2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111110111"
        )
    port map (
            in0 => \N__17811\,
            in1 => \N__16224\,
            in2 => \N__15472\,
            in3 => \N__17563\,
            lcout => \this_vga_signals.g1_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15469\,
            in1 => \N__15451\,
            in2 => \_gnd_net_\,
            in3 => \N__27822\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15436\,
            in1 => \N__15421\,
            in2 => \_gnd_net_\,
            in3 => \N__27821\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_wclke_3_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__25723\,
            in1 => \N__24576\,
            in2 => \N__23350\,
            in3 => \N__20800\,
            lcout => \this_sprites_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101010011"
        )
    port map (
            in0 => \N__16869\,
            in1 => \N__16803\,
            in2 => \N__16673\,
            in3 => \N__16739\,
            lcout => \this_vga_ramdac.m6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__15379\,
            in1 => \N__27459\,
            in2 => \N__15369\,
            in3 => \N__15861\,
            lcout => \this_vga_ramdac.N_2871_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.G_384_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15799\,
            in1 => \N__15816\,
            in2 => \_gnd_net_\,
            in3 => \N__15807\,
            lcout => \G_384\,
            ltout => \G_384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__15339\,
            in1 => \N__16594\,
            in2 => \N__15352\,
            in3 => \N__27461\,
            lcout => \this_vga_ramdac.N_2872_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__16031\,
            in1 => \N__16016\,
            in2 => \_gnd_net_\,
            in3 => \N__16000\,
            lcout => \this_vga_signals.line_clk_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__16879\,
            in1 => \N__27460\,
            in2 => \N__15834\,
            in3 => \N__15862\,
            lcout => \this_vga_ramdac.N_2873_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15817\,
            in2 => \_gnd_net_\,
            in3 => \N__15808\,
            lcout => \M_this_vga_signals_pixel_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIBSKN5_1_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15659\,
            in1 => \N__15513\,
            in2 => \_gnd_net_\,
            in3 => \N__21972\,
            lcout => \this_ppu.un1_M_vaddress_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_6_0_wclke_3_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__25716\,
            in1 => \N__24567\,
            in2 => \N__23349\,
            in3 => \N__20808\,
            lcout => \this_sprites_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_0_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22008\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15648\,
            lcout => \M_this_ppu_vram_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32016\,
            ce => 'H',
            sr => \N__21466\
        );

    \this_ppu.M_vaddress_q_1_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__22009\,
            in1 => \N__15647\,
            in2 => \_gnd_net_\,
            in3 => \N__15505\,
            lcout => \M_this_ppu_sprites_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32016\,
            ce => 'H',
            sr => \N__21466\
        );

    \this_ppu.M_vaddress_q_2_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__15655\,
            in1 => \N__15512\,
            in2 => \N__20352\,
            in3 => \N__22023\,
            lcout => \M_this_ppu_sprites_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32032\,
            ce => 'H',
            sr => \N__21492\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGE761_6_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__18104\,
            in1 => \N__19693\,
            in2 => \_gnd_net_\,
            in3 => \N__19513\,
            lcout => \this_vga_signals.vaddress_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_2_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17343\,
            lcout => \this_vga_signals.vaddress_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000001111"
        )
    port map (
            in0 => \N__16183\,
            in1 => \N__17235\,
            in2 => \N__16141\,
            in3 => \N__17915\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110100101"
        )
    port map (
            in0 => \N__19707\,
            in1 => \N__16087\,
            in2 => \N__16078\,
            in3 => \N__17461\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNINM635_5_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011110110010"
        )
    port map (
            in0 => \N__19141\,
            in1 => \N__19752\,
            in2 => \N__19706\,
            in3 => \N__16075\,
            lcout => \this_vga_signals.i2_mux\,
            ltout => \this_vga_signals.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5BS7N_5_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101100110"
        )
    port map (
            in0 => \N__19675\,
            in1 => \N__17836\,
            in2 => \N__16060\,
            in3 => \N__17465\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNI5BS7NZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m4_0_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__18972\,
            in1 => \N__19525\,
            in2 => \_gnd_net_\,
            in3 => \N__18330\,
            lcout => \this_vga_signals.if_i2_mux\,
            ltout => \this_vga_signals.if_i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_17_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100111111001"
        )
    port map (
            in0 => \N__17092\,
            in1 => \N__19680\,
            in2 => \N__16057\,
            in3 => \N__17350\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_7_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__19138\,
            in1 => \N__17650\,
            in2 => \_gnd_net_\,
            in3 => \N__18328\,
            lcout => \this_vga_signals.g1_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001001010101"
        )
    port map (
            in0 => \N__16050\,
            in1 => \N__17234\,
            in2 => \N__17508\,
            in3 => \N__17916\,
            lcout => \this_vga_signals.g1_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_23_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__19139\,
            in1 => \N__19671\,
            in2 => \_gnd_net_\,
            in3 => \N__19751\,
            lcout => \this_vga_signals.if_N_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110011011101"
        )
    port map (
            in0 => \N__18329\,
            in1 => \N__19140\,
            in2 => \N__19704\,
            in3 => \N__16246\,
            lcout => \this_vga_signals.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIVRE454_5_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16240\,
            in1 => \N__16234\,
            in2 => \N__16228\,
            in3 => \N__16971\,
            lcout => \this_vga_signals.i14_mux_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x0_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000110110"
        )
    port map (
            in0 => \N__16311\,
            in1 => \N__19000\,
            in2 => \N__18389\,
            in3 => \N__19523\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_axb1_0_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_ns_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__17658\,
            in1 => \_gnd_net_\,
            in2 => \N__16210\,
            in3 => \N__16204\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_0\,
            ltout => \this_vga_signals.mult1_un68_sum_axb1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_6_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111110111"
        )
    port map (
            in0 => \N__17804\,
            in1 => \N__16252\,
            in2 => \N__16207\,
            in3 => \N__17518\,
            lcout => \this_vga_signals.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000011111001"
        )
    port map (
            in0 => \N__19521\,
            in1 => \N__18964\,
            in2 => \N__16282\,
            in3 => \N__17589\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_4_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18965\,
            in1 => \N__19522\,
            in2 => \_gnd_net_\,
            in3 => \N__17657\,
            lcout => \this_vga_signals.g0_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x1_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001001011"
        )
    port map (
            in0 => \N__19524\,
            in1 => \N__18356\,
            in2 => \N__19014\,
            in3 => \N__16312\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_0_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100101100110"
        )
    port map (
            in0 => \N__16384\,
            in1 => \N__16375\,
            in2 => \N__19005\,
            in3 => \N__18421\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHM0ARA_5_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100111000011"
        )
    port map (
            in0 => \N__16366\,
            in1 => \N__16360\,
            in2 => \N__17689\,
            in3 => \N__16354\,
            lcout => \this_vga_signals.i13_mux_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI3HO5K_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110011"
        )
    port map (
            in0 => \N__17647\,
            in1 => \N__16348\,
            in2 => \N__19527\,
            in3 => \N__18355\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_N_4L5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5E1_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100110110"
        )
    port map (
            in0 => \N__19356\,
            in1 => \N__16327\,
            in2 => \N__16318\,
            in3 => \N__17649\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5EZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIAO8TO2_2_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101101001101"
        )
    port map (
            in0 => \N__17805\,
            in1 => \N__19010\,
            in2 => \N__16315\,
            in3 => \N__18230\,
            lcout => \this_vga_signals.m21_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_520_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110010011001"
        )
    port map (
            in0 => \N__16308\,
            in1 => \N__17646\,
            in2 => \N__19526\,
            in3 => \N__18327\,
            lcout => if_generate_plus_mult1_un68_sum_axb1_520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_1_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__17648\,
            in1 => \_gnd_net_\,
            in2 => \N__19253\,
            in3 => \N__19009\,
            lcout => \this_vga_signals.g0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18354\,
            in1 => \N__16281\,
            in2 => \_gnd_net_\,
            in3 => \N__16261\,
            lcout => \this_vga_signals.mult1_un61_sum_c3\,
            ltout => \this_vga_signals.mult1_un61_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_7_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19221\,
            in1 => \N__19008\,
            in2 => \N__16255\,
            in3 => \N__18264\,
            lcout => \this_vga_signals.g0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011010000"
        )
    port map (
            in0 => \N__17403\,
            in1 => \N__16467\,
            in2 => \N__16402\,
            in3 => \N__16560\,
            lcout => \this_ppu.line_clk.M_last_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31973\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010101010"
        )
    port map (
            in0 => \N__16972\,
            in1 => \N__16957\,
            in2 => \N__16939\,
            in3 => \N__17595\,
            lcout => \this_vga_signals.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIKBOI74_4_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16924\,
            in1 => \N__18268\,
            in2 => \N__19258\,
            in3 => \N__16918\,
            lcout => \this_vga_signals.m21_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__16912\,
            in1 => \N__16900\,
            in2 => \N__23203\,
            in3 => \N__19312\,
            lcout => \M_this_ppu_vram_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIMRAD5_5_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20028\,
            lcout => \this_ppu.M_last_q_RNIMRAD5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110100010111"
        )
    port map (
            in0 => \N__16644\,
            in1 => \N__16743\,
            in2 => \N__16804\,
            in3 => \N__16855\,
            lcout => \this_vga_ramdac.m16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011101"
        )
    port map (
            in0 => \N__16854\,
            in1 => \N__16791\,
            in2 => \N__16752\,
            in3 => \N__16645\,
            lcout => \this_vga_ramdac.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIUNVB4_7_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101100000000"
        )
    port map (
            in0 => \N__16586\,
            in1 => \N__17404\,
            in2 => \N__16503\,
            in3 => \N__16395\,
            lcout => \M_this_vga_signals_line_clk_0\,
            ltout => \M_this_vga_signals_line_clk_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIMRAD5_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18750\,
            in1 => \N__20608\,
            in2 => \N__17086\,
            in3 => \N__20098\,
            lcout => \this_ppu.M_state_d_0_sqmuxa\,
            ltout => \this_ppu.M_state_d_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_1_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__18457\,
            in1 => \N__20184\,
            in2 => \N__17083\,
            in3 => \N__27482\,
            lcout => \this_ppu.M_count_qZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31988\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_0_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__27481\,
            in1 => \N__20100\,
            in2 => \_gnd_net_\,
            in3 => \N__21994\,
            lcout => \this_ppu.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31988\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17080\,
            in1 => \N__17065\,
            in2 => \_gnd_net_\,
            in3 => \N__27820\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIMRAD5_4_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20107\,
            in2 => \_gnd_net_\,
            in3 => \N__20023\,
            lcout => \this_ppu.M_last_q_RNIMRAD5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_0_c_RNO_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20106\,
            in2 => \_gnd_net_\,
            in3 => \N__20022\,
            lcout => \this_ppu.un1_M_count_q_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17053\,
            in1 => \N__17041\,
            in2 => \_gnd_net_\,
            in3 => \N__27800\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIQKTIG_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001010"
        )
    port map (
            in0 => \N__22001\,
            in1 => \N__21641\,
            in2 => \N__17028\,
            in3 => \N__27480\,
            lcout => \this_ppu.M_last_q_RNIQKTIG\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_1_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001011111"
        )
    port map (
            in0 => \N__19217\,
            in1 => \_gnd_net_\,
            in2 => \N__19714\,
            in3 => \N__18103\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17509\,
            in1 => \N__17386\,
            in2 => \N__17482\,
            in3 => \N__17236\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18527\,
            in2 => \_gnd_net_\,
            in3 => \N__18579\,
            lcout => \this_vga_signals.M_vcounter_d7lt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111000011"
        )
    port map (
            in0 => \N__17479\,
            in1 => \N__17473\,
            in2 => \N__19705\,
            in3 => \N__17466\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIJPU72_2_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__17801\,
            in1 => \N__17440\,
            in2 => \N__19006\,
            in3 => \N__19517\,
            lcout => \this_vga_signals.M_vcounter_d7lt9_1\,
            ltout => \this_vga_signals.M_vcounter_d7lt9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIAEPU2_6_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110101"
        )
    port map (
            in0 => \N__19676\,
            in1 => \_gnd_net_\,
            in2 => \N__17407\,
            in3 => \N__18102\,
            lcout => \this_vga_signals.un4_lvisibility_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_1_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19518\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17338\,
            lcout => \this_vga_signals.vaddress_1_5\,
            ltout => \this_vga_signals.vaddress_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_18_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__17382\,
            in1 => \N__17365\,
            in2 => \N__17353\,
            in3 => \N__17233\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__19519\,
            in1 => \N__18101\,
            in2 => \_gnd_net_\,
            in3 => \N__17339\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_4_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000001111"
        )
    port map (
            in0 => \N__17242\,
            in1 => \N__17232\,
            in2 => \N__17095\,
            in3 => \N__17929\,
            lcout => \this_vga_signals.g1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNITP439_0_2_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101001100101"
        )
    port map (
            in0 => \N__18371\,
            in1 => \N__18978\,
            in2 => \N__19249\,
            in3 => \N__17803\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_RNITP439_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIFPMH71_2_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18834\,
            in2 => \N__17692\,
            in3 => \N__17551\,
            lcout => \this_vga_signals.m16_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__17674\,
            in1 => \N__18368\,
            in2 => \N__19247\,
            in3 => \N__17599\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18976\,
            in2 => \N__17566\,
            in3 => \N__18262\,
            lcout => \this_vga_signals.g0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNITP439_2_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011000111001"
        )
    port map (
            in0 => \N__18977\,
            in1 => \N__17802\,
            in2 => \N__19248\,
            in3 => \N__18369\,
            lcout => \this_vga_signals.M_vcounter_q_RNITP439Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18370\,
            in1 => \N__18263\,
            in2 => \N__18842\,
            in3 => \N__18217\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_0_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__17545\,
            in1 => \N__17536\,
            in2 => \N__17530\,
            in3 => \N__18218\,
            lcout => \this_vga_signals.g0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18835\,
            in1 => \N__18265\,
            in2 => \_gnd_net_\,
            in3 => \N__18219\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_1_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100110011100"
        )
    port map (
            in0 => \N__19012\,
            in1 => \N__19216\,
            in2 => \N__17512\,
            in3 => \N__17806\,
            lcout => \this_vga_signals.mult1_un82_sum_c3_0_N_4L5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_3_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110010011001"
        )
    port map (
            in0 => \N__18439\,
            in1 => \N__18427\,
            in2 => \N__19254\,
            in3 => \N__18393\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_21_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110111011010"
        )
    port map (
            in0 => \N__18420\,
            in1 => \N__19011\,
            in2 => \N__18409\,
            in3 => \N__18221\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__18406\,
            in1 => \N__17807\,
            in2 => \N__18400\,
            in3 => \N__18169\,
            lcout => \this_vga_signals.N_5_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18392\,
            in1 => \N__18266\,
            in2 => \N__18843\,
            in3 => \N__18220\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18805\,
            in2 => \N__18178\,
            in3 => \N__18175\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011000011"
        )
    port map (
            in0 => \N__18163\,
            in1 => \N__18145\,
            in2 => \N__18130\,
            in3 => \N__17944\,
            lcout => \this_vga_signals.g1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI1RPOO2_1_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000101000"
        )
    port map (
            in0 => \N__17824\,
            in1 => \N__17817\,
            in2 => \N__18548\,
            in3 => \N__17722\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_25_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5P1Q0M_4_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101011001"
        )
    port map (
            in0 => \N__17713\,
            in1 => \N__17707\,
            in2 => \N__17695\,
            in3 => \N__18625\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIGBAMTL1_9_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__21000\,
            in1 => \N__18619\,
            in2 => \N__18610\,
            in3 => \N__18481\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__18586\,
            in1 => \N__18844\,
            in2 => \N__18549\,
            in3 => \N__18556\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_N_4L5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_m2_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18544\,
            in2 => \N__18490\,
            in3 => \N__18487\,
            lcout => \this_vga_signals.mult1_un82_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_2_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27450\,
            in1 => \N__21990\,
            in2 => \N__20188\,
            in3 => \N__18448\,
            lcout => \this_ppu.M_count_qZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18475\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_0_c_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18463\,
            in2 => \N__19812\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \this_ppu.un1_M_count_q_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_1_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18721\,
            in2 => \N__19851\,
            in3 => \N__18451\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_0\,
            carryout => \this_ppu.un1_M_count_q_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18637\,
            in2 => \N__19834\,
            in3 => \N__18442\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_3_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20272\,
            in2 => \N__20259\,
            in3 => \N__18670\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_2\,
            carryout => \this_ppu.un1_M_count_q_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_4_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18667\,
            in2 => \N__20242\,
            in3 => \N__18661\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_3\,
            carryout => \this_ppu.un1_M_count_q_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_5_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18643\,
            in2 => \N__20122\,
            in3 => \N__18658\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_4\,
            carryout => \this_ppu.un1_M_count_q_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_6_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18655\,
            in2 => \N__20227\,
            in3 => \N__18649\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_5\,
            carryout => \this_ppu.un1_M_count_q_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_7_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101010100"
        )
    port map (
            in0 => \N__20159\,
            in1 => \N__19990\,
            in2 => \N__22011\,
            in3 => \N__18646\,
            lcout => \this_ppu.M_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31981\,
            ce => 'H',
            sr => \N__32392\
        );

    \this_ppu.line_clk.M_last_q_RNIMRAD5_1_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20025\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20094\,
            lcout => \this_ppu.M_last_q_RNIMRAD5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIMRAD5_0_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20092\,
            in2 => \_gnd_net_\,
            in3 => \N__20024\,
            lcout => \this_ppu.M_last_q_RNIMRAD5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_4_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27452\,
            in1 => \N__21988\,
            in2 => \N__20177\,
            in3 => \N__18631\,
            lcout => \this_ppu.M_count_qZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31989\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_0_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__19813\,
            in1 => \N__20093\,
            in2 => \_gnd_net_\,
            in3 => \N__20026\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_count_q_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_0_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27451\,
            in1 => \N__20160\,
            in2 => \N__18760\,
            in3 => \N__21989\,
            lcout => \this_ppu.M_count_qZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31989\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_6_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__21987\,
            in1 => \N__27453\,
            in2 => \N__20175\,
            in3 => \N__18757\,
            lcout => \this_ppu.M_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31989\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIMMU35_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__18751\,
            in1 => \N__20601\,
            in2 => \_gnd_net_\,
            in3 => \N__18730\,
            lcout => \this_ppu.N_82_i\,
            ltout => \this_ppu.N_82_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIMRAD5_3_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18724\,
            in3 => \N__20091\,
            lcout => \this_ppu.M_last_q_RNIMRAD5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_3_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20357\,
            in1 => \N__20482\,
            in2 => \_gnd_net_\,
            in3 => \N__20304\,
            lcout => \M_this_ppu_map_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32008\,
            ce => 'H',
            sr => \N__21467\
        );

    \this_ppu.M_vaddress_q_4_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__20525\,
            in1 => \N__20483\,
            in2 => \N__20356\,
            in3 => \N__20305\,
            lcout => \M_this_ppu_map_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32017\,
            ce => 'H',
            sr => \N__21493\
        );

    \this_reset_cond.M_stage_q_4_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__28471\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18715\,
            lcout => \this_reset_cond.M_stage_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__28470\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20710\,
            lcout => \this_reset_cond.M_stage_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27823\,
            in1 => \N__18709\,
            in2 => \_gnd_net_\,
            in3 => \N__18691\,
            lcout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27824\,
            in1 => \N__19789\,
            in2 => \_gnd_net_\,
            in3 => \N__19768\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_13_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19753\,
            in1 => \N__19710\,
            in2 => \_gnd_net_\,
            in3 => \N__19528\,
            lcout => \this_vga_signals.if_N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_5_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__28481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19333\,
            lcout => \this_reset_cond.M_stage_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31951\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__23185\,
            in1 => \N__19324\,
            in2 => \N__29672\,
            in3 => \N__19318\,
            lcout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_6_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__19300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28482\,
            lcout => \this_reset_cond.M_stage_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31951\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27825\,
            in1 => \N__19294\,
            in2 => \_gnd_net_\,
            in3 => \N__19279\,
            lcout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011011101"
        )
    port map (
            in0 => \N__19256\,
            in1 => \N__19007\,
            in2 => \_gnd_net_\,
            in3 => \N__18830\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27762\,
            in1 => \N__18799\,
            in2 => \_gnd_net_\,
            in3 => \N__18781\,
            lcout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27826\,
            in1 => \N__19978\,
            in2 => \_gnd_net_\,
            in3 => \N__19960\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__29645\,
            in1 => \N__23161\,
            in2 => \N__19945\,
            in3 => \N__19942\,
            lcout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__23198\,
            in1 => \N__20668\,
            in2 => \N__29673\,
            in3 => \N__19936\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__23192\,
            in1 => \N__19927\,
            in2 => \N__19915\,
            in3 => \N__19861\,
            lcout => \M_this_ppu_vram_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19897\,
            in1 => \N__19882\,
            in2 => \_gnd_net_\,
            in3 => \N__27819\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_1_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20203\,
            in1 => \N__20209\,
            in2 => \_gnd_net_\,
            in3 => \N__20097\,
            lcout => OPEN,
            ltout => \this_ppu.N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_1_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__20613\,
            in1 => \N__20577\,
            in2 => \N__19855\,
            in3 => \N__32436\,
            lcout => \this_ppu.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNI230G_0_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19852\,
            in1 => \N__19833\,
            in2 => \N__20260\,
            in3 => \N__19808\,
            lcout => \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI05C9_1_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20576\,
            lcout => \this_ppu.M_state_q_i_1\,
            ltout => \this_ppu.M_state_q_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIMRAD5_2_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20275\,
            in3 => \N__20027\,
            lcout => \this_ppu.M_last_q_RNIMRAD5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_3_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27496\,
            in1 => \N__22010\,
            in2 => \N__20176\,
            in3 => \N__20266\,
            lcout => \this_ppu.M_count_qZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIIJ0G_7_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20238\,
            in1 => \N__20220\,
            in2 => \N__20041\,
            in3 => \N__20118\,
            lcout => \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4\,
            ltout => \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIJVOI1_0_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20202\,
            in1 => \N__20617\,
            in2 => \N__20191\,
            in3 => \N__20095\,
            lcout => \this_ppu.M_state_d_0_sqmuxa_1\,
            ltout => \this_ppu.M_state_d_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_5_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27495\,
            in1 => \N__22022\,
            in2 => \N__20131\,
            in3 => \N__20128\,
            lcout => \this_ppu.M_count_qZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31982\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_7_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20096\,
            in1 => \N__20040\,
            in2 => \_gnd_net_\,
            in3 => \N__20029\,
            lcout => \this_ppu.un1_M_count_q_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28467\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__28468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19984\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__28469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20716\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__25789\,
            in1 => \N__27554\,
            in2 => \N__27002\,
            in3 => \N__32830\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31956\,
            ce => 'H',
            sr => \N__32390\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27818\,
            in1 => \N__20704\,
            in2 => \_gnd_net_\,
            in3 => \N__20686\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__20662\,
            in1 => \N__20653\,
            in2 => \N__23199\,
            in3 => \N__20641\,
            lcout => \M_this_ppu_vram_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIV8OI_1_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20612\,
            in2 => \_gnd_net_\,
            in3 => \N__20578\,
            lcout => \M_this_ppu_vram_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_7_0_wclke_3_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25708\,
            in1 => \N__24561\,
            in2 => \N__23319\,
            in3 => \N__20788\,
            lcout => \this_sprites_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_m_2_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30306\,
            in2 => \_gnd_net_\,
            in3 => \N__30597\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNI25476_4_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20529\,
            in1 => \N__20493\,
            in2 => \N__20364\,
            in3 => \N__20303\,
            lcout => \this_ppu.un1_M_vaddress_q_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_6_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__21551\,
            in1 => \N__21522\,
            in2 => \_gnd_net_\,
            in3 => \N__23885\,
            lcout => \this_ppu.M_vaddress_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32009\,
            ce => 'H',
            sr => \N__21503\
        );

    \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23712\,
            in2 => \_gnd_net_\,
            in3 => \N__24469\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20878\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_en_0_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27924\,
            in1 => \N__27207\,
            in2 => \_gnd_net_\,
            in3 => \N__32638\,
            lcout => \M_this_sprites_ram_write_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI2S2S_13_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27925\,
            in1 => \N__27208\,
            in2 => \N__31327\,
            in3 => \N__28017\,
            lcout => \M_this_state_q_RNI2S2SZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_fast_15_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__27216\,
            in1 => \N__27169\,
            in2 => \N__27096\,
            in3 => \N__27052\,
            lcout => \M_this_state_q_fastZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31949\,
            ce => 'H',
            sr => \N__32388\
        );

    \M_this_state_q_14_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001010"
        )
    port map (
            in0 => \N__27226\,
            in1 => \N__28528\,
            in2 => \N__32851\,
            in3 => \N__25768\,
            lcout => \M_this_state_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31949\,
            ce => 'H',
            sr => \N__32388\
        );

    \this_vga_signals.M_this_state_q_tr43_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__27215\,
            in1 => \N__27168\,
            in2 => \N__27097\,
            in3 => \N__27051\,
            lcout => \this_vga_signals.M_this_state_q_ns_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_wclke_3_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__25725\,
            in1 => \N__24562\,
            in2 => \N__23339\,
            in3 => \N__20769\,
            lcout => \this_sprites_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_wclke_3_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20770\,
            in1 => \N__23323\,
            in2 => \N__24575\,
            in3 => \N__25726\,
            lcout => \this_sprites_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__25727\,
            in1 => \N__24566\,
            in2 => \N__23340\,
            in3 => \N__20771\,
            lcout => \this_sprites_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_0_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__22653\,
            in1 => \N__33818\,
            in2 => \N__33340\,
            in3 => \N__21104\,
            lcout => \M_this_sprites_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_1_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__21105\,
            in1 => \N__33982\,
            in2 => \N__33642\,
            in3 => \N__22654\,
            lcout => \M_this_sprites_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010101"
        )
    port map (
            in0 => \N__27945\,
            in1 => \N__25392\,
            in2 => \N__27227\,
            in3 => \N__32786\,
            lcout => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\,
            ltout => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_2_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__33512\,
            in1 => \N__34212\,
            in2 => \N__21205\,
            in3 => \N__22655\,
            lcout => \M_this_sprites_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__24594\,
            in1 => \N__32785\,
            in2 => \N__24042\,
            in3 => \N__30598\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31961\,
            ce => 'H',
            sr => \N__32389\
        );

    \M_this_state_q_12_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100010000"
        )
    port map (
            in0 => \N__32784\,
            in1 => \N__28524\,
            in2 => \N__23995\,
            in3 => \N__27994\,
            lcout => \M_this_state_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31961\,
            ce => 'H',
            sr => \N__32389\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_3_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__34347\,
            in1 => \N__22662\,
            in2 => \N__33427\,
            in3 => \N__21109\,
            lcout => \M_this_sprites_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNICRTO5_9_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20991\,
            in2 => \_gnd_net_\,
            in3 => \N__20920\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_0_5_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__27003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26856\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_0_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__22252\,
            in1 => \N__22219\,
            in2 => \_gnd_net_\,
            in3 => \N__22027\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31987\,
            ce => 'H',
            sr => \N__25036\
        );

    \this_ppu.M_haddress_q_1_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110001111000"
        )
    port map (
            in0 => \N__22026\,
            in1 => \N__22251\,
            in2 => \N__22066\,
            in3 => \N__22220\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31987\,
            ce => 'H',
            sr => \N__25036\
        );

    \this_ppu.M_vaddress_q_5_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21521\,
            in2 => \_gnd_net_\,
            in3 => \N__21547\,
            lcout => \M_this_ppu_map_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31993\,
            ce => 'H',
            sr => \N__21505\
        );

    \this_ppu.M_vaddress_q_7_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__21445\,
            in1 => \N__23886\,
            in2 => \N__21555\,
            in3 => \N__21523\,
            lcout => \this_ppu.M_vaddress_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32001\,
            ce => 'H',
            sr => \N__21504\
        );

    \this_ppu.M_vaddress_q_RNI1DAA_7_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21444\,
            in2 => \_gnd_net_\,
            in3 => \N__23881\,
            lcout => \M_this_ppu_map_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__24016\,
            in1 => \N__28198\,
            in2 => \N__26877\,
            in3 => \N__32790\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31946\,
            ce => 'H',
            sr => \N__32391\
        );

    \this_vga_signals.M_this_sprites_address_q_m_1_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25501\,
            in2 => \_gnd_net_\,
            in3 => \N__24474\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32431\,
            lcout => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__22855\,
            in1 => \N__24473\,
            in2 => \N__34213\,
            in3 => \N__32777\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_8_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23002\,
            in2 => \_gnd_net_\,
            in3 => \N__28161\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_8_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__21673\,
            in1 => \N__24151\,
            in2 => \N__21664\,
            in3 => \N__22978\,
            lcout => \M_this_sprites_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31952\,
            ce => 'H',
            sr => \N__27289\
        );

    \this_vga_signals.un23_i_a2_x1_0_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31202\,
            in1 => \N__29616\,
            in2 => \N__31323\,
            in3 => \N__25382\,
            lcout => OPEN,
            ltout => \this_vga_signals.un23_i_a2_x1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un23_i_a2_ns_0_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21655\,
            in3 => \N__21685\,
            lcout => dma_axb0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dma_ac0_5_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__31252\,
            in1 => \N__21592\,
            in2 => \N__25447\,
            in3 => \N__21607\,
            lcout => \dma_ac0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un23_i_a2_4_2_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29617\,
            in1 => \N__30784\,
            in2 => \N__27607\,
            in3 => \N__30609\,
            lcout => this_vga_signals_un23_i_a2_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un23_i_a2_1_3_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__25383\,
            in1 => \_gnd_net_\,
            in2 => \N__28040\,
            in3 => \N__32924\,
            lcout => this_vga_signals_un23_i_a2_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un23_i_a2_3_2_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31316\,
            in1 => \N__27206\,
            in2 => \N__27946\,
            in3 => \N__28027\,
            lcout => OPEN,
            ltout => \this_vga_signals_un23_i_a2_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dma_c3_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__21601\,
            in1 => \N__24061\,
            in2 => \N__21595\,
            in3 => \N__21585\,
            lcout => dma_c3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNITS9I4_7_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101110111"
        )
    port map (
            in0 => \N__21679\,
            in1 => \N__21586\,
            in2 => \N__24076\,
            in3 => \N__25445\,
            lcout => OPEN,
            ltout => \M_this_state_q_RNITS9I4Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIV6UJ7_8_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__21910\,
            in1 => \N__25446\,
            in2 => \N__21901\,
            in3 => \N__22393\,
            lcout => dma_ac0_5_i,
            ltout => \dma_ac0_5_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIV6UJ7_0_8_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21874\,
            in3 => \_gnd_net_\,
            lcout => dma_ac0_5_i_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_3_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__24052\,
            in1 => \N__26399\,
            in2 => \N__22387\,
            in3 => \N__32788\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31964\,
            ce => 'H',
            sr => \N__32382\
        );

    \this_vga_signals.un23_i_a2_4_0_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24403\,
            in1 => \N__30578\,
            in2 => \N__26425\,
            in3 => \N__25461\,
            lcout => \this_vga_signals.un23_i_a2_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__24012\,
            in1 => \N__26873\,
            in2 => \N__24467\,
            in3 => \N__32787\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31964\,
            ce => 'H',
            sr => \N__32382\
        );

    \M_this_state_q_RNI6Q0S_7_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29620\,
            in1 => \N__27621\,
            in2 => \N__30648\,
            in3 => \N__30847\,
            lcout => \M_this_state_q_RNI6Q0SZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__32774\,
            in1 => \N__23009\,
            in2 => \N__33981\,
            in3 => \N__24431\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__22715\,
            in1 => \N__34333\,
            in2 => \N__24466\,
            in3 => \N__32776\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__32775\,
            in1 => \N__23271\,
            in2 => \N__33538\,
            in3 => \N__24435\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_0_3_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__27004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26863\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_13_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23272\,
            in2 => \_gnd_net_\,
            in3 => \N__28211\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_10_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__22378\,
            in1 => \N__24175\,
            in2 => \N__22408\,
            in3 => \N__22681\,
            lcout => \M_this_sprites_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31976\,
            ce => 'H',
            sr => \N__27284\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__25663\,
            in1 => \N__24455\,
            in2 => \N__33641\,
            in3 => \N__32826\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_4_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24454\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26165\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNI21NK5_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27494\,
            in2 => \_gnd_net_\,
            in3 => \N__22024\,
            lcout => \this_ppu.M_last_q_RNI21NK5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIEKA06_1_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__22262\,
            in1 => \N__22224\,
            in2 => \N__22076\,
            in3 => \N__22025\,
            lcout => \this_ppu.un1_M_haddress_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_2_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23428\,
            in2 => \_gnd_net_\,
            in3 => \N__23976\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32018\,
            ce => 'H',
            sr => \N__25030\
        );

    \this_vga_signals.M_this_sprites_address_q_m_9_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28160\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_3_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28258\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24480\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_1_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__25474\,
            in1 => \N__24170\,
            in2 => \N__22456\,
            in3 => \N__22630\,
            lcout => \M_this_sprites_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31953\,
            ce => 'H',
            sr => \N__27291\
        );

    \M_this_sprites_address_q_9_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__24171\,
            in1 => \N__22447\,
            in2 => \N__22441\,
            in3 => \N__22831\,
            lcout => \M_this_sprites_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31953\,
            ce => 'H',
            sr => \N__27291\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__22507\,
            in1 => \N__28170\,
            in2 => \N__34220\,
            in3 => \N__32639\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_2_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__22426\,
            in1 => \N__24142\,
            in2 => \N__22429\,
            in3 => \N__22486\,
            lcout => \M_this_sprites_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31957\,
            ce => 'H',
            sr => \N__27290\
        );

    \this_vga_signals.M_this_sprites_address_q_m_2_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24465\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_3_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__24143\,
            in1 => \N__28093\,
            in2 => \N__22420\,
            in3 => \N__22474\,
            lcout => \M_this_sprites_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31957\,
            ce => 'H',
            sr => \N__27290\
        );

    \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24436\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_10_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22719\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIMJ231_8_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__25391\,
            in1 => \N__32923\,
            in2 => \N__31258\,
            in3 => \N__28031\,
            lcout => \M_this_state_q_RNIMJ231Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_19_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27940\,
            in1 => \N__25390\,
            in2 => \N__22663\,
            in3 => \N__24096\,
            lcout => \this_vga_signals.un1_M_this_state_q_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un23_i_a2_1_1_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__26400\,
            in1 => \N__31200\,
            in2 => \_gnd_net_\,
            in3 => \N__28162\,
            lcout => this_vga_signals_un23_i_a2_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNI1DGI7_0_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25962\,
            in2 => \N__24097\,
            in3 => \N__24095\,
            lcout => \M_this_sprites_address_q_RNI1DGI7Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25514\,
            in2 => \_gnd_net_\,
            in3 => \N__22621\,
            lcout => \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_0\,
            carryout => \un1_M_this_sprites_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22515\,
            in2 => \_gnd_net_\,
            in3 => \N__22477\,
            lcout => \un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_1\,
            carryout => \un1_M_this_sprites_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28262\,
            in2 => \_gnd_net_\,
            in3 => \N__22465\,
            lcout => \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_2\,
            carryout => \un1_M_this_sprites_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26166\,
            in3 => \N__22462\,
            lcout => \un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_3\,
            carryout => \un1_M_this_sprites_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24873\,
            in3 => \N__22459\,
            lcout => \un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_4\,
            carryout => \un1_M_this_sprites_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23711\,
            in2 => \_gnd_net_\,
            in3 => \N__23119\,
            lcout => \un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_5\,
            carryout => \un1_M_this_sprites_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24240\,
            in2 => \_gnd_net_\,
            in3 => \N__23116\,
            lcout => \un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_6\,
            carryout => \un1_M_this_sprites_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23010\,
            in2 => \_gnd_net_\,
            in3 => \N__22969\,
            lcout => \un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22860\,
            in2 => \_gnd_net_\,
            in3 => \N__22822\,
            lcout => \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_8\,
            carryout => \un1_M_this_sprites_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22708\,
            in2 => \_gnd_net_\,
            in3 => \N__22675\,
            lcout => \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_9\,
            carryout => \un1_M_this_sprites_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24523\,
            in2 => \_gnd_net_\,
            in3 => \N__22672\,
            lcout => \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_10\,
            carryout => \un1_M_this_sprites_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25683\,
            in3 => \N__22669\,
            lcout => \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_11\,
            carryout => \un1_M_this_sprites_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23293\,
            in2 => \_gnd_net_\,
            in3 => \N__22666\,
            lcout => \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o2_0_0_0_0_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32925\,
            in1 => \N__29595\,
            in2 => \_gnd_net_\,
            in3 => \N__24419\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_o2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_11_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__24487\,
            in1 => \N__24172\,
            in2 => \N__24607\,
            in3 => \N__23392\,
            lcout => \M_this_sprites_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31983\,
            ce => 'H',
            sr => \N__27287\
        );

    \M_this_sprites_address_q_12_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__23386\,
            in1 => \N__24173\,
            in2 => \N__25633\,
            in3 => \N__23380\,
            lcout => \M_this_sprites_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31983\,
            ce => 'H',
            sr => \N__27287\
        );

    \M_this_sprites_address_q_13_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__24174\,
            in1 => \N__23374\,
            in2 => \N__23368\,
            in3 => \N__23356\,
            lcout => \M_this_sprites_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31983\,
            ce => 'H',
            sr => \N__27287\
        );

    \this_vga_signals.M_this_map_address_q_m_9_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25218\,
            in2 => \_gnd_net_\,
            in3 => \N__27611\,
            lcout => \this_vga_signals.M_this_map_address_q_mZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o2_0_1_0_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26436\,
            in1 => \N__25396\,
            in2 => \N__27625\,
            in3 => \N__28207\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_ns_0_o2_0_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__23236\,
            in1 => \N__27960\,
            in2 => \N__23227\,
            in3 => \N__32849\,
            lcout => \N_435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_0_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__25924\,
            in1 => \N__24181\,
            in2 => \N__23671\,
            in3 => \N__23224\,
            lcout => \M_this_sprites_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31996\,
            ce => 'H',
            sr => \N__27283\
        );

    \this_sprites_ram.mem_radreg_11_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23215\,
            lcout => \this_sprites_ram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32003\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_d_5_m_9_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__25210\,
            in1 => \N__26464\,
            in2 => \N__33311\,
            in3 => \N__32850\,
            lcout => \this_vga_signals.M_this_map_address_d_5_mZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_7_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__26325\,
            in1 => \N__25177\,
            in2 => \N__25129\,
            in3 => \N__25246\,
            lcout => \M_this_map_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32010\,
            ce => 'H',
            sr => \N__27281\
        );

    \this_vga_signals.M_this_map_address_q_m_2_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24786\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26471\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_map_address_q_mZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_2_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__23623\,
            in1 => \N__26324\,
            in2 => \N__23626\,
            in3 => \N__24763\,
            lcout => \M_this_map_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32010\,
            ce => 'H',
            sr => \N__27281\
        );

    \this_vga_signals.M_this_map_address_d_8_m_2_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__24785\,
            in1 => \N__27626\,
            in2 => \N__34222\,
            in3 => \N__32848\,
            lcout => \this_vga_signals.M_this_map_address_d_8_mZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_9_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__26326\,
            in1 => \N__23617\,
            in2 => \N__23605\,
            in3 => \N__25183\,
            lcout => \M_this_map_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32010\,
            ce => 'H',
            sr => \N__27281\
        );

    \this_ppu.M_haddress_q_RNIR3M06_4_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23569\,
            in1 => \N__23919\,
            in2 => \N__23438\,
            in3 => \N__23975\,
            lcout => \this_ppu.un1_M_haddress_q_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_5_LC_18_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25080\,
            in2 => \_gnd_net_\,
            in3 => \N__25049\,
            lcout => \M_this_ppu_map_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32033\,
            ce => 'H',
            sr => \N__25034\
        );

    \this_ppu.M_haddress_q_6_LC_18_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__25050\,
            in1 => \_gnd_net_\,
            in2 => \N__25093\,
            in3 => \N__33115\,
            lcout => \M_this_ppu_vram_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32033\,
            ce => 'H',
            sr => \N__25034\
        );

    \this_ppu.M_haddress_q_4_LC_18_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__23983\,
            in1 => \N__23426\,
            in2 => \N__23930\,
            in3 => \N__23570\,
            lcout => \M_this_ppu_map_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32033\,
            ce => 'H',
            sr => \N__25034\
        );

    \this_ppu.M_haddress_q_3_LC_18_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__23427\,
            in1 => \N__23920\,
            in2 => \_gnd_net_\,
            in3 => \N__23982\,
            lcout => \M_this_ppu_map_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32033\,
            ce => 'H',
            sr => \N__25034\
        );

    \this_ppu.M_vaddress_q_RNI0655_6_LC_18_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23893\,
            lcout => \this_ppu_M_vaddress_q_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__24595\,
            in1 => \N__30754\,
            in2 => \N__23638\,
            in3 => \N__32624\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31958\,
            ce => 'H',
            sr => \N__32386\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__23695\,
            in1 => \N__28220\,
            in2 => \N__33536\,
            in3 => \N__32620\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_6_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__24150\,
            in1 => \N__23836\,
            in2 => \N__23824\,
            in3 => \N__23821\,
            lcout => \M_this_sprites_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31965\,
            ce => 'H',
            sr => \N__27292\
        );

    \this_vga_signals.M_this_sprites_address_q_m_0_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25961\,
            in2 => \_gnd_net_\,
            in3 => \N__24475\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_5_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__24835\,
            in1 => \N__24149\,
            in2 => \N__23656\,
            in3 => \N__23647\,
            lcout => \M_this_sprites_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31965\,
            ce => 'H',
            sr => \N__27292\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_0_6_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26978\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26890\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_6_0_a2_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__28199\,
            in1 => \N__24468\,
            in2 => \N__25381\,
            in3 => \N__25424\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_14_1_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001111"
        )
    port map (
            in0 => \N__34058\,
            in1 => \N__32588\,
            in2 => \N__24103\,
            in3 => \N__29181\,
            lcout => OPEN,
            ltout => \this_vga_signals.un1_M_this_state_q_14Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_14_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110000"
        )
    port map (
            in0 => \N__32589\,
            in1 => \N__27231\,
            in2 => \N__24100\,
            in3 => \N__25379\,
            lcout => \un1_M_this_state_q_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un23_i_a2_1_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__25423\,
            in1 => \N__24072\,
            in2 => \N__29606\,
            in3 => \N__30756\,
            lcout => un23_i_a2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a3_3_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__26733\,
            in1 => \N__26791\,
            in2 => \N__25903\,
            in3 => \N__25811\,
            lcout => \this_vga_signals.N_486\,
            ltout => \this_vga_signals.N_486_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__24043\,
            in1 => \N__29596\,
            in2 => \N__24019\,
            in3 => \N__32825\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31977\,
            ce => 'H',
            sr => \N__32375\
        );

    \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__26732\,
            in1 => \N__26974\,
            in2 => \N__28578\,
            in3 => \N__26790\,
            lcout => \N_465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_1_9_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__26734\,
            in1 => \N__26878\,
            in2 => \N__26991\,
            in3 => \N__26792\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_1_1_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__26786\,
            in1 => \N__25898\,
            in2 => \N__24640\,
            in3 => \N__25812\,
            lcout => \this_vga_signals.N_438_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_i_o2_0_14_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28078\,
            in2 => \_gnd_net_\,
            in3 => \N__31319\,
            lcout => \this_vga_signals_M_this_state_q_ns_i_o2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_i_o2_0_12_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28077\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31201\,
            lcout => \this_vga_signals_M_this_state_q_ns_i_o2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_11_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28226\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_1_5_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__25813\,
            in1 => \N__26716\,
            in2 => \N__26796\,
            in3 => \N__25902\,
            lcout => \this_vga_signals.N_446_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__24524\,
            in1 => \N__24476\,
            in2 => \N__33336\,
            in3 => \N__32822\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__24232\,
            in1 => \N__33794\,
            in2 => \N__24481\,
            in3 => \N__32823\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_7_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__24180\,
            in1 => \N__24211\,
            in2 => \N__24352\,
            in3 => \N__24349\,
            lcout => \M_this_sprites_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31990\,
            ce => 'H',
            sr => \N__27288\
        );

    \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28227\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_4_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__26125\,
            in1 => \N__24205\,
            in2 => \N__24196\,
            in3 => \N__24179\,
            lcout => \M_this_sprites_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31990\,
            ce => 'H',
            sr => \N__27288\
        );

    \this_vga_signals.M_this_map_address_d_5_m_5_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__24731\,
            in1 => \N__26462\,
            in2 => \N__33841\,
            in3 => \N__32755\,
            lcout => \this_vga_signals.M_this_map_address_d_5_mZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_q_m_0_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26463\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26096\,
            lcout => \this_vga_signals.M_this_map_address_q_mZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d_1_sqmuxa_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33692\,
            in1 => \N__32754\,
            in2 => \_gnd_net_\,
            in3 => \N__29190\,
            lcout => \this_vga_signals.M_this_state_d_1_sqmuxaZ0\,
            ltout => \this_vga_signals.M_this_state_d_1_sqmuxaZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_12_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__29191\,
            in1 => \N__25915\,
            in2 => \N__24643\,
            in3 => \N__27871\,
            lcout => \un1_M_this_state_q_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__26953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26715\,
            lcout => \this_vga_signals.N_399_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_8_0_a2_1_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30755\,
            in2 => \_gnd_net_\,
            in3 => \N__30636\,
            lcout => \this_vga_signals.N_293_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_q_m_6_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24677\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27627\,
            lcout => \this_vga_signals.M_this_map_address_q_mZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_q_m_5_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24732\,
            in2 => \_gnd_net_\,
            in3 => \N__27624\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_map_address_q_mZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_5_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__26328\,
            in1 => \N__24625\,
            in2 => \N__24619\,
            in3 => \N__24706\,
            lcout => \M_this_map_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32004\,
            ce => 'H',
            sr => \N__27285\
        );

    \M_this_map_address_q_0_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__26068\,
            in1 => \N__26327\,
            in2 => \N__24616\,
            in3 => \N__24817\,
            lcout => \M_this_map_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32004\,
            ce => 'H',
            sr => \N__27285\
        );

    \this_vga_signals.M_this_map_address_d_5_m_6_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__24678\,
            in1 => \N__26474\,
            in2 => \N__33990\,
            in3 => \N__32824\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_map_address_d_5_mZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_6_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__26329\,
            in1 => \N__24829\,
            in2 => \N__24820\,
            in3 => \N__24652\,
            lcout => \M_this_map_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32004\,
            ce => 'H',
            sr => \N__27285\
        );

    \M_this_map_address_q_RNICF7V6_0_LC_19_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26092\,
            in2 => \N__26362\,
            in3 => \N__26360\,
            lcout => \M_this_map_address_q_RNICF7V6Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_19_22_0_\,
            carryout => \un1_M_this_map_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_0_c_RNI6GRR_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26626\,
            in2 => \_gnd_net_\,
            in3 => \N__24811\,
            lcout => \un1_M_this_map_address_q_cry_0_c_RNI6GRRZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_0\,
            carryout => \un1_M_this_map_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_1_c_RNI8JSR_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24784\,
            in2 => \_gnd_net_\,
            in3 => \N__24757\,
            lcout => \un1_M_this_map_address_q_cry_1_c_RNI8JSRZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_1\,
            carryout => \un1_M_this_map_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_2_c_RNIAMTR_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26572\,
            in2 => \_gnd_net_\,
            in3 => \N__24754\,
            lcout => \un1_M_this_map_address_q_cry_2_c_RNIAMTRZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_2\,
            carryout => \un1_M_this_map_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_3_c_RNICPUR_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26497\,
            in2 => \_gnd_net_\,
            in3 => \N__24751\,
            lcout => \un1_M_this_map_address_q_cry_3_c_RNICPURZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_3\,
            carryout => \un1_M_this_map_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_4_c_RNIESVR_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24730\,
            in2 => \_gnd_net_\,
            in3 => \N__24700\,
            lcout => \un1_M_this_map_address_q_cry_4_c_RNIESVRZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_4\,
            carryout => \un1_M_this_map_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_5_c_RNIGV0S_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24676\,
            in2 => \_gnd_net_\,
            in3 => \N__24646\,
            lcout => \un1_M_this_map_address_q_cry_5_c_RNIGV0SZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_5\,
            carryout => \un1_M_this_map_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_6_c_RNII22S_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25161\,
            in3 => \N__25240\,
            lcout => \un1_M_this_map_address_q_cry_6_c_RNII22SZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_6\,
            carryout => \un1_M_this_map_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_7_c_RNIK53S_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27655\,
            in2 => \_gnd_net_\,
            in3 => \N__25237\,
            lcout => \un1_M_this_map_address_q_cry_7_c_RNIK53SZ0\,
            ltout => OPEN,
            carryin => \bfn_19_23_0_\,
            carryout => \un1_M_this_map_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_8_c_RNIM84S_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25214\,
            in2 => \_gnd_net_\,
            in3 => \N__25186\,
            lcout => \un1_M_this_map_address_q_cry_8_c_RNIM84SZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_d_5_m_7_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__32821\,
            in1 => \N__25156\,
            in2 => \N__34221\,
            in3 => \N__26475\,
            lcout => \this_vga_signals.M_this_map_address_d_5_mZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_q_m_7_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25157\,
            in2 => \_gnd_net_\,
            in3 => \N__27623\,
            lcout => \this_vga_signals.M_this_map_address_q_mZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_7_LC_19_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__33174\,
            in1 => \N__33116\,
            in2 => \N__25097\,
            in3 => \N__25051\,
            lcout => \this_ppu.M_haddress_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32039\,
            ce => 'H',
            sr => \N__25035\
        );

    \this_reset_cond.M_stage_q_7_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__28483\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24991\,
            lcout => \this_reset_cond.M_stage_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24982\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__24866\,
            in1 => \N__28213\,
            in2 => \N__33646\,
            in3 => \N__32746\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_i_o3_0_12_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__27030\,
            in1 => \N__27119\,
            in2 => \_gnd_net_\,
            in3 => \N__27160\,
            lcout => \this_vga_signals.N_390_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__27118\,
            in1 => \N__27158\,
            in2 => \_gnd_net_\,
            in3 => \N__27029\,
            lcout => \N_389_0\,
            ltout => \N_389_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__33999\,
            in1 => \N__25518\,
            in2 => \N__25477\,
            in3 => \N__28212\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_8_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__32916\,
            in1 => \N__25782\,
            in2 => \N__26995\,
            in3 => \N__32622\,
            lcout => \M_this_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31978\,
            ce => 'H',
            sr => \N__32376\
        );

    \this_vga_signals.un23_i_a2_0_1_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__29160\,
            in1 => \N__25462\,
            in2 => \_gnd_net_\,
            in3 => \N__25746\,
            lcout => \N_297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_9_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__32621\,
            in1 => \N__27246\,
            in2 => \N__25405\,
            in3 => \N__25380\,
            lcout => \M_this_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31978\,
            ce => 'H',
            sr => \N__32376\
        );

    \this_vga_signals.M_this_state_q_ns_0_a3_sx_9_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__25332\,
            in1 => \N__28574\,
            in2 => \N__25269\,
            in3 => \N__28076\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_ns_0_a3_sxZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a3_9_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25881\,
            in1 => \N__25839\,
            in2 => \N__25336\,
            in3 => \N__25308\,
            lcout => \this_vga_signals.N_469\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o3_8_3_0_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__25333\,
            in1 => \N__25309\,
            in2 => \N__25270\,
            in3 => \N__28075\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_5_0_a2_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28036\,
            in1 => \N__26426\,
            in2 => \N__27622\,
            in3 => \N__29162\,
            lcout => \this_vga_signals.N_291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a3_1_0_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__25810\,
            in1 => \N__25852\,
            in2 => \N__25882\,
            in3 => \N__28561\,
            lcout => \N_466\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_1_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__25876\,
            in1 => \N__25850\,
            in2 => \_gnd_net_\,
            in3 => \N__28559\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_4_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__25877\,
            in1 => \N__25851\,
            in2 => \N__26889\,
            in3 => \N__28560\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_1_4_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__26717\,
            in1 => \N__26769\,
            in2 => \N__25816\,
            in3 => \N__25809\,
            lcout => \this_vga_signals.N_444_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_14_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111110101"
        )
    port map (
            in0 => \N__26269\,
            in1 => \N__30470\,
            in2 => \N__27330\,
            in3 => \N__28804\,
            lcout => \M_this_external_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31997\,
            ce => 'H',
            sr => \N__32380\
        );

    \this_vga_signals.M_this_external_address_d_5_14_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33537\,
            in1 => \N__28825\,
            in2 => \_gnd_net_\,
            in3 => \N__32756\,
            lcout => \this_vga_signals.M_this_external_address_d_5Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_fast_14_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100010000"
        )
    port map (
            in0 => \N__32757\,
            in1 => \N__28523\,
            in2 => \N__25764\,
            in3 => \N__25747\,
            lcout => \M_this_state_q_fastZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31997\,
            ce => 'H',
            sr => \N__32380\
        );

    \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25724\,
            in3 => \N__28203\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d_0_sqmuxa_1_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__34057\,
            in1 => \N__32770\,
            in2 => \_gnd_net_\,
            in3 => \N__29188\,
            lcout => \this_vga_signals.M_this_state_d_0_sqmuxaZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_3_iv_0_14_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__30843\,
            in1 => \N__26275\,
            in2 => \N__28838\,
            in3 => \N__30675\,
            lcout => \this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__26152\,
            in1 => \N__33319\,
            in2 => \N__28222\,
            in3 => \N__32771\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_m_5_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28744\,
            in2 => \_gnd_net_\,
            in3 => \N__30676\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_d_8_m_1_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__32759\,
            in1 => \N__26627\,
            in2 => \N__33991\,
            in3 => \N__27599\,
            lcout => \this_vga_signals.M_this_map_address_d_8_mZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_d_8_m_0_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__26100\,
            in1 => \N__27597\,
            in2 => \N__33836\,
            in3 => \N__32760\,
            lcout => \this_vga_signals.M_this_map_address_d_8_mZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_q_m_4_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26499\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26453\,
            lcout => \this_vga_signals.M_this_map_address_q_mZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_d_8_m_4_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__26498\,
            in1 => \N__27598\,
            in2 => \N__33329\,
            in3 => \N__32761\,
            lcout => \this_vga_signals.M_this_map_address_d_8_mZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__32758\,
            in1 => \N__25951\,
            in2 => \N__28228\,
            in3 => \N__33827\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_q_m_1_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26473\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26628\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_map_address_q_mZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_1_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__26662\,
            in1 => \N__26306\,
            in2 => \N__26656\,
            in3 => \N__26653\,
            lcout => \M_this_map_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32019\,
            ce => 'H',
            sr => \N__27286\
        );

    \this_vga_signals.M_this_map_address_d_8_m_3_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__26574\,
            in1 => \N__27603\,
            in2 => \N__34362\,
            in3 => \N__32772\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_map_address_d_8_mZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_3_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__26307\,
            in1 => \N__26548\,
            in2 => \N__26602\,
            in3 => \N__26599\,
            lcout => \M_this_map_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32019\,
            ce => 'H',
            sr => \N__27286\
        );

    \this_vga_signals.M_this_map_address_q_m_3_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26573\,
            in2 => \_gnd_net_\,
            in3 => \N__26472\,
            lcout => \this_vga_signals.M_this_map_address_q_mZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_4_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__26542\,
            in1 => \N__26308\,
            in2 => \N__26536\,
            in3 => \N__26524\,
            lcout => \M_this_map_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32019\,
            ce => 'H',
            sr => \N__27286\
        );

    \this_vga_signals.M_this_map_address_d_5_m_8_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__27656\,
            in1 => \N__26476\,
            in2 => \N__34332\,
            in3 => \N__32854\,
            lcout => \this_vga_signals.M_this_map_address_d_5_mZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_map_ram_write_en_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33001\,
            in2 => \_gnd_net_\,
            in3 => \N__26361\,
            lcout => \this_vga_signals.un1_M_this_map_ram_write_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_8_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__26335\,
            in1 => \N__26309\,
            in2 => \N__27511\,
            in3 => \N__26281\,
            lcout => \M_this_map_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32034\,
            ce => 'H',
            sr => \N__27282\
        );

    \M_this_state_q_10_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__27250\,
            in1 => \N__32623\,
            in2 => \N__26674\,
            in3 => \N__29159\,
            lcout => \M_this_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31968\,
            ce => 'H',
            sr => \N__32381\
        );

    \M_this_state_q_15_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__27235\,
            in1 => \N__27167\,
            in2 => \N__27126\,
            in3 => \N__27042\,
            lcout => \M_this_state_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31979\,
            ce => 'H',
            sr => \N__32377\
        );

    \this_vga_signals.M_this_data_count_q_3_bm_10_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__32616\,
            in1 => \N__32432\,
            in2 => \N__33697\,
            in3 => \N__29163\,
            lcout => \this_vga_signals.M_this_data_count_q_3_bmZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_m_6_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28698\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30683\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_tr37_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001010"
        )
    port map (
            in0 => \N__28035\,
            in1 => \N__27159\,
            in2 => \N__27098\,
            in3 => \N__27043\,
            lcout => \this_vga_signals.M_this_map_ram_write_data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_21_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27044\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27086\,
            lcout => \this_start_data_delay_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31984\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_tr35_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__28041\,
            in1 => \N__27161\,
            in2 => \N__27127\,
            in3 => \N__27045\,
            lcout => \M_this_map_ram_write_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_1_10_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__26947\,
            in1 => \N__26882\,
            in2 => \N__26800\,
            in3 => \N__26724\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_2_sqmuxa_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__32625\,
            in1 => \N__33693\,
            in2 => \N__34063\,
            in3 => \N__29161\,
            lcout => \this_vga_signals.M_this_external_address_d_2_sqmuxaZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_5_13_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28876\,
            in1 => \N__33614\,
            in2 => \_gnd_net_\,
            in3 => \N__32637\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_d_5Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_3_iv_0_13_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__30669\,
            in1 => \N__30800\,
            in2 => \N__27337\,
            in3 => \N__28877\,
            lcout => \this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_bm_13_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__32750\,
            in1 => \N__32433\,
            in2 => \N__34050\,
            in3 => \N__29187\,
            lcout => \this_vga_signals.M_this_data_count_q_3_bmZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_13_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__27936\,
            in1 => \N__31150\,
            in2 => \N__27313\,
            in3 => \N__31295\,
            lcout => \M_this_state_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32005\,
            ce => 'H',
            sr => \N__32378\
        );

    \M_this_state_q_11_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__27334\,
            in1 => \N__31149\,
            in2 => \N__31199\,
            in3 => \N__32985\,
            lcout => \M_this_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32005\,
            ce => 'H',
            sr => \N__32378\
        );

    \this_vga_signals.un1_M_this_state_q_21_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__32984\,
            in1 => \N__27935\,
            in2 => \_gnd_net_\,
            in3 => \N__28785\,
            lcout => \this_vga_signals.un1_M_this_state_q_21_0\,
            ltout => \this_vga_signals.un1_M_this_state_q_21_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_13_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111011111111"
        )
    port map (
            in0 => \N__27309\,
            in1 => \N__28861\,
            in2 => \N__27301\,
            in3 => \N__27298\,
            lcout => \M_this_external_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32005\,
            ce => 'H',
            sr => \N__32378\
        );

    \this_vga_signals.M_this_external_address_q_m_4_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30685\,
            in2 => \_gnd_net_\,
            in3 => \N__30237\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_8_m_5_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__30841\,
            in1 => \N__33630\,
            in2 => \N__28749\,
            in3 => \N__32752\,
            lcout => \this_vga_signals.M_this_external_address_d_8_mZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_8_m_4_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__32751\,
            in1 => \N__30236\,
            in2 => \N__33328\,
            in3 => \N__30840\,
            lcout => \this_vga_signals.M_this_external_address_d_8_mZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_8_0_a2_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__28042\,
            in1 => \N__27961\,
            in2 => \N__27944\,
            in3 => \N__29164\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_16_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27864\,
            in2 => \N__27847\,
            in3 => \N__29082\,
            lcout => \un1_M_this_state_q_16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_13_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27844\,
            lcout => \this_sprites_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32011\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_5_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__27703\,
            in1 => \N__30487\,
            in2 => \N__27697\,
            in3 => \N__28717\,
            lcout => \M_this_external_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32020\,
            ce => 'H',
            sr => \N__32383\
        );

    \this_vga_signals.M_this_external_address_d_8_m_6_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__30842\,
            in1 => \N__28694\,
            in2 => \N__33532\,
            in3 => \N__32753\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_d_8_mZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_6_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__30488\,
            in1 => \N__27688\,
            in2 => \N__27679\,
            in3 => \N__28669\,
            lcout => \M_this_external_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32020\,
            ce => 'H',
            sr => \N__32383\
        );

    \this_vga_signals.M_this_map_address_q_m_8_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27657\,
            in2 => \_gnd_net_\,
            in3 => \N__27631\,
            lcout => \this_vga_signals.M_this_map_address_q_mZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_9_LC_22_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28466\,
            in2 => \_gnd_net_\,
            in3 => \N__28372\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_8_LC_22_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28465\,
            in2 => \_gnd_net_\,
            in3 => \N__28384\,
            lcout => \this_reset_cond.M_stage_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__28266\,
            in1 => \N__28221\,
            in2 => \N__34363\,
            in3 => \N__32773\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIV6TA_2_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29537\,
            in2 => \_gnd_net_\,
            in3 => \N__29321\,
            lcout => OPEN,
            ltout => \M_this_state_d88_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNI44LB1_0_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__29356\,
            in1 => \N__29377\,
            in2 => \N__28081\,
            in3 => \N__29065\,
            lcout => \M_this_state_d88_12\,
            ltout => \M_this_state_d88_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d_1_sqmuxa_1_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__28654\,
            in1 => \N__28074\,
            in2 => \N__28048\,
            in3 => \N__31567\,
            lcout => \this_vga_signals.N_387_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_m_7_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30978\,
            in2 => \_gnd_net_\,
            in3 => \N__30682\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32252\,
            in1 => \N__29203\,
            in2 => \N__29059\,
            in3 => \N__32154\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31991\,
            ce => \N__31676\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_1_LC_22_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33989\,
            in1 => \N__31116\,
            in2 => \_gnd_net_\,
            in3 => \N__29355\,
            lcout => OPEN,
            ltout => \N_507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_1_LC_22_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32253\,
            in1 => \N__29335\,
            in2 => \N__28045\,
            in3 => \N__32155\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31991\,
            ce => \N__31676\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_2_LC_22_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34192\,
            in1 => \N__31117\,
            in2 => \_gnd_net_\,
            in3 => \N__29325\,
            lcout => OPEN,
            ltout => \N_508_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_2_LC_22_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32254\,
            in1 => \N__29548\,
            in2 => \N__28657\,
            in3 => \N__32156\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31991\,
            ce => \N__31676\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_3_LC_22_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34358\,
            in1 => \N__31115\,
            in2 => \_gnd_net_\,
            in3 => \N__29539\,
            lcout => \N_509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a2_0_0_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33682\,
            in1 => \N__32789\,
            in2 => \N__34059\,
            in3 => \N__29180\,
            lcout => \N_436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNI60TF_15_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31404\,
            in1 => \N__32092\,
            in2 => \N__31372\,
            in3 => \N__31437\,
            lcout => \M_this_state_d88_11\,
            ltout => \M_this_state_d88_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNII1EE2_10_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31566\,
            in2 => \N__28645\,
            in3 => \N__28642\,
            lcout => \M_this_state_d88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_0_0_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__28633\,
            in1 => \N__31254\,
            in2 => \_gnd_net_\,
            in3 => \N__28504\,
            lcout => OPEN,
            ltout => \M_this_state_qsr_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__28624\,
            in1 => \N__28609\,
            in2 => \N__28597\,
            in3 => \N__28594\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32006\,
            ce => 'H',
            sr => \N__32373\
        );

    \this_vga_signals.N_570_0_i_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__31253\,
            in1 => \N__28505\,
            in2 => \_gnd_net_\,
            in3 => \N__32434\,
            lcout => \N_570_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_5_m_9_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__30891\,
            in1 => \N__30684\,
            in2 => \N__33966\,
            in3 => \N__32834\,
            lcout => \this_vga_signals.M_this_external_address_d_5_mZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNIE44V9_0_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28971\,
            in2 => \N__28786\,
            in3 => \N__28784\,
            lcout => \M_this_external_address_q_RNIE44V9Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_22_20_0_\,
            carryout => \un1_M_this_external_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_0_c_RNIGGGB_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30361\,
            in2 => \_gnd_net_\,
            in3 => \N__28765\,
            lcout => \un1_M_this_external_address_q_cry_0_c_RNIGGGBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_0\,
            carryout => \un1_M_this_external_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_1_c_RNIIJHB_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30292\,
            in2 => \_gnd_net_\,
            in3 => \N__28762\,
            lcout => \un1_M_this_external_address_q_cry_1_c_RNIIJHBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_1\,
            carryout => \un1_M_this_external_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_2_c_RNIKMIB_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29237\,
            in2 => \_gnd_net_\,
            in3 => \N__28759\,
            lcout => \un1_M_this_external_address_q_cry_2_c_RNIKMIBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_2\,
            carryout => \un1_M_this_external_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_3_c_RNIMPJB_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30227\,
            in2 => \_gnd_net_\,
            in3 => \N__28756\,
            lcout => \un1_M_this_external_address_q_cry_3_c_RNIMPJBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_3\,
            carryout => \un1_M_this_external_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_4_c_RNIOSKB_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28748\,
            in3 => \N__28711\,
            lcout => \un1_M_this_external_address_q_cry_4_c_RNIOSKBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_4\,
            carryout => \un1_M_this_external_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_5_c_RNIQVLB_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28690\,
            in2 => \_gnd_net_\,
            in3 => \N__28663\,
            lcout => \un1_M_this_external_address_q_cry_5_c_RNIQVLBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_5\,
            carryout => \un1_M_this_external_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_6_c_RNIS2NB_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30965\,
            in2 => \_gnd_net_\,
            in3 => \N__28660\,
            lcout => \un1_M_this_external_address_q_cry_6_c_RNIS2NBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_6\,
            carryout => \un1_M_this_external_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29020\,
            in2 => \_gnd_net_\,
            in3 => \N__28909\,
            lcout => \un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0\,
            ltout => OPEN,
            carryin => \bfn_22_21_0_\,
            carryout => \un1_M_this_external_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30883\,
            in2 => \_gnd_net_\,
            in3 => \N__28906\,
            lcout => \un1_M_this_external_address_q_cry_8_c_RNI09PBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_8\,
            carryout => \un1_M_this_external_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30928\,
            in2 => \_gnd_net_\,
            in3 => \N__28903\,
            lcout => \un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_9\,
            carryout => \un1_M_this_external_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29295\,
            in2 => \_gnd_net_\,
            in3 => \N__28900\,
            lcout => \un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_10\,
            carryout => \un1_M_this_external_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30426\,
            in2 => \_gnd_net_\,
            in3 => \N__28897\,
            lcout => \un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_11\,
            carryout => \un1_M_this_external_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28884\,
            in2 => \_gnd_net_\,
            in3 => \N__28852\,
            lcout => \un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_12\,
            carryout => \un1_M_this_external_address_q_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28842\,
            in2 => \_gnd_net_\,
            in3 => \N__28792\,
            lcout => \un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_13\,
            carryout => \un1_M_this_external_address_q_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30195\,
            in2 => \_gnd_net_\,
            in3 => \N__28789\,
            lcout => \un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_m_8_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29028\,
            in3 => \N__30859\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_q_mZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_8_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__30522\,
            in1 => \N__29047\,
            in2 => \N__29041\,
            in3 => \N__29002\,
            lcout => \M_this_external_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32035\,
            ce => 'H',
            sr => \N__32384\
        );

    \this_vga_signals.M_this_external_address_d_5_m_8_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__29021\,
            in1 => \N__33828\,
            in2 => \N__30698\,
            in3 => \N__32828\,
            lcout => \this_vga_signals.M_this_external_address_d_5_mZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_8_m_0_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__32829\,
            in1 => \N__28967\,
            in2 => \N__33837\,
            in3 => \N__30860\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_d_8_mZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_0_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__28945\,
            in1 => \N__30521\,
            in2 => \N__28996\,
            in3 => \N__28993\,
            lcout => \M_this_external_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32035\,
            ce => 'H',
            sr => \N__32384\
        );

    \this_vga_signals.M_this_external_address_q_m_0_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30671\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28966\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_9_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__30523\,
            in1 => \N__30706\,
            in2 => \N__28939\,
            in3 => \N__28927\,
            lcout => \M_this_external_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32035\,
            ce => 'H',
            sr => \N__32384\
        );

    \this_vga_signals.M_this_external_address_d_5_m_11_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__32853\,
            in1 => \N__29291\,
            in2 => \N__34331\,
            in3 => \N__30700\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_d_5_mZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_11_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__29269\,
            in1 => \N__30527\,
            in2 => \N__28921\,
            in3 => \N__28918\,
            lcout => \M_this_external_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32040\,
            ce => 'H',
            sr => \N__32387\
        );

    \this_vga_signals.M_this_external_address_q_m_11_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30848\,
            in2 => \_gnd_net_\,
            in3 => \N__29290\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_m_3_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29238\,
            in3 => \N__30699\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_q_mZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_3_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__30528\,
            in1 => \N__29209\,
            in2 => \N__29263\,
            in3 => \N__29260\,
            lcout => \M_this_external_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32040\,
            ce => 'H',
            sr => \N__32387\
        );

    \this_vga_signals.M_this_external_address_d_8_m_3_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__29230\,
            in1 => \N__34306\,
            in2 => \N__30861\,
            in3 => \N__32852\,
            lcout => \this_vga_signals.M_this_external_address_d_8_mZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_0_LC_22_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__29827\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29389\,
            lcout => \M_this_data_count_q_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_7_0_a2_LC_23_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__31231\,
            in1 => \N__29618\,
            in2 => \N__32932\,
            in3 => \N__29189\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_292_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_18_1_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__31128\,
            in1 => \N__31318\,
            in2 => \N__29089\,
            in3 => \N__29086\,
            lcout => \this_vga_signals.un1_M_this_state_q_18Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIAQQL_4_LC_23_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29504\,
            in1 => \N__29447\,
            in2 => \N__31057\,
            in3 => \N__29477\,
            lcout => \M_this_state_d88_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_0_LC_23_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33813\,
            in1 => \N__31100\,
            in2 => \_gnd_net_\,
            in3 => \N__29382\,
            lcout => \N_506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_5_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33637\,
            in1 => \N__31101\,
            in2 => \_gnd_net_\,
            in3 => \N__29478\,
            lcout => \N_511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_6_LC_23_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29448\,
            in1 => \N__33496\,
            in2 => \_gnd_net_\,
            in3 => \N__31102\,
            lcout => \N_512\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_3_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__29410\,
            in1 => \N__32238\,
            in2 => \N__29521\,
            in3 => \N__32157\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31998\,
            ce => \N__31668\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_4_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31107\,
            in1 => \N__33327\,
            in2 => \_gnd_net_\,
            in3 => \N__29508\,
            lcout => OPEN,
            ltout => \N_510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_4_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__29488\,
            in1 => \N__32239\,
            in2 => \N__29404\,
            in3 => \N__32158\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31998\,
            ce => \N__31668\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_5_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__32240\,
            in1 => \N__29401\,
            in2 => \N__29464\,
            in3 => \N__32159\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31998\,
            ce => \N__31668\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_6_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__32241\,
            in1 => \N__29395\,
            in2 => \N__29434\,
            in3 => \N__32160\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31998\,
            ce => \N__31668\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_c_0_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29378\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_23_17_0_\,
            carryout => \M_this_data_count_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_1_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29354\,
            in2 => \N__30071\,
            in3 => \N__29329\,
            lcout => \M_this_data_count_q_s_1\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_0\,
            carryout => \M_this_data_count_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_2_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29997\,
            in2 => \N__29326\,
            in3 => \N__29542\,
            lcout => \M_this_data_count_q_s_2\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_1\,
            carryout => \M_this_data_count_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_3_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29538\,
            in2 => \N__30072\,
            in3 => \N__29512\,
            lcout => \M_this_data_count_q_s_3\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_2\,
            carryout => \M_this_data_count_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_4_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30001\,
            in2 => \N__29509\,
            in3 => \N__29482\,
            lcout => \M_this_data_count_q_s_4\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_3\,
            carryout => \M_this_data_count_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_5_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29479\,
            in2 => \N__30073\,
            in3 => \N__29455\,
            lcout => \M_this_data_count_q_s_5\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_4\,
            carryout => \M_this_data_count_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_6_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30005\,
            in2 => \N__29452\,
            in3 => \N__29425\,
            lcout => \M_this_data_count_q_s_6\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_5\,
            carryout => \M_this_data_count_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_7_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31052\,
            in2 => \N__30074\,
            in3 => \N__29422\,
            lcout => \M_this_data_count_q_s_7\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_6\,
            carryout => \M_this_data_count_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_8_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30014\,
            in2 => \N__31591\,
            in3 => \N__29419\,
            lcout => \M_this_data_count_q_s_8\,
            ltout => OPEN,
            carryin => \bfn_23_18_0_\,
            carryout => \M_this_data_count_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_9_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31634\,
            in2 => \N__30076\,
            in3 => \N__29416\,
            lcout => \M_this_data_count_q_s_9\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_8\,
            carryout => \M_this_data_count_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_9_THRU_LUT4_0_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30021\,
            in2 => \N__31546\,
            in3 => \N__29413\,
            lcout => \M_this_data_count_q_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_9\,
            carryout => \M_this_data_count_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_11_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31610\,
            in2 => \N__30075\,
            in3 => \N__30169\,
            lcout => \M_this_data_count_q_s_11\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_10\,
            carryout => \M_this_data_count_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_12_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30012\,
            in2 => \N__31438\,
            in3 => \N__30166\,
            lcout => \M_this_data_count_q_s_12\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_11\,
            carryout => \M_this_data_count_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_12_THRU_LUT4_0_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32086\,
            in2 => \N__30077\,
            in3 => \N__30163\,
            lcout => \M_this_data_count_q_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_12\,
            carryout => \M_this_data_count_q_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_14_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30013\,
            in2 => \N__31405\,
            in3 => \N__29695\,
            lcout => \M_this_data_count_q_s_14\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_13\,
            carryout => \M_this_data_count_q_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_15_LC_23_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31367\,
            in2 => \_gnd_net_\,
            in3 => \N__29692\,
            lcout => \M_this_data_count_q_s_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_12_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29689\,
            lcout => \this_sprites_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_m_1_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30362\,
            in2 => \_gnd_net_\,
            in3 => \N__30695\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_sn_m1_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__32929\,
            in1 => \N__29619\,
            in2 => \_gnd_net_\,
            in3 => \N__32430\,
            lcout => \M_this_data_count_q_3_sn_N_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_8_m_1_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__32843\,
            in1 => \N__30363\,
            in2 => \N__33992\,
            in3 => \N__30839\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_d_8_mZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_1_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__30391\,
            in1 => \N__30518\,
            in2 => \N__30385\,
            in3 => \N__30382\,
            lcout => \M_this_external_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32026\,
            ce => 'H',
            sr => \N__32374\
        );

    \this_vga_signals.M_this_external_address_d_8_m_2_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__30838\,
            in1 => \N__30299\,
            in2 => \N__34202\,
            in3 => \N__32844\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_d_8_mZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_2_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__30519\,
            in1 => \N__30340\,
            in2 => \N__30325\,
            in3 => \N__30322\,
            lcout => \M_this_external_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32026\,
            ce => 'H',
            sr => \N__32374\
        );

    \M_this_external_address_q_4_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__30274\,
            in1 => \N__30520\,
            in2 => \N__30265\,
            in3 => \N__30253\,
            lcout => \M_this_external_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32026\,
            ce => 'H',
            sr => \N__32374\
        );

    \this_vga_signals.M_this_external_address_d_5_i_m_15_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000101010"
        )
    port map (
            in0 => \N__30696\,
            in1 => \N__32846\,
            in2 => \N__33426\,
            in3 => \N__30194\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_d_5_i_mZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_15_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__30175\,
            in1 => \N__30525\,
            in2 => \N__30214\,
            in3 => \N__30211\,
            lcout => \M_this_external_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32036\,
            ce => 'H',
            sr => \N__32379\
        );

    \this_vga_signals.M_this_external_address_q_i_m_15_LC_23_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30193\,
            in2 => \_gnd_net_\,
            in3 => \N__30852\,
            lcout => \this_vga_signals.M_this_external_address_q_i_mZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_8_m_7_LC_23_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__32845\,
            in1 => \N__33421\,
            in2 => \N__30862\,
            in3 => \N__30971\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_d_8_mZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_7_LC_23_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__30526\,
            in1 => \N__31015\,
            in2 => \N__31003\,
            in3 => \N__31000\,
            lcout => \M_this_external_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32036\,
            ce => 'H',
            sr => \N__32379\
        );

    \this_vga_signals.M_this_external_address_d_5_m_10_LC_23_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__30697\,
            in1 => \N__32847\,
            in2 => \N__34150\,
            in3 => \N__30932\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_external_address_d_5_mZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_10_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__30907\,
            in1 => \N__30524\,
            in2 => \N__30949\,
            in3 => \N__30946\,
            lcout => \M_this_external_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32036\,
            ce => 'H',
            sr => \N__32379\
        );

    \this_vga_signals.M_this_external_address_q_m_10_LC_23_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30936\,
            in2 => \_gnd_net_\,
            in3 => \N__30856\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_m_12_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30422\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_m_9_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30887\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30858\,
            lcout => \this_vga_signals.M_this_external_address_q_mZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_5_m_12_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__30421\,
            in1 => \N__30670\,
            in2 => \N__33326\,
            in3 => \N__32827\,
            lcout => \this_vga_signals.M_this_external_address_d_5_mZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_12_LC_23_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__30535\,
            in1 => \N__30529\,
            in2 => \N__30454\,
            in3 => \N__30445\,
            lcout => \M_this_external_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32044\,
            ce => 'H',
            sr => \N__32385\
        );

    \this_vga_signals.M_this_map_ram_write_data_3_LC_23_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34318\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33022\,
            lcout => \M_this_map_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_e_0_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__32931\,
            in1 => \N__32723\,
            in2 => \_gnd_net_\,
            in3 => \N__32429\,
            lcout => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o3_7_0_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31317\,
            in2 => \_gnd_net_\,
            in3 => \N__31203\,
            lcout => \N_391_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qe_0_i_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100101010"
        )
    port map (
            in0 => \N__31210\,
            in1 => \N__31204\,
            in2 => \N__31148\,
            in3 => \N__32435\,
            lcout => \M_this_data_count_qe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_7_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33390\,
            in1 => \N__31053\,
            in2 => \_gnd_net_\,
            in3 => \N__31103\,
            lcout => \N_513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_7_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__32249\,
            in1 => \N__31072\,
            in2 => \N__31066\,
            in3 => \N__32165\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32012\,
            ce => \N__31677\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_8_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33835\,
            in1 => \N__31589\,
            in2 => \_gnd_net_\,
            in3 => \N__31515\,
            lcout => OPEN,
            ltout => \N_514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_8_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32250\,
            in1 => \N__31033\,
            in2 => \N__31027\,
            in3 => \N__32166\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32012\,
            ce => \N__31677\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_9_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34000\,
            in1 => \N__31635\,
            in2 => \_gnd_net_\,
            in3 => \N__31516\,
            lcout => OPEN,
            ltout => \N_515_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_9_LC_24_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32251\,
            in1 => \N__31024\,
            in2 => \N__31018\,
            in3 => \N__32167\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32012\,
            ce => \N__31677\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_11_LC_24_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__32234\,
            in1 => \N__31348\,
            in2 => \N__31456\,
            in3 => \N__32161\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32022\,
            ce => \N__31669\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_12_LC_24_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33312\,
            in1 => \N__31436\,
            in2 => \_gnd_net_\,
            in3 => \N__31506\,
            lcout => OPEN,
            ltout => \N_518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_12_LC_24_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32235\,
            in1 => \N__31447\,
            in2 => \N__31441\,
            in3 => \N__32162\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32022\,
            ce => \N__31669\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_14_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33480\,
            in1 => \N__31403\,
            in2 => \_gnd_net_\,
            in3 => \N__31507\,
            lcout => OPEN,
            ltout => \N_520_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_14_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32236\,
            in1 => \N__31414\,
            in2 => \N__31408\,
            in3 => \N__32163\,
            lcout => \M_this_data_count_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32022\,
            ce => \N__31669\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_15_LC_24_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33406\,
            in1 => \N__31368\,
            in2 => \_gnd_net_\,
            in3 => \N__31508\,
            lcout => OPEN,
            ltout => \N_521_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_15_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32237\,
            in1 => \N__31381\,
            in2 => \N__31375\,
            in3 => \N__32164\,
            lcout => \M_this_data_count_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32022\,
            ce => \N__31669\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_11_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34357\,
            in1 => \N__31611\,
            in2 => \_gnd_net_\,
            in3 => \N__31505\,
            lcout => \N_517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_ns_10_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31342\,
            in1 => \N__32203\,
            in2 => \_gnd_net_\,
            in3 => \N__31480\,
            lcout => OPEN,
            ltout => \M_this_data_count_q_3_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_10_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010011001"
        )
    port map (
            in0 => \N__31544\,
            in1 => \N__32941\,
            in2 => \N__32935\,
            in3 => \N__32136\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32027\,
            ce => \N__31678\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_e_8_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__32930\,
            in1 => \N__32791\,
            in2 => \_gnd_net_\,
            in3 => \N__32428\,
            lcout => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8\,
            ltout => \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_am_13_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__33578\,
            in1 => \_gnd_net_\,
            in2 => \N__32269\,
            in3 => \N__32087\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_data_count_q_3_amZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_ns_13_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32266\,
            in2 => \N__32257\,
            in3 => \N__32204\,
            lcout => OPEN,
            ltout => \M_this_data_count_q_3_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010011001"
        )
    port map (
            in0 => \N__32088\,
            in1 => \N__32176\,
            in2 => \N__32170\,
            in3 => \N__32137\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32027\,
            ce => \N__31678\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNI8TRI_10_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31537\,
            in1 => \N__31636\,
            in2 => \N__31615\,
            in3 => \N__31590\,
            lcout => \M_this_state_d88_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_am_10_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34129\,
            in1 => \N__31545\,
            in2 => \_gnd_net_\,
            in3 => \N__31514\,
            lcout => \this_vga_signals.M_this_data_count_q_3_amZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_6_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33005\,
            lcout => \M_this_map_ram_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_7_LC_24_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33006\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33422\,
            lcout => \M_this_map_ram_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI5S7_7_LC_24_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33175\,
            in2 => \_gnd_net_\,
            in3 => \N__33125\,
            lcout => \M_this_ppu_map_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIIT3_6_LC_24_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33126\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_ppu_vram_addr_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_2_LC_24_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34144\,
            lcout => \M_this_map_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_1_LC_24_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33945\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33023\,
            lcout => \M_this_map_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_LC_24_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__33043\,
            in1 => \N__33814\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_map_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_5_LC_24_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33046\,
            in3 => \N__33613\,
            lcout => \M_this_map_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_4_LC_24_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33039\,
            in2 => \_gnd_net_\,
            in3 => \N__33266\,
            lcout => \M_this_map_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d21_2_LC_26_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__34343\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34151\,
            lcout => \this_vga_signals.M_this_external_address_d21Z0Z_2\,
            ltout => \this_vga_signals.M_this_external_address_d21Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d21_LC_26_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33198\,
            in1 => \N__33970\,
            in2 => \N__34066\,
            in3 => \N__33822\,
            lcout => \this_vga_signals.M_this_external_address_dZ0Z21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d22_LC_26_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33199\,
            in1 => \N__33971\,
            in2 => \N__33850\,
            in3 => \N__33823\,
            lcout => \this_vga_signals.M_this_external_address_dZ0Z22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d21_6_LC_26_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33595\,
            in1 => \N__33519\,
            in2 => \N__33389\,
            in3 => \N__33248\,
            lcout => \this_vga_signals.M_this_external_address_d21Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
