// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 8 2022 20:03:30

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    rgb,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    debug,
    clk);

    input [15:0] port_address;
    input [7:0] port_data;
    output [5:0] rgb;
    output vsync;
    output vblank;
    input rst_n;
    input port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    output debug;
    input clk;

    wire N__20240;
    wire N__20239;
    wire N__20238;
    wire N__20229;
    wire N__20228;
    wire N__20227;
    wire N__20220;
    wire N__20219;
    wire N__20218;
    wire N__20211;
    wire N__20210;
    wire N__20209;
    wire N__20202;
    wire N__20201;
    wire N__20200;
    wire N__20193;
    wire N__20192;
    wire N__20191;
    wire N__20184;
    wire N__20183;
    wire N__20182;
    wire N__20175;
    wire N__20174;
    wire N__20173;
    wire N__20166;
    wire N__20165;
    wire N__20164;
    wire N__20157;
    wire N__20156;
    wire N__20155;
    wire N__20148;
    wire N__20147;
    wire N__20146;
    wire N__20139;
    wire N__20138;
    wire N__20137;
    wire N__20130;
    wire N__20129;
    wire N__20128;
    wire N__20121;
    wire N__20120;
    wire N__20119;
    wire N__20112;
    wire N__20111;
    wire N__20110;
    wire N__20103;
    wire N__20102;
    wire N__20101;
    wire N__20094;
    wire N__20093;
    wire N__20092;
    wire N__20085;
    wire N__20084;
    wire N__20083;
    wire N__20076;
    wire N__20075;
    wire N__20074;
    wire N__20067;
    wire N__20066;
    wire N__20065;
    wire N__20058;
    wire N__20057;
    wire N__20056;
    wire N__20049;
    wire N__20048;
    wire N__20047;
    wire N__20040;
    wire N__20039;
    wire N__20038;
    wire N__20031;
    wire N__20030;
    wire N__20029;
    wire N__20022;
    wire N__20021;
    wire N__20020;
    wire N__20013;
    wire N__20012;
    wire N__20011;
    wire N__20004;
    wire N__20003;
    wire N__20002;
    wire N__19995;
    wire N__19994;
    wire N__19993;
    wire N__19986;
    wire N__19985;
    wire N__19984;
    wire N__19977;
    wire N__19976;
    wire N__19975;
    wire N__19968;
    wire N__19967;
    wire N__19966;
    wire N__19959;
    wire N__19958;
    wire N__19957;
    wire N__19950;
    wire N__19949;
    wire N__19948;
    wire N__19941;
    wire N__19940;
    wire N__19939;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19908;
    wire N__19905;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19887;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19853;
    wire N__19852;
    wire N__19851;
    wire N__19850;
    wire N__19849;
    wire N__19846;
    wire N__19839;
    wire N__19836;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19723;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19708;
    wire N__19705;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19686;
    wire N__19685;
    wire N__19680;
    wire N__19677;
    wire N__19676;
    wire N__19675;
    wire N__19672;
    wire N__19671;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19649;
    wire N__19646;
    wire N__19641;
    wire N__19640;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19613;
    wire N__19610;
    wire N__19609;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19601;
    wire N__19598;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19574;
    wire N__19571;
    wire N__19570;
    wire N__19567;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19535;
    wire N__19534;
    wire N__19533;
    wire N__19532;
    wire N__19531;
    wire N__19524;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19511;
    wire N__19510;
    wire N__19509;
    wire N__19506;
    wire N__19505;
    wire N__19504;
    wire N__19501;
    wire N__19496;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19481;
    wire N__19480;
    wire N__19479;
    wire N__19478;
    wire N__19477;
    wire N__19476;
    wire N__19475;
    wire N__19474;
    wire N__19473;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19469;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19449;
    wire N__19446;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19434;
    wire N__19429;
    wire N__19426;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19379;
    wire N__19378;
    wire N__19377;
    wire N__19376;
    wire N__19375;
    wire N__19370;
    wire N__19363;
    wire N__19358;
    wire N__19353;
    wire N__19346;
    wire N__19341;
    wire N__19336;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19316;
    wire N__19311;
    wire N__19308;
    wire N__19303;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19280;
    wire N__19277;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19269;
    wire N__19264;
    wire N__19261;
    wire N__19260;
    wire N__19255;
    wire N__19252;
    wire N__19251;
    wire N__19250;
    wire N__19245;
    wire N__19242;
    wire N__19241;
    wire N__19238;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19222;
    wire N__19221;
    wire N__19220;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19202;
    wire N__19201;
    wire N__19200;
    wire N__19199;
    wire N__19198;
    wire N__19197;
    wire N__19196;
    wire N__19195;
    wire N__19194;
    wire N__19193;
    wire N__19192;
    wire N__19191;
    wire N__19190;
    wire N__19189;
    wire N__19188;
    wire N__19187;
    wire N__19186;
    wire N__19185;
    wire N__19184;
    wire N__19183;
    wire N__19182;
    wire N__19181;
    wire N__19180;
    wire N__19179;
    wire N__19178;
    wire N__19177;
    wire N__19176;
    wire N__19175;
    wire N__19174;
    wire N__19173;
    wire N__19172;
    wire N__19171;
    wire N__19170;
    wire N__19169;
    wire N__19168;
    wire N__19167;
    wire N__19166;
    wire N__19165;
    wire N__19164;
    wire N__19163;
    wire N__19162;
    wire N__19161;
    wire N__19160;
    wire N__19159;
    wire N__19158;
    wire N__19157;
    wire N__19156;
    wire N__19155;
    wire N__19154;
    wire N__19153;
    wire N__19152;
    wire N__19151;
    wire N__19150;
    wire N__19149;
    wire N__19148;
    wire N__19147;
    wire N__19146;
    wire N__19145;
    wire N__19144;
    wire N__19143;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19139;
    wire N__19138;
    wire N__19137;
    wire N__19136;
    wire N__19135;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19131;
    wire N__19130;
    wire N__19129;
    wire N__19128;
    wire N__19127;
    wire N__19126;
    wire N__19125;
    wire N__19124;
    wire N__19123;
    wire N__19122;
    wire N__19121;
    wire N__19120;
    wire N__19119;
    wire N__19118;
    wire N__19117;
    wire N__19116;
    wire N__19115;
    wire N__19114;
    wire N__19113;
    wire N__19112;
    wire N__19111;
    wire N__19110;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18859;
    wire N__18856;
    wire N__18853;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18603;
    wire N__18598;
    wire N__18595;
    wire N__18594;
    wire N__18589;
    wire N__18586;
    wire N__18585;
    wire N__18580;
    wire N__18577;
    wire N__18576;
    wire N__18575;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18559;
    wire N__18556;
    wire N__18555;
    wire N__18554;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18318;
    wire N__18317;
    wire N__18316;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18301;
    wire N__18296;
    wire N__18291;
    wire N__18288;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18156;
    wire N__18151;
    wire N__18148;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18021;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17881;
    wire N__17880;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17869;
    wire N__17868;
    wire N__17865;
    wire N__17860;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17816;
    wire N__17815;
    wire N__17812;
    wire N__17809;
    wire N__17808;
    wire N__17807;
    wire N__17806;
    wire N__17805;
    wire N__17804;
    wire N__17803;
    wire N__17802;
    wire N__17801;
    wire N__17800;
    wire N__17799;
    wire N__17798;
    wire N__17797;
    wire N__17796;
    wire N__17795;
    wire N__17794;
    wire N__17793;
    wire N__17792;
    wire N__17791;
    wire N__17788;
    wire N__17785;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17725;
    wire N__17724;
    wire N__17721;
    wire N__17720;
    wire N__17715;
    wire N__17712;
    wire N__17709;
    wire N__17706;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17662;
    wire N__17659;
    wire N__17658;
    wire N__17655;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17644;
    wire N__17643;
    wire N__17640;
    wire N__17639;
    wire N__17638;
    wire N__17637;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17622;
    wire N__17619;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17351;
    wire N__17348;
    wire N__17347;
    wire N__17346;
    wire N__17345;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17331;
    wire N__17330;
    wire N__17327;
    wire N__17322;
    wire N__17319;
    wire N__17318;
    wire N__17317;
    wire N__17314;
    wire N__17309;
    wire N__17304;
    wire N__17297;
    wire N__17294;
    wire N__17293;
    wire N__17292;
    wire N__17291;
    wire N__17290;
    wire N__17289;
    wire N__17288;
    wire N__17285;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17255;
    wire N__17252;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17232;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17218;
    wire N__17217;
    wire N__17216;
    wire N__17215;
    wire N__17214;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17202;
    wire N__17195;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17164;
    wire N__17161;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17146;
    wire N__17143;
    wire N__17132;
    wire N__17129;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16972;
    wire N__16969;
    wire N__16968;
    wire N__16967;
    wire N__16966;
    wire N__16965;
    wire N__16962;
    wire N__16959;
    wire N__16956;
    wire N__16955;
    wire N__16954;
    wire N__16947;
    wire N__16944;
    wire N__16939;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16923;
    wire N__16916;
    wire N__16913;
    wire N__16912;
    wire N__16909;
    wire N__16906;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16735;
    wire N__16734;
    wire N__16733;
    wire N__16732;
    wire N__16731;
    wire N__16730;
    wire N__16725;
    wire N__16722;
    wire N__16717;
    wire N__16712;
    wire N__16711;
    wire N__16704;
    wire N__16701;
    wire N__16698;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16601;
    wire N__16598;
    wire N__16597;
    wire N__16594;
    wire N__16591;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16519;
    wire N__16516;
    wire N__16515;
    wire N__16514;
    wire N__16513;
    wire N__16512;
    wire N__16509;
    wire N__16508;
    wire N__16507;
    wire N__16506;
    wire N__16505;
    wire N__16502;
    wire N__16497;
    wire N__16492;
    wire N__16489;
    wire N__16480;
    wire N__16479;
    wire N__16478;
    wire N__16477;
    wire N__16476;
    wire N__16475;
    wire N__16474;
    wire N__16469;
    wire N__16466;
    wire N__16461;
    wire N__16452;
    wire N__16447;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16405;
    wire N__16402;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16387;
    wire N__16382;
    wire N__16379;
    wire N__16378;
    wire N__16377;
    wire N__16372;
    wire N__16371;
    wire N__16370;
    wire N__16369;
    wire N__16366;
    wire N__16365;
    wire N__16364;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16349;
    wire N__16348;
    wire N__16347;
    wire N__16346;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16334;
    wire N__16329;
    wire N__16326;
    wire N__16321;
    wire N__16314;
    wire N__16311;
    wire N__16310;
    wire N__16309;
    wire N__16308;
    wire N__16305;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16293;
    wire N__16290;
    wire N__16285;
    wire N__16282;
    wire N__16275;
    wire N__16272;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16252;
    wire N__16241;
    wire N__16240;
    wire N__16239;
    wire N__16238;
    wire N__16237;
    wire N__16236;
    wire N__16235;
    wire N__16220;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16199;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15905;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15865;
    wire N__15864;
    wire N__15863;
    wire N__15860;
    wire N__15857;
    wire N__15856;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15835;
    wire N__15832;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15814;
    wire N__15811;
    wire N__15808;
    wire N__15803;
    wire N__15800;
    wire N__15799;
    wire N__15796;
    wire N__15793;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15731;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15611;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15593;
    wire N__15590;
    wire N__15589;
    wire N__15588;
    wire N__15585;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15567;
    wire N__15566;
    wire N__15565;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15469;
    wire N__15468;
    wire N__15467;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15459;
    wire N__15458;
    wire N__15457;
    wire N__15456;
    wire N__15455;
    wire N__15454;
    wire N__15453;
    wire N__15452;
    wire N__15447;
    wire N__15444;
    wire N__15439;
    wire N__15434;
    wire N__15429;
    wire N__15424;
    wire N__15419;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15397;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15376;
    wire N__15373;
    wire N__15370;
    wire N__15365;
    wire N__15362;
    wire N__15361;
    wire N__15356;
    wire N__15353;
    wire N__15352;
    wire N__15351;
    wire N__15350;
    wire N__15349;
    wire N__15348;
    wire N__15347;
    wire N__15346;
    wire N__15345;
    wire N__15340;
    wire N__15335;
    wire N__15334;
    wire N__15333;
    wire N__15330;
    wire N__15329;
    wire N__15328;
    wire N__15323;
    wire N__15322;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15301;
    wire N__15300;
    wire N__15299;
    wire N__15298;
    wire N__15297;
    wire N__15294;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15264;
    wire N__15255;
    wire N__15250;
    wire N__15241;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15207;
    wire N__15206;
    wire N__15205;
    wire N__15204;
    wire N__15201;
    wire N__15200;
    wire N__15197;
    wire N__15192;
    wire N__15191;
    wire N__15190;
    wire N__15189;
    wire N__15188;
    wire N__15187;
    wire N__15186;
    wire N__15185;
    wire N__15180;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15159;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15125;
    wire N__15124;
    wire N__15123;
    wire N__15122;
    wire N__15121;
    wire N__15120;
    wire N__15119;
    wire N__15118;
    wire N__15117;
    wire N__15114;
    wire N__15113;
    wire N__15112;
    wire N__15111;
    wire N__15106;
    wire N__15105;
    wire N__15102;
    wire N__15101;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15093;
    wire N__15092;
    wire N__15091;
    wire N__15090;
    wire N__15089;
    wire N__15086;
    wire N__15085;
    wire N__15084;
    wire N__15083;
    wire N__15082;
    wire N__15079;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15055;
    wire N__15050;
    wire N__15047;
    wire N__15046;
    wire N__15045;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15033;
    wire N__15026;
    wire N__15019;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__15001;
    wire N__15000;
    wire N__14999;
    wire N__14996;
    wire N__14991;
    wire N__14984;
    wire N__14977;
    wire N__14964;
    wire N__14961;
    wire N__14958;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14936;
    wire N__14931;
    wire N__14920;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14875;
    wire N__14874;
    wire N__14873;
    wire N__14872;
    wire N__14871;
    wire N__14870;
    wire N__14867;
    wire N__14862;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14831;
    wire N__14830;
    wire N__14829;
    wire N__14828;
    wire N__14827;
    wire N__14826;
    wire N__14825;
    wire N__14824;
    wire N__14823;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14801;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14782;
    wire N__14779;
    wire N__14768;
    wire N__14767;
    wire N__14766;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14758;
    wire N__14757;
    wire N__14756;
    wire N__14755;
    wire N__14754;
    wire N__14753;
    wire N__14750;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14724;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14708;
    wire N__14707;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14672;
    wire N__14671;
    wire N__14670;
    wire N__14669;
    wire N__14668;
    wire N__14667;
    wire N__14666;
    wire N__14665;
    wire N__14664;
    wire N__14661;
    wire N__14660;
    wire N__14657;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14645;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14629;
    wire N__14626;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14593;
    wire N__14592;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14570;
    wire N__14567;
    wire N__14566;
    wire N__14565;
    wire N__14558;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14528;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14516;
    wire N__14515;
    wire N__14512;
    wire N__14511;
    wire N__14510;
    wire N__14509;
    wire N__14508;
    wire N__14507;
    wire N__14506;
    wire N__14505;
    wire N__14504;
    wire N__14503;
    wire N__14502;
    wire N__14501;
    wire N__14500;
    wire N__14499;
    wire N__14498;
    wire N__14497;
    wire N__14496;
    wire N__14495;
    wire N__14494;
    wire N__14493;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14482;
    wire N__14481;
    wire N__14478;
    wire N__14477;
    wire N__14476;
    wire N__14475;
    wire N__14472;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14454;
    wire N__14449;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14437;
    wire N__14436;
    wire N__14427;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14413;
    wire N__14406;
    wire N__14403;
    wire N__14400;
    wire N__14397;
    wire N__14394;
    wire N__14391;
    wire N__14388;
    wire N__14385;
    wire N__14382;
    wire N__14377;
    wire N__14374;
    wire N__14367;
    wire N__14364;
    wire N__14351;
    wire N__14340;
    wire N__14339;
    wire N__14336;
    wire N__14329;
    wire N__14324;
    wire N__14321;
    wire N__14316;
    wire N__14313;
    wire N__14310;
    wire N__14307;
    wire N__14302;
    wire N__14299;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14199;
    wire N__14196;
    wire N__14193;
    wire N__14190;
    wire N__14189;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14177;
    wire N__14172;
    wire N__14169;
    wire N__14166;
    wire N__14165;
    wire N__14160;
    wire N__14157;
    wire N__14154;
    wire N__14153;
    wire N__14152;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14133;
    wire N__14130;
    wire N__14127;
    wire N__14126;
    wire N__14119;
    wire N__14116;
    wire N__14111;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14100;
    wire N__14099;
    wire N__14094;
    wire N__14093;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14082;
    wire N__14077;
    wire N__14072;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14058;
    wire N__14051;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14036;
    wire N__14033;
    wire N__14032;
    wire N__14031;
    wire N__14030;
    wire N__14029;
    wire N__14028;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14020;
    wire N__14017;
    wire N__14010;
    wire N__14007;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13991;
    wire N__13986;
    wire N__13979;
    wire N__13976;
    wire N__13975;
    wire N__13974;
    wire N__13973;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13965;
    wire N__13964;
    wire N__13963;
    wire N__13962;
    wire N__13961;
    wire N__13960;
    wire N__13959;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13948;
    wire N__13945;
    wire N__13944;
    wire N__13941;
    wire N__13936;
    wire N__13933;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13915;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13896;
    wire N__13895;
    wire N__13894;
    wire N__13891;
    wire N__13882;
    wire N__13879;
    wire N__13878;
    wire N__13871;
    wire N__13866;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13850;
    wire N__13847;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13828;
    wire N__13825;
    wire N__13820;
    wire N__13817;
    wire N__13816;
    wire N__13815;
    wire N__13812;
    wire N__13811;
    wire N__13810;
    wire N__13809;
    wire N__13806;
    wire N__13805;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13778;
    wire N__13763;
    wire N__13762;
    wire N__13761;
    wire N__13760;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13720;
    wire N__13717;
    wire N__13706;
    wire N__13705;
    wire N__13704;
    wire N__13703;
    wire N__13696;
    wire N__13693;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13678;
    wire N__13677;
    wire N__13674;
    wire N__13673;
    wire N__13670;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13659;
    wire N__13658;
    wire N__13657;
    wire N__13656;
    wire N__13655;
    wire N__13654;
    wire N__13653;
    wire N__13652;
    wire N__13651;
    wire N__13648;
    wire N__13645;
    wire N__13640;
    wire N__13637;
    wire N__13628;
    wire N__13617;
    wire N__13604;
    wire N__13601;
    wire N__13600;
    wire N__13599;
    wire N__13596;
    wire N__13595;
    wire N__13592;
    wire N__13591;
    wire N__13588;
    wire N__13585;
    wire N__13582;
    wire N__13581;
    wire N__13580;
    wire N__13579;
    wire N__13578;
    wire N__13577;
    wire N__13576;
    wire N__13575;
    wire N__13574;
    wire N__13573;
    wire N__13570;
    wire N__13567;
    wire N__13562;
    wire N__13559;
    wire N__13552;
    wire N__13547;
    wire N__13542;
    wire N__13537;
    wire N__13520;
    wire N__13517;
    wire N__13516;
    wire N__13515;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13507;
    wire N__13504;
    wire N__13503;
    wire N__13502;
    wire N__13501;
    wire N__13498;
    wire N__13497;
    wire N__13494;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13483;
    wire N__13480;
    wire N__13477;
    wire N__13476;
    wire N__13475;
    wire N__13472;
    wire N__13471;
    wire N__13470;
    wire N__13465;
    wire N__13462;
    wire N__13459;
    wire N__13456;
    wire N__13453;
    wire N__13450;
    wire N__13445;
    wire N__13436;
    wire N__13431;
    wire N__13426;
    wire N__13409;
    wire N__13406;
    wire N__13405;
    wire N__13404;
    wire N__13403;
    wire N__13402;
    wire N__13399;
    wire N__13398;
    wire N__13395;
    wire N__13392;
    wire N__13387;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13383;
    wire N__13382;
    wire N__13381;
    wire N__13380;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13365;
    wire N__13354;
    wire N__13347;
    wire N__13344;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13213;
    wire N__13210;
    wire N__13209;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13187;
    wire N__13186;
    wire N__13185;
    wire N__13184;
    wire N__13181;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13169;
    wire N__13168;
    wire N__13167;
    wire N__13166;
    wire N__13165;
    wire N__13162;
    wire N__13159;
    wire N__13154;
    wire N__13149;
    wire N__13146;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13129;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13110;
    wire N__13105;
    wire N__13102;
    wire N__13099;
    wire N__13094;
    wire N__13093;
    wire N__13092;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13079;
    wire N__13074;
    wire N__13067;
    wire N__13066;
    wire N__13065;
    wire N__13064;
    wire N__13063;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13052;
    wire N__13047;
    wire N__13046;
    wire N__13045;
    wire N__13042;
    wire N__13039;
    wire N__13034;
    wire N__13031;
    wire N__13028;
    wire N__13023;
    wire N__13018;
    wire N__13015;
    wire N__13004;
    wire N__13003;
    wire N__12998;
    wire N__12995;
    wire N__12994;
    wire N__12991;
    wire N__12990;
    wire N__12989;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12975;
    wire N__12972;
    wire N__12965;
    wire N__12964;
    wire N__12963;
    wire N__12962;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12949;
    wire N__12940;
    wire N__12935;
    wire N__12934;
    wire N__12931;
    wire N__12928;
    wire N__12923;
    wire N__12920;
    wire N__12919;
    wire N__12918;
    wire N__12917;
    wire N__12912;
    wire N__12907;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12892;
    wire N__12887;
    wire N__12886;
    wire N__12883;
    wire N__12882;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12870;
    wire N__12863;
    wire N__12862;
    wire N__12861;
    wire N__12860;
    wire N__12859;
    wire N__12858;
    wire N__12857;
    wire N__12852;
    wire N__12845;
    wire N__12840;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12808;
    wire N__12805;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12787;
    wire N__12782;
    wire N__12779;
    wire N__12778;
    wire N__12775;
    wire N__12772;
    wire N__12767;
    wire N__12764;
    wire N__12763;
    wire N__12760;
    wire N__12757;
    wire N__12754;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12739;
    wire N__12738;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12726;
    wire N__12719;
    wire N__12718;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12701;
    wire N__12700;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12664;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12646;
    wire N__12645;
    wire N__12642;
    wire N__12637;
    wire N__12632;
    wire N__12631;
    wire N__12630;
    wire N__12629;
    wire N__12628;
    wire N__12627;
    wire N__12624;
    wire N__12623;
    wire N__12622;
    wire N__12621;
    wire N__12620;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12608;
    wire N__12607;
    wire N__12606;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12598;
    wire N__12595;
    wire N__12594;
    wire N__12593;
    wire N__12588;
    wire N__12587;
    wire N__12586;
    wire N__12585;
    wire N__12584;
    wire N__12581;
    wire N__12576;
    wire N__12573;
    wire N__12568;
    wire N__12565;
    wire N__12564;
    wire N__12563;
    wire N__12560;
    wire N__12559;
    wire N__12558;
    wire N__12557;
    wire N__12556;
    wire N__12555;
    wire N__12554;
    wire N__12549;
    wire N__12546;
    wire N__12541;
    wire N__12538;
    wire N__12535;
    wire N__12526;
    wire N__12519;
    wire N__12514;
    wire N__12509;
    wire N__12502;
    wire N__12495;
    wire N__12492;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12454;
    wire N__12451;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12431;
    wire N__12428;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12420;
    wire N__12417;
    wire N__12416;
    wire N__12413;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12399;
    wire N__12398;
    wire N__12393;
    wire N__12388;
    wire N__12385;
    wire N__12380;
    wire N__12377;
    wire N__12368;
    wire N__12367;
    wire N__12364;
    wire N__12363;
    wire N__12362;
    wire N__12359;
    wire N__12358;
    wire N__12357;
    wire N__12356;
    wire N__12355;
    wire N__12354;
    wire N__12353;
    wire N__12352;
    wire N__12349;
    wire N__12348;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12332;
    wire N__12329;
    wire N__12324;
    wire N__12323;
    wire N__12322;
    wire N__12319;
    wire N__12318;
    wire N__12317;
    wire N__12316;
    wire N__12315;
    wire N__12314;
    wire N__12313;
    wire N__12312;
    wire N__12311;
    wire N__12310;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12291;
    wire N__12290;
    wire N__12289;
    wire N__12288;
    wire N__12287;
    wire N__12286;
    wire N__12285;
    wire N__12284;
    wire N__12279;
    wire N__12274;
    wire N__12271;
    wire N__12266;
    wire N__12259;
    wire N__12256;
    wire N__12247;
    wire N__12236;
    wire N__12229;
    wire N__12226;
    wire N__12217;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12073;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12044;
    wire N__12043;
    wire N__12040;
    wire N__12037;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12019;
    wire N__12016;
    wire N__12015;
    wire N__12012;
    wire N__12007;
    wire N__12004;
    wire N__11999;
    wire N__11996;
    wire N__11995;
    wire N__11992;
    wire N__11989;
    wire N__11986;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11962;
    wire N__11959;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11942;
    wire N__11941;
    wire N__11940;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11906;
    wire N__11903;
    wire N__11900;
    wire N__11897;
    wire N__11896;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11867;
    wire N__11864;
    wire N__11863;
    wire N__11862;
    wire N__11857;
    wire N__11854;
    wire N__11849;
    wire N__11848;
    wire N__11843;
    wire N__11842;
    wire N__11841;
    wire N__11838;
    wire N__11833;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11812;
    wire N__11811;
    wire N__11808;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11796;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11765;
    wire N__11764;
    wire N__11763;
    wire N__11758;
    wire N__11755;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11714;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11702;
    wire N__11701;
    wire N__11700;
    wire N__11699;
    wire N__11698;
    wire N__11695;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11678;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11651;
    wire N__11648;
    wire N__11641;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11494;
    wire N__11493;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11459;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11441;
    wire N__11438;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11414;
    wire N__11413;
    wire N__11410;
    wire N__11409;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11397;
    wire N__11390;
    wire N__11389;
    wire N__11386;
    wire N__11383;
    wire N__11378;
    wire N__11375;
    wire N__11374;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11366;
    wire N__11363;
    wire N__11362;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11278;
    wire N__11277;
    wire N__11272;
    wire N__11269;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11194;
    wire N__11193;
    wire N__11188;
    wire N__11185;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10928;
    wire N__10927;
    wire N__10924;
    wire N__10921;
    wire N__10916;
    wire N__10913;
    wire N__10912;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10882;
    wire N__10881;
    wire N__10880;
    wire N__10879;
    wire N__10878;
    wire N__10875;
    wire N__10874;
    wire N__10873;
    wire N__10868;
    wire N__10867;
    wire N__10866;
    wire N__10863;
    wire N__10862;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10858;
    wire N__10855;
    wire N__10854;
    wire N__10851;
    wire N__10848;
    wire N__10843;
    wire N__10840;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10824;
    wire N__10815;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10744;
    wire N__10743;
    wire N__10742;
    wire N__10735;
    wire N__10734;
    wire N__10733;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10706;
    wire N__10703;
    wire N__10702;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10579;
    wire N__10578;
    wire N__10577;
    wire N__10576;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10564;
    wire N__10559;
    wire N__10556;
    wire N__10547;
    wire N__10546;
    wire N__10545;
    wire N__10544;
    wire N__10539;
    wire N__10534;
    wire N__10529;
    wire N__10526;
    wire N__10525;
    wire N__10524;
    wire N__10523;
    wire N__10522;
    wire N__10519;
    wire N__10516;
    wire N__10509;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10387;
    wire N__10384;
    wire N__10383;
    wire N__10378;
    wire N__10375;
    wire N__10370;
    wire N__10369;
    wire N__10368;
    wire N__10367;
    wire N__10360;
    wire N__10357;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10342;
    wire N__10339;
    wire N__10336;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10204;
    wire N__10203;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10181;
    wire N__10178;
    wire N__10177;
    wire N__10176;
    wire N__10175;
    wire N__10174;
    wire N__10171;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10030;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10006;
    wire N__10005;
    wire N__10002;
    wire N__10001;
    wire N__10000;
    wire N__9999;
    wire N__9996;
    wire N__9995;
    wire N__9992;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9957;
    wire N__9944;
    wire N__9941;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9933;
    wire N__9932;
    wire N__9925;
    wire N__9924;
    wire N__9923;
    wire N__9922;
    wire N__9921;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9901;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9874;
    wire N__9871;
    wire N__9868;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9832;
    wire N__9831;
    wire N__9828;
    wire N__9825;
    wire N__9824;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9816;
    wire N__9813;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9774;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9595;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9575;
    wire N__9572;
    wire N__9571;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9551;
    wire N__9548;
    wire N__9547;
    wire N__9546;
    wire N__9545;
    wire N__9542;
    wire N__9537;
    wire N__9534;
    wire N__9527;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9521;
    wire N__9520;
    wire N__9517;
    wire N__9512;
    wire N__9507;
    wire N__9506;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9481;
    wire N__9480;
    wire N__9477;
    wire N__9472;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9409;
    wire N__9404;
    wire N__9401;
    wire N__9396;
    wire N__9389;
    wire N__9386;
    wire N__9385;
    wire N__9382;
    wire N__9381;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9365;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9353;
    wire N__9350;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9338;
    wire N__9335;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9320;
    wire N__9317;
    wire N__9316;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9299;
    wire N__9296;
    wire N__9295;
    wire N__9294;
    wire N__9293;
    wire N__9290;
    wire N__9283;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8960;
    wire N__8957;
    wire N__8956;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8929;
    wire N__8928;
    wire N__8925;
    wire N__8920;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8908;
    wire N__8907;
    wire N__8906;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8869;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8851;
    wire N__8850;
    wire N__8847;
    wire N__8842;
    wire N__8837;
    wire N__8836;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8819;
    wire N__8816;
    wire N__8815;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8800;
    wire N__8799;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8787;
    wire N__8780;
    wire N__8779;
    wire N__8778;
    wire N__8775;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8747;
    wire N__8744;
    wire N__8743;
    wire N__8738;
    wire N__8735;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8723;
    wire N__8720;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8708;
    wire N__8707;
    wire N__8704;
    wire N__8701;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8614;
    wire N__8613;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8592;
    wire N__8585;
    wire N__8584;
    wire N__8583;
    wire N__8582;
    wire N__8581;
    wire N__8578;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8559;
    wire N__8552;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8540;
    wire N__8537;
    wire N__8536;
    wire N__8535;
    wire N__8534;
    wire N__8531;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8517;
    wire N__8510;
    wire N__8509;
    wire N__8508;
    wire N__8507;
    wire N__8506;
    wire N__8503;
    wire N__8502;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8480;
    wire N__8477;
    wire N__8476;
    wire N__8473;
    wire N__8472;
    wire N__8471;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8454;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8416;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8408;
    wire N__8407;
    wire N__8406;
    wire N__8403;
    wire N__8398;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8378;
    wire N__8377;
    wire N__8376;
    wire N__8373;
    wire N__8372;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8339;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8331;
    wire N__8330;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8309;
    wire N__8304;
    wire N__8297;
    wire N__8296;
    wire N__8295;
    wire N__8294;
    wire N__8291;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8242;
    wire N__8239;
    wire N__8234;
    wire N__8231;
    wire N__8230;
    wire N__8229;
    wire N__8228;
    wire N__8227;
    wire N__8222;
    wire N__8217;
    wire N__8214;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8159;
    wire N__8158;
    wire N__8155;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8096;
    wire N__8095;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8078;
    wire N__8077;
    wire N__8076;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8054;
    wire N__8053;
    wire N__8050;
    wire N__8049;
    wire N__8046;
    wire N__8045;
    wire N__8042;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7936;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7890;
    wire N__7887;
    wire N__7884;
    wire N__7881;
    wire N__7880;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7843;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7804;
    wire N__7799;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7762;
    wire N__7761;
    wire N__7756;
    wire N__7753;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7739;
    wire N__7736;
    wire N__7733;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7639;
    wire N__7638;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7621;
    wire N__7618;
    wire N__7615;
    wire N__7612;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7589;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7417;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7406;
    wire N__7405;
    wire N__7404;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7390;
    wire N__7389;
    wire N__7386;
    wire N__7385;
    wire N__7384;
    wire N__7377;
    wire N__7374;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7360;
    wire N__7359;
    wire N__7354;
    wire N__7351;
    wire N__7350;
    wire N__7349;
    wire N__7346;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7332;
    wire N__7331;
    wire N__7330;
    wire N__7329;
    wire N__7324;
    wire N__7321;
    wire N__7320;
    wire N__7317;
    wire N__7316;
    wire N__7315;
    wire N__7314;
    wire N__7305;
    wire N__7302;
    wire N__7299;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7287;
    wire N__7284;
    wire N__7283;
    wire N__7282;
    wire N__7281;
    wire N__7278;
    wire N__7275;
    wire N__7274;
    wire N__7273;
    wire N__7270;
    wire N__7269;
    wire N__7266;
    wire N__7259;
    wire N__7256;
    wire N__7255;
    wire N__7252;
    wire N__7245;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7218;
    wire N__7215;
    wire N__7210;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7185;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7147;
    wire N__7144;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7115;
    wire N__7112;
    wire N__7109;
    wire N__7104;
    wire N__7101;
    wire VCCG0;
    wire GNDG0;
    wire port_rw_c_i;
    wire CONSTANT_ONE_NET;
    wire this_vga_signals_M_hstate_q_i_1;
    wire port_nmib_c_i;
    wire rgb_c_2;
    wire rgb_c_5;
    wire this_vga_signals_M_hstate_q_i_4;
    wire rgb_c_4;
    wire rgb_c_0;
    wire m5;
    wire rgb_c_1;
    wire rgb_2_5_0__i2_mux_0;
    wire rgb_2_5_0__i2_mux;
    wire m19;
    wire rgb72;
    wire rgb_c_3;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_0 ;
    wire port_clk_c;
    wire this_start_data_delay_this_edge_detector_M_last_q;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_0 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_1 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_2 ;
    wire m16;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_8 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_6 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_7 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_5 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_3 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_4 ;
    wire bfn_13_17_0_;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_7 ;
    wire bfn_13_18_0_;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_CO ;
    wire \this_vga_signals.N_238_0_cascade_ ;
    wire \this_vga_signals.N_221_0_cascade_ ;
    wire \this_vga_signals.N_232_0 ;
    wire \this_vga_signals.N_237_0_cascade_ ;
    wire \this_vga_signals.M_vstate_d_0_sqmuxa ;
    wire \this_vga_signals.N_221_0 ;
    wire \this_vga_signals.N_225_0 ;
    wire \this_vga_signals.N_225_0_cascade_ ;
    wire \this_vga_signals.N_239_0 ;
    wire \this_vga_signals.N_239_0_cascade_ ;
    wire port_nmib_c;
    wire \this_vga_signals.N_258_cascade_ ;
    wire \this_vga_signals.N_238_0 ;
    wire \this_vga_signals.M_vstate_qZ0Z_2 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_1 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_6 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_2 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_3 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_4 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_5 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_13 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_11 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_12 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_9 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_10 ;
    wire \this_vga_signals.M_vstate_q_RNI3M6M4Z0Z_0 ;
    wire \this_vga_signals.N_251_cascade_ ;
    wire \this_vga_signals.N_237_0 ;
    wire \this_vga_signals.M_vstate_qZ0Z_0 ;
    wire \this_vga_signals.M_vstate_q_srsts_0_a4_0_4_cascade_ ;
    wire \this_vga_signals.M_vstate_q_srsts_0_a4_0_4 ;
    wire \this_vga_signals.N_230_0_cascade_ ;
    wire vsync_c;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.N_230_0 ;
    wire \this_vga_signals.M_vstate_q_srsts_0_o2_2_5_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.N_248_0 ;
    wire \this_vga_signals.N_248_0_cascade_ ;
    wire \this_vga_signals.M_vstate_qZ0Z_5 ;
    wire \this_vga_signals.N_252 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_vstate_q_srsts_0_o2_2_3_cascade_ ;
    wire \this_vga_signals.N_255 ;
    wire \this_vga_signals.M_vstate_q_srsts_0_o2_2_3 ;
    wire \this_vga_signals.M_vstate_qZ0Z_3 ;
    wire \this_vga_signals.N_226_0 ;
    wire \this_vga_signals.N_256 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_7 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_10 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_11 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_8 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_9 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_14 ;
    wire \this_vga_signals.N_417_cascade_ ;
    wire \this_vga_signals.N_412_cascade_ ;
    wire \this_vga_signals.N_390_0_cascade_ ;
    wire \this_vga_signals.N_390_0 ;
    wire \this_vga_signals.M_hstate_qZ0Z_2 ;
    wire \this_vga_signals.N_413_cascade_ ;
    wire \this_vga_signals.N_398_0 ;
    wire \this_vga_signals.M_hstate_qZ0Z_3 ;
    wire \this_vga_signals.M_hstate_q_srsts_0_a3_0_4 ;
    wire \this_vga_signals.N_416 ;
    wire \this_vga_signals.M_hstate_q_srsts_0_a3_0_4_cascade_ ;
    wire \this_vga_signals.M_hstate_qZ0Z_4 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_12 ;
    wire \this_vga_signals.M_hstate_d_0_sqmuxa_cascade_ ;
    wire \this_vga_signals.N_405_0 ;
    wire \this_vga_signals.M_hstate_qZ0Z_0 ;
    wire \this_vga_signals.N_405_0_cascade_ ;
    wire \this_vga_signals.N_409 ;
    wire \this_vga_signals.N_397_0 ;
    wire \this_vga_signals.M_hstate_qZ0Z_5 ;
    wire \this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5_cascade_ ;
    wire \this_vga_signals.N_385_0 ;
    wire \this_vga_signals.N_385_0_cascade_ ;
    wire \this_vga_signals.N_391_0 ;
    wire \this_vga_signals.N_386_0 ;
    wire \this_vga_signals.N_386_0_cascade_ ;
    wire \this_vga_signals.M_hstate_q_srsts_0_o3_2_1 ;
    wire \this_vga_signals.N_388_0 ;
    wire \this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5 ;
    wire \this_vga_signals.N_393_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire \this_vga_signals.g2_2_cascade_ ;
    wire \this_vga_signals.g1_cascade_ ;
    wire \this_vga_signals.g2_5_cascade_ ;
    wire \this_vga_signals.g1_1_4 ;
    wire \this_vga_signals.g0_14_N_8L16_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_c3_0_0_cascade_ ;
    wire this_vga_signals_un14_address_if_generate_plus_mult1_un75_sum_i_3;
    wire \this_vga_signals.if_N_2_6_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c3_0 ;
    wire \this_vga_signals.g0_14_N_7L14 ;
    wire \this_vga_signals.if_N_9_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb1 ;
    wire \this_vga_signals.mult1_un61_sum_axb1_cascade_ ;
    wire \this_vga_signals.if_m3_1_2_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_3_out ;
    wire \this_vga_signals.if_i2_mux_0 ;
    wire \this_vga_signals.if_N_6_0_0_cascade_ ;
    wire this_vga_signals_un6_address_if_generate_plus_mult1_un75_sum_i_3;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_13 ;
    wire \this_vga_signals.mult1_un40_sum_0_ac0_3_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_0_ac0_3_0_a1_0_cascade_ ;
    wire \this_vga_signals.if_m3_0_0 ;
    wire \this_vga_signals.mult1_un40_sum_0_ac0_3_1 ;
    wire \this_vga_signals.mult1_un40_sum_0_ac0_3_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_0_ac0_3_2 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_14 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_15 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire bfn_17_17_0_;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire bfn_17_18_0_;
    wire \this_vga_signals.M_hcounter_qZ0Z_10 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_9 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_10 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_11 ;
    wire \this_vga_signals.g1_1_1 ;
    wire \this_vga_signals.g2_1_0_cascade_ ;
    wire \this_vga_signals.g2_3_0_cascade_ ;
    wire \this_vga_signals.if_N_2_4_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c3_2_cascade_ ;
    wire \this_vga_signals.g0_0_6_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3 ;
    wire \this_vga_signals.g0_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb2_i ;
    wire \this_vga_signals.g0_14_N_4L6 ;
    wire \this_vga_signals.g1_2_1 ;
    wire \this_vga_signals.g2_5_0 ;
    wire \this_vga_signals.M_vaddress_q_RNI85LKP4Z0Z_2 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c3_1_1_0_cascade_ ;
    wire \this_vga_signals.g3_0_0_0_1_cascade_ ;
    wire \this_vga_signals.g1_2 ;
    wire \this_vga_signals.g2 ;
    wire \this_vga_signals.g1_0_1_0_0 ;
    wire \this_vga_signals.N_4_i ;
    wire \this_vga_signals.g0_14_N_7L14_1 ;
    wire \this_vga_signals.if_m2_0_1 ;
    wire \this_vga_signals.if_N_3_0_i ;
    wire \this_vga_signals.if_N_3_0_i_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_c3_0 ;
    wire \this_vga_signals.if_i1_mux_0 ;
    wire \this_vga_signals.if_m2 ;
    wire \this_vga_signals.M_haddress_q_RNILVKM8Z0Z_6_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_cascade_ ;
    wire \this_vga_signals.if_N_8_i ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_3_1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_1_0_cascade_ ;
    wire \this_vga_signals.if_N_4_i ;
    wire this_vga_signals_un6_address_if_N_5_mux_0_cascade_;
    wire \this_vga_signals.mult1_un47_sum_c3_cascade_ ;
    wire \this_vga_signals.if_m1_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_ ;
    wire \this_vga_signals.if_m1_9_1 ;
    wire \this_vga_signals.M_hstate_qZ0Z_1 ;
    wire \this_vga_signals.M_haddress_qZ0Z_0 ;
    wire bfn_18_15_0_;
    wire \this_vga_signals.M_haddress_qZ0Z_1 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_0 ;
    wire \this_vga_signals.M_haddress_qZ0Z_2 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_1 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_2 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_3 ;
    wire \this_vga_signals.M_haddress_qZ0Z_5 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_4 ;
    wire \this_vga_signals.M_haddress_qZ0Z_6 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_5 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_6 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_7 ;
    wire bfn_18_16_0_;
    wire \this_vga_signals.un1_M_haddress_q_cry_8 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_9 ;
    wire \this_vga_signals.un1_M_haddress_q_cry_10 ;
    wire \this_vga_signals.M_hstate_q_RNIFIH84Z0Z_5 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_16 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_17 ;
    wire \this_vga_signals.mult1_un54_sum_c3 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_0_i ;
    wire this_vga_signals_un6_address_if_generate_plus_mult1_un54_sum_i_3;
    wire \this_vga_signals.g1_3_1_cascade_ ;
    wire \this_vga_signals.if_N_7_cascade_ ;
    wire \this_vga_signals.if_m1_3 ;
    wire \this_vga_signals.if_m1_3_cascade_ ;
    wire \this_vga_signals.if_m8_am_cascade_ ;
    wire \this_vga_signals.if_m8_bm ;
    wire \this_vga_signals.g1_0_0 ;
    wire \this_vga_signals.g0_0_2_cascade_ ;
    wire \this_vga_signals.g0_0_3_0 ;
    wire \this_vga_signals.g3_2 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_0_0_1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_cascade_ ;
    wire \this_vga_signals.if_m1 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_2 ;
    wire \this_vga_signals.g1_N_2L1 ;
    wire \this_vga_signals.G_5_0_x2_1 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_cascade_ ;
    wire \this_vga_signals.g2_4_cascade_ ;
    wire \this_vga_signals.g1_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_1 ;
    wire \this_vga_signals.g0_0_0_2 ;
    wire \this_vga_signals.g0_29_1 ;
    wire \this_vga_signals.N_3_0_0_0 ;
    wire \this_vga_signals.if_N_7 ;
    wire \this_vga_signals.mult1_un54_sum_axb1 ;
    wire \this_vga_signals.mult1_un40_sum_m_2 ;
    wire this_vga_signals_un6_address_if_N_5_mux_0;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_c3 ;
    wire this_vga_signals_un6_address_if_generate_plus_mult1_un47_sum_i_3;
    wire \this_vga_signals.mult1_un40_sum_m_1 ;
    wire \this_vga_signals.CO1_1_0 ;
    wire \this_vga_signals.mult1_un40_sum_1_axb1 ;
    wire \this_vga_signals.mult1_un40_sum_1_c2_0 ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc2_0 ;
    wire \this_vga_signals.N_2_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_a4_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_0 ;
    wire \this_vga_signals.mult1_un40_sum1_0_3 ;
    wire \this_vga_signals.M_haddress_qZ0Z_7 ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_a5 ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_1 ;
    wire \this_vga_signals.mult1_un40_sum_1_ac0_2 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_15 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_18 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_16 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_17 ;
    wire M_state_qZ0Z_5;
    wire \this_start_data_delay.this_edge_detector.N_252_0 ;
    wire \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0 ;
    wire \this_start_data_delay.this_edge_detector.N_252_0_cascade_ ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_18 ;
    wire \this_start_data_delay.this_edge_detector.N_267_cascade_ ;
    wire \this_vga_signals.if_m12_bm ;
    wire \this_vga_signals.if_m12_am ;
    wire \this_vga_signals.if_m13_ns_1 ;
    wire if_m13_ns;
    wire \this_vga_signals.N_9_0_0_cascade_ ;
    wire \this_vga_signals.g0_4_2 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_0_0_1_1 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_d_cascade_ ;
    wire \this_vga_signals.if_N_2_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_2_cascade_ ;
    wire \this_vga_signals.N_3_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_1_x ;
    wire \this_vga_signals.g0_3_0_cascade_ ;
    wire \this_vga_signals.if_N_2_5 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_ ;
    wire \this_vga_signals.g0_0_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_0 ;
    wire \this_vga_signals.g0_0_5_1_cascade_ ;
    wire \this_vga_signals.g0_3_1 ;
    wire \this_vga_signals.if_N_2_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_0_0 ;
    wire M_this_vram_read_data_3;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0 ;
    wire \this_start_data_delay.this_edge_detector.N_253_0 ;
    wire \this_vga_signals.M_haddress_qZ0Z_3 ;
    wire \this_start_data_delay.this_edge_detector.N_261_cascade_ ;
    wire \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0Z0Z_0 ;
    wire M_this_start_address_delay_out_0;
    wire \this_start_data_delay.this_edge_detector.N_267 ;
    wire \this_start_data_delay.this_edge_detector.N_275_cascade_ ;
    wire \this_start_data_delay.this_edge_detector.N_263_cascade_ ;
    wire M_state_qZ0Z_0;
    wire port_address_c_0;
    wire port_address_c_1;
    wire \this_start_data_delay.this_edge_detector.N_275 ;
    wire \this_start_data_delay.this_edge_detector.N_259_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un68_sum_i_1_3 ;
    wire \this_vga_signals.M_haddress_qZ0Z_4 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_2 ;
    wire this_vga_signals_un6_address_if_generate_plus_mult1_un68_sum_i_3;
    wire \this_vga_signals.g0_14_N_8L16_sx ;
    wire \this_vga_signals.mult1_un40_sum1_3_cascade_ ;
    wire \this_vga_signals.g0_4_0 ;
    wire M_this_vram_read_data_1;
    wire \this_vga_signals.g0_1_1_1_cascade_ ;
    wire \this_vga_signals.g0_3_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_1_1 ;
    wire \this_vga_signals.N_2_1_0 ;
    wire \this_vga_signals.g0_3_2_1 ;
    wire \this_vga_signals.mult1_un40_sum_m_am_x_2_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_m_ns_2 ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_5_3 ;
    wire \this_vga_signals.mult1_un40_sum_m_x1_3_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_m_ns_3_cascade_ ;
    wire \this_vga_signals.N_6_i ;
    wire \this_vga_signals.mult1_un40_sum_m_am_2 ;
    wire \this_vga_signals.mult1_un40_sum1_3 ;
    wire \this_vga_signals.N_6_i_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0 ;
    wire \this_vga_signals.if_m5_0_s ;
    wire \this_vga_signals.if_m1_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ;
    wire \this_vga_signals.if_N_2_2_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1_3 ;
    wire \this_vga_signals.mult1_un61_sum_c3_1_0 ;
    wire M_state_qZ0Z_2;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_d ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_1 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_0 ;
    wire this_vga_signals_un14_address_if_generate_plus_mult1_un54_sum_i_3;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_5_4 ;
    wire \this_vga_signals.M_vaddress_q_fastZ0Z_7 ;
    wire \this_vga_signals.mult1_un40_sum_0_axb1 ;
    wire \this_vga_signals.mult1_un40_sum_m_1_1 ;
    wire \this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_m_0_1 ;
    wire \this_vga_signals.M_vaddress_q_fastZ0Z_6 ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_5_2_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_5_2 ;
    wire \this_vga_signals.mult1_un40_sum_1_axbxc3_a4_1_0 ;
    wire \this_vga_signals.M_vaddress_q_fastZ0Z_5 ;
    wire \this_vga_signals.M_vaddress_q_fastZ0Z_9 ;
    wire \this_vga_signals.M_vaddress_q_fastZ0Z_8 ;
    wire \this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8 ;
    wire \this_vga_signals.N_353_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_m_bm_2 ;
    wire \this_vga_signals.mult1_un40_sum_0_axbxc3_5_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_0_axbxc3_5_3 ;
    wire \this_vga_signals.mult1_un40_sum0_3 ;
    wire \this_vga_signals.M_vaddress_q_5_repZ0Z1 ;
    wire \this_vga_signals.N_9_0 ;
    wire \this_vga_signals.M_vaddress_q_6_repZ0Z1 ;
    wire \this_vga_signals.M_vaddress_q_7_repZ0Z1 ;
    wire \this_vga_signals.N_15_0 ;
    wire \this_vga_signals.N_15_0_0_cascade_ ;
    wire \this_vga_signals.M_haddress_qZ0Z_9 ;
    wire \this_vga_signals.M_haddress_qZ0Z_8 ;
    wire \this_vga_signals.M_haddress_qZ0Z_10 ;
    wire \this_vga_signals.CO0_0 ;
    wire M_haddress_q_RNI8ARU_11;
    wire M_state_qZ0Z_1;
    wire port_enb_c;
    wire M_state_qZ0Z_3;
    wire M_this_start_data_delay_out_0;
    wire \this_vram.mem_WE_2 ;
    wire port_address_c_5;
    wire port_address_c_2;
    wire port_address_c_6;
    wire \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3Z0Z_0 ;
    wire M_current_data_qZ0Z_1;
    wire \this_vga_signals.M_hstate_d_0_sqmuxa ;
    wire \this_vga_signals.M_vaddress_qZ0Z_0 ;
    wire bfn_23_9_0_;
    wire \this_vga_signals.M_vaddress_qZ0Z_1 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_0 ;
    wire \this_vga_signals.M_vaddress_qZ0Z_2 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_1 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_2 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_3 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_4 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNEZ0 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_5 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOEZ0 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_6 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_7 ;
    wire bfn_23_10_0_;
    wire \this_vga_signals.un1_M_vaddress_q_cry_8 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01REZ0 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPEZ0 ;
    wire \this_vga_signals.M_vaddress_qZ0Z_3 ;
    wire \this_vga_signals.N_1253_0_cascade_ ;
    wire \this_vga_signals.g1_1_cascade_ ;
    wire \this_vga_signals.N_15_0_0 ;
    wire \this_vga_signals.N_353_0 ;
    wire \this_vga_signals.N_3520_0_cascade_ ;
    wire \this_vga_signals.CO1_2_1 ;
    wire \this_vga_signals.mult1_un40_sum_0_2 ;
    wire \this_vga_signals.g0_1_N_2L1 ;
    wire \this_vga_signals.N_1253_0 ;
    wire \this_vga_signals.mult1_un40_sum_0_2_cascade_ ;
    wire \this_vga_signals.N_3_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_0_0 ;
    wire \this_vga_signals.g0_1_N_5L7_x0_cascade_ ;
    wire \this_vga_signals.g0_1_N_5L7_x1 ;
    wire \this_vga_signals.mult1_un40_sum_m_ns_3 ;
    wire \this_vga_signals.M_vaddress_qZ0Z_4 ;
    wire \this_vga_signals.g0_1_N_5L7_ns_cascade_ ;
    wire \this_vga_signals.g0_1_1_0 ;
    wire \this_vga_signals.N_355_0 ;
    wire \this_vga_signals.g1_4 ;
    wire \this_vga_signals.M_vaddress_qZ0Z_7 ;
    wire \this_vga_signals.M_vaddress_qZ0Z_8 ;
    wire \this_vga_signals.M_vaddress_qZ0Z_6 ;
    wire \this_vga_signals.CO0 ;
    wire \this_vga_signals.if_i2_mux ;
    wire M_this_vram_read_data_2;
    wire \this_vram.mem_WE_6 ;
    wire M_current_address_qZ1Z_0;
    wire M_current_address_qZ0Z_0;
    wire \this_vram.mem_out_bus5_0 ;
    wire \this_vram.mem_out_bus1_0 ;
    wire \this_vram.mem_mem_1_0_RNISSKZ0Z11 ;
    wire \this_vram.mem_radregZ0Z_11 ;
    wire \this_vram.mem_N_109_cascade_ ;
    wire M_this_vram_read_data_0;
    wire \this_vram.mem_out_bus0_0 ;
    wire \this_vram.mem_out_bus4_0 ;
    wire \this_vram.mem_mem_0_0_RNIQOIZ0Z11_cascade_ ;
    wire \this_vram.mem_N_112 ;
    wire \this_vram.mem_out_bus2_0 ;
    wire \this_vram.mem_out_bus6_0 ;
    wire \this_vram.mem_mem_2_0_RNIU0NZ0Z11 ;
    wire \this_vram.mem_out_bus1_1 ;
    wire \this_vram.mem_out_bus5_1 ;
    wire \this_vram.mem_mem_1_0_RNISSK11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_88 ;
    wire \this_vram.mem_out_bus4_2 ;
    wire \this_vram.mem_out_bus0_2 ;
    wire \this_vram.mem_out_bus6_2 ;
    wire \this_vram.mem_out_bus2_2 ;
    wire \this_vram.mem_mem_0_1_RNISOIZ0Z11 ;
    wire \this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_ ;
    wire \this_vram.mem_N_98 ;
    wire \this_vram.mem_out_bus6_1 ;
    wire \this_vram.mem_out_bus2_1 ;
    wire \this_vram.mem_out_bus4_1 ;
    wire \this_vram.mem_out_bus0_1 ;
    wire \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_ ;
    wire \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0 ;
    wire \this_vram.mem_N_91 ;
    wire \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKMEZ0 ;
    wire \this_vga_signals.M_vaddress_qZ0Z_5 ;
    wire \this_vga_signals.N_583_g ;
    wire \this_vram.mem_out_bus6_3 ;
    wire \this_vram.mem_out_bus2_3 ;
    wire \this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_105 ;
    wire \this_vram.mem_out_bus0_3 ;
    wire \this_vram.mem_out_bus4_3 ;
    wire \this_vram.mem_mem_0_1_RNISOI11Z0Z_0 ;
    wire \this_vram.mem_WE_12 ;
    wire \this_vram.mem_out_bus7_1 ;
    wire \this_vram.mem_out_bus3_1 ;
    wire \this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ;
    wire \this_vram.mem_out_bus5_3 ;
    wire \this_vram.mem_out_bus1_3 ;
    wire \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_102 ;
    wire \this_vram.mem_out_bus1_2 ;
    wire \this_vram.mem_out_bus5_2 ;
    wire \this_vram.mem_radregZ0Z_12 ;
    wire \this_vram.mem_mem_1_1_RNIUSKZ0Z11_cascade_ ;
    wire \this_vram.mem_N_95 ;
    wire \this_vram.mem_out_bus3_0 ;
    wire \this_vram.mem_out_bus7_0 ;
    wire \this_vram.mem_mem_3_0_RNI05PZ0Z11 ;
    wire \this_vram.mem_WE_10 ;
    wire \this_vram.mem_WE_8 ;
    wire \this_vram.mem_WE_14 ;
    wire \this_vram.mem_out_bus7_3 ;
    wire \this_vram.mem_out_bus3_3 ;
    wire \this_vram.mem_mem_3_1_RNI25P11Z0Z_0 ;
    wire \this_vram.mem_out_bus3_2 ;
    wire \this_vram.mem_out_bus7_2 ;
    wire \this_vram.mem_radregZ0Z_13 ;
    wire \this_vram.mem_mem_3_1_RNI25PZ0Z11 ;
    wire port_data_c_6;
    wire M_current_address_qZ0Z_6;
    wire \this_vram.mem_WE_4 ;
    wire M_current_address_qZ0Z_12;
    wire M_current_address_qZ0Z_13;
    wire debug_c;
    wire \this_vram.mem_WE_0 ;
    wire port_data_c_5;
    wire M_current_address_qZ0Z_5;
    wire M_current_address_qZ0Z_11;
    wire port_data_c_4;
    wire M_current_address_qZ0Z_4;
    wire M_current_address_qZ0Z_2;
    wire M_current_address_qZ0Z_9;
    wire M_current_data_qZ0Z_0;
    wire M_current_address_qZ0Z_1;
    wire M_current_address_qZ0Z_3;
    wire M_current_address_q_0_0;
    wire M_current_address_qZ0Z_10;
    wire port_data_c_0;
    wire M_current_address_qZ0Z_7;
    wire port_data_c_1;
    wire M_current_address_qZ0Z_8;
    wire M_current_address_q_0_6_0;
    wire N_631_g;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_2 ;
    wire \this_vga_signals.mult1_un61_sum_c3 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_0 ;
    wire this_vga_signals_un14_address_if_generate_plus_mult1_un61_sum_i_3;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_i ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3 ;
    wire this_vga_signals_un6_address_if_generate_plus_mult1_un61_sum_i_3;
    wire port_data_c_2;
    wire M_current_data_qZ0Z_2;
    wire M_current_data_d_0_sqmuxa;
    wire port_data_c_3;
    wire M_this_reset_cond_out_0;
    wire M_current_data_qZ0Z_3;
    wire clk_c_g;
    wire port_address_c_4;
    wire port_address_c_7;
    wire port_address_c_3;
    wire port_rw_c;
    wire \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4Z0Z_0 ;
    wire _gnd_net_;

    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,\this_vram.mem_out_bus0_1 ,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,\this_vram.mem_out_bus0_0 ,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__12194,N__17591,N__11120,N__9092,N__13331,N__10685,N__10502,N__10151,N__19829,N__11618,N__9221}),
            .WADDR({N__18278,N__18722,N__17987,N__18137,N__17474,N__17084,N__16889,N__18431,N__18830,N__18536,N__15770}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,N__14210,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__18614,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .RCLKE(),
            .RCLK(N__19111),
            .RE(N__7404),
            .WCLKE(N__16601),
            .WCLK(N__19112),
            .WE(N__7314));
    defparam \this_vram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,\this_vram.mem_out_bus0_3 ,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,\this_vram.mem_out_bus0_2 ,dangling_wire_55,dangling_wire_56,dangling_wire_57}),
            .RADDR({N__12188,N__17585,N__11114,N__9086,N__13325,N__10679,N__10496,N__10145,N__19823,N__11612,N__9215}),
            .WADDR({N__18272,N__18716,N__17981,N__18131,N__17468,N__17078,N__16883,N__18425,N__18824,N__18530,N__15764}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,N__19280,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,N__19697,dangling_wire_85,dangling_wire_86,dangling_wire_87}),
            .RCLKE(),
            .RCLK(N__19114),
            .RE(N__7385),
            .WCLKE(N__16597),
            .WCLK(N__19115),
            .WE(N__7389));
    defparam \this_vram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,\this_vram.mem_out_bus1_1 ,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,\this_vram.mem_out_bus1_0 ,dangling_wire_99,dangling_wire_100,dangling_wire_101}),
            .RADDR({N__12182,N__17579,N__11108,N__9080,N__13319,N__10673,N__10490,N__10139,N__19817,N__11606,N__9209}),
            .WADDR({N__18266,N__18710,N__17975,N__18125,N__17462,N__17072,N__16877,N__18419,N__18818,N__18524,N__15758}),
            .MASK({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .WDATA({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__14206,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__18610,dangling_wire_129,dangling_wire_130,dangling_wire_131}),
            .RCLKE(),
            .RCLK(N__19119),
            .RE(N__7384),
            .WCLKE(N__16142),
            .WCLK(N__19120),
            .WE(N__7255));
    defparam \this_vram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,\this_vram.mem_out_bus1_3 ,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,\this_vram.mem_out_bus1_2 ,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .RADDR({N__12176,N__17573,N__11102,N__9074,N__13313,N__10667,N__10484,N__10133,N__19811,N__11600,N__9203}),
            .WADDR({N__18260,N__18704,N__17969,N__18119,N__17456,N__17066,N__16871,N__18413,N__18812,N__18518,N__15752}),
            .MASK({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161}),
            .WDATA({dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__19276,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,N__19693,dangling_wire_173,dangling_wire_174,dangling_wire_175}),
            .RCLKE(),
            .RCLK(N__19130),
            .RE(N__7360),
            .WCLKE(N__16138),
            .WCLK(N__19131),
            .WE(N__7421));
    defparam \this_vram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,\this_vram.mem_out_bus2_1 ,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,\this_vram.mem_out_bus2_0 ,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .RADDR({N__12170,N__17567,N__11096,N__9068,N__13307,N__10661,N__10478,N__10127,N__19805,N__11594,N__9197}),
            .WADDR({N__18254,N__18698,N__17963,N__18113,N__17450,N__17060,N__16865,N__18407,N__18806,N__18512,N__15746}),
            .MASK({dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205}),
            .WDATA({dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,N__14199,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,N__18603,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .RCLKE(),
            .RCLK(N__19145),
            .RE(N__7359),
            .WCLKE(N__16640),
            .WCLK(N__19144),
            .WE(N__7417));
    defparam \this_vram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,\this_vram.mem_out_bus2_3 ,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,\this_vram.mem_out_bus2_2 ,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .RADDR({N__12164,N__17561,N__11090,N__9062,N__13301,N__10655,N__10472,N__10121,N__19799,N__11588,N__9191}),
            .WADDR({N__18248,N__18692,N__17957,N__18107,N__17444,N__17054,N__16859,N__18401,N__18800,N__18506,N__15740}),
            .MASK({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .WDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,N__19269,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,N__19686,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RCLKE(),
            .RCLK(N__19158),
            .RE(N__7332),
            .WCLKE(N__16636),
            .WCLK(N__19159),
            .WE(N__7416));
    defparam \this_vram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,\this_vram.mem_out_bus3_1 ,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,\this_vram.mem_out_bus3_0 ,dangling_wire_275,dangling_wire_276,dangling_wire_277}),
            .RADDR({N__12158,N__17555,N__11084,N__9056,N__13295,N__10649,N__10466,N__10115,N__19793,N__11582,N__9185}),
            .WADDR({N__18242,N__18686,N__17951,N__18101,N__17438,N__17048,N__16853,N__18395,N__18794,N__18500,N__15734}),
            .MASK({dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293}),
            .WDATA({dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,N__14189,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,N__18594,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .RCLKE(),
            .RCLK(N__19166),
            .RE(N__7331),
            .WCLKE(N__16612),
            .WCLK(N__19167),
            .WE(N__7406));
    defparam \this_vram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,\this_vram.mem_out_bus3_3 ,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,\this_vram.mem_out_bus3_2 ,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .RADDR({N__12152,N__17549,N__11078,N__9050,N__13289,N__10643,N__10460,N__10109,N__19787,N__11576,N__9179}),
            .WADDR({N__18236,N__18680,N__17945,N__18095,N__17432,N__17042,N__16847,N__18389,N__18788,N__18494,N__15728}),
            .MASK({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .WDATA({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,N__19260,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,N__19676,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .RCLKE(),
            .RCLK(N__19170),
            .RE(N__7298),
            .WCLKE(N__16619),
            .WCLK(N__19171),
            .WE(N__7405));
    defparam \this_vram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,\this_vram.mem_out_bus4_1 ,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,\this_vram.mem_out_bus4_0 ,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .RADDR({N__12146,N__17543,N__11072,N__9044,N__13283,N__10637,N__10454,N__10103,N__19781,N__11570,N__9173}),
            .WADDR({N__18230,N__18674,N__17939,N__18089,N__17426,N__17036,N__16841,N__18383,N__18782,N__18488,N__15722}),
            .MASK({dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381}),
            .WDATA({dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,N__14177,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,N__18585,dangling_wire_393,dangling_wire_394,dangling_wire_395}),
            .RCLKE(),
            .RCLK(N__19173),
            .RE(N__7390),
            .WCLKE(N__15799),
            .WCLK(N__19174),
            .WE(N__7209));
    defparam \this_vram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,\this_vram.mem_out_bus4_3 ,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,\this_vram.mem_out_bus4_2 ,dangling_wire_407,dangling_wire_408,dangling_wire_409}),
            .RADDR({N__12140,N__17537,N__11066,N__9038,N__13277,N__10631,N__10448,N__10097,N__19775,N__11564,N__9167}),
            .WADDR({N__18224,N__18668,N__17933,N__18083,N__17420,N__17030,N__16835,N__18377,N__18776,N__18482,N__15716}),
            .MASK({dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425}),
            .WDATA({dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,N__19251,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,N__19675,dangling_wire_437,dangling_wire_438,dangling_wire_439}),
            .RCLKE(),
            .RCLK(N__19176),
            .RE(N__7349),
            .WCLKE(N__15800),
            .WCLK(N__19177),
            .WE(N__7373));
    defparam \this_vram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,\this_vram.mem_out_bus5_1 ,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,\this_vram.mem_out_bus5_0 ,dangling_wire_451,dangling_wire_452,dangling_wire_453}),
            .RADDR({N__12134,N__17531,N__11060,N__9032,N__13271,N__10625,N__10442,N__10091,N__19769,N__11558,N__9161}),
            .WADDR({N__18218,N__18662,N__17927,N__18077,N__17414,N__17024,N__16829,N__18371,N__18770,N__18476,N__15710}),
            .MASK({dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469}),
            .WDATA({dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,N__14165,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,N__18576,dangling_wire_481,dangling_wire_482,dangling_wire_483}),
            .RCLKE(),
            .RCLK(N__19180),
            .RE(N__7350),
            .WCLKE(N__17362),
            .WCLK(N__19181),
            .WE(N__7329));
    defparam \this_vram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,\this_vram.mem_out_bus5_3 ,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,\this_vram.mem_out_bus5_2 ,dangling_wire_495,dangling_wire_496,dangling_wire_497}),
            .RADDR({N__12128,N__17525,N__11054,N__9026,N__13265,N__10619,N__10436,N__10085,N__19763,N__11552,N__9155}),
            .WADDR({N__18212,N__18656,N__17921,N__18071,N__17408,N__17018,N__16823,N__18365,N__18764,N__18470,N__15704}),
            .MASK({dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513}),
            .WDATA({dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,N__19241,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,N__19640,dangling_wire_525,dangling_wire_526,dangling_wire_527}),
            .RCLKE(),
            .RCLK(N__19184),
            .RE(N__7316),
            .WCLKE(N__17366),
            .WCLK(N__19185),
            .WE(N__7320));
    defparam \this_vram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,\this_vram.mem_out_bus6_1 ,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,\this_vram.mem_out_bus6_0 ,dangling_wire_539,dangling_wire_540,dangling_wire_541}),
            .RADDR({N__12122,N__17519,N__11048,N__9020,N__13259,N__10613,N__10430,N__10079,N__19757,N__11546,N__9149}),
            .WADDR({N__18206,N__18650,N__17915,N__18065,N__17402,N__17012,N__16817,N__18359,N__18758,N__18464,N__15698}),
            .MASK({dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557}),
            .WDATA({dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,N__14153,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,N__18555,dangling_wire_569,dangling_wire_570,dangling_wire_571}),
            .RCLKE(),
            .RCLK(N__19190),
            .RE(N__7283),
            .WCLKE(N__14281),
            .WCLK(N__19191),
            .WE(N__7274));
    defparam \this_vram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,\this_vram.mem_out_bus6_3 ,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,\this_vram.mem_out_bus6_2 ,dangling_wire_583,dangling_wire_584,dangling_wire_585}),
            .RADDR({N__12116,N__17513,N__11042,N__9014,N__13253,N__10607,N__10424,N__10073,N__19751,N__11540,N__9143}),
            .WADDR({N__18200,N__18644,N__17909,N__18059,N__17396,N__17006,N__16811,N__18353,N__18752,N__18458,N__15692}),
            .MASK({dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601}),
            .WDATA({dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,N__19221,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,N__19671,dangling_wire_613,dangling_wire_614,dangling_wire_615}),
            .RCLKE(),
            .RCLK(N__19195),
            .RE(N__7315),
            .WCLKE(N__14285),
            .WCLK(N__19196),
            .WE(N__7273));
    defparam \this_vram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,\this_vram.mem_out_bus7_1 ,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,\this_vram.mem_out_bus7_0 ,dangling_wire_627,dangling_wire_628,dangling_wire_629}),
            .RADDR({N__12110,N__17507,N__11036,N__9008,N__13247,N__10601,N__10418,N__10067,N__19745,N__11534,N__9137}),
            .WADDR({N__18194,N__18638,N__17903,N__18053,N__17390,N__17000,N__16805,N__18347,N__18746,N__18452,N__15686}),
            .MASK({dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645}),
            .WDATA({dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,N__14152,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,N__18575,dangling_wire_657,dangling_wire_658,dangling_wire_659}),
            .RCLKE(),
            .RCLK(N__19199),
            .RE(N__7218),
            .WCLKE(N__17128),
            .WCLK(N__19200),
            .WE(N__7269));
    defparam \this_vram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,\this_vram.mem_out_bus7_3 ,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,\this_vram.mem_out_bus7_2 ,dangling_wire_671,dangling_wire_672,dangling_wire_673}),
            .RADDR({N__12104,N__17501,N__11030,N__9002,N__13241,N__10595,N__10412,N__10061,N__19739,N__11528,N__9131}),
            .WADDR({N__18188,N__18632,N__17897,N__18047,N__17384,N__16994,N__16799,N__18341,N__18740,N__18446,N__15680}),
            .MASK({dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689}),
            .WDATA({dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,N__19250,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,N__19685,dangling_wire_701,dangling_wire_702,dangling_wire_703}),
            .RCLKE(),
            .RCLK(N__19201),
            .RE(N__7282),
            .WCLKE(N__17132),
            .WCLK(N__19202),
            .WE(N__7281));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__20238),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__20240),
            .DIN(N__20239),
            .DOUT(N__20238),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__20240),
            .PADOUT(N__20239),
            .PADIN(N__20238),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_iopad (
            .OE(N__20229),
            .DIN(N__20228),
            .DOUT(N__20227),
            .PACKAGEPIN(debug));
    defparam debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_preio (
            .PADOEN(N__20229),
            .PADOUT(N__20228),
            .PADIN(N__20227),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__17225),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__20220),
            .DIN(N__20219),
            .DOUT(N__20218),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__20220),
            .PADOUT(N__20219),
            .PADIN(N__20218),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7556),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__20211),
            .DIN(N__20210),
            .DOUT(N__20209),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__20211),
            .PADOUT(N__20210),
            .PADIN(N__20209),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7499),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_0_iopad (
            .OE(N__20202),
            .DIN(N__20201),
            .DOUT(N__20200),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_0_preio (
            .PADOEN(N__20202),
            .PADOUT(N__20201),
            .PADIN(N__20200),
            .CLOCKENABLE(),
            .DIN0(port_address_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_1_iopad (
            .OE(N__20193),
            .DIN(N__20192),
            .DOUT(N__20191),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_1_preio (
            .PADOEN(N__20193),
            .PADOUT(N__20192),
            .PADIN(N__20191),
            .CLOCKENABLE(),
            .DIN0(port_address_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_2_iopad (
            .OE(N__20184),
            .DIN(N__20183),
            .DOUT(N__20182),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_2_preio (
            .PADOEN(N__20184),
            .PADOUT(N__20183),
            .PADIN(N__20182),
            .CLOCKENABLE(),
            .DIN0(port_address_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_3_iopad (
            .OE(N__20175),
            .DIN(N__20174),
            .DOUT(N__20173),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_3_preio (
            .PADOEN(N__20175),
            .PADOUT(N__20174),
            .PADIN(N__20173),
            .CLOCKENABLE(),
            .DIN0(port_address_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_4_iopad (
            .OE(N__20166),
            .DIN(N__20165),
            .DOUT(N__20164),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_4_preio (
            .PADOEN(N__20166),
            .PADOUT(N__20165),
            .PADIN(N__20164),
            .CLOCKENABLE(),
            .DIN0(port_address_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_5_iopad (
            .OE(N__20157),
            .DIN(N__20156),
            .DOUT(N__20155),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_5_preio (
            .PADOEN(N__20157),
            .PADOUT(N__20156),
            .PADIN(N__20155),
            .CLOCKENABLE(),
            .DIN0(port_address_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_6_iopad (
            .OE(N__20148),
            .DIN(N__20147),
            .DOUT(N__20146),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_6_preio (
            .PADOEN(N__20148),
            .PADOUT(N__20147),
            .PADIN(N__20146),
            .CLOCKENABLE(),
            .DIN0(port_address_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_7_iopad (
            .OE(N__20139),
            .DIN(N__20138),
            .DOUT(N__20137),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_7_preio (
            .PADOEN(N__20139),
            .PADOUT(N__20138),
            .PADIN(N__20137),
            .CLOCKENABLE(),
            .DIN0(port_address_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__20130),
            .DIN(N__20129),
            .DOUT(N__20128),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__20130),
            .PADOUT(N__20129),
            .PADIN(N__20128),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__20121),
            .DIN(N__20120),
            .DOUT(N__20119),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__20121),
            .PADOUT(N__20120),
            .PADIN(N__20119),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__20112),
            .DIN(N__20111),
            .DOUT(N__20110),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__20112),
            .PADOUT(N__20111),
            .PADIN(N__20110),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__20103),
            .DIN(N__20102),
            .DOUT(N__20101),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__20103),
            .PADOUT(N__20102),
            .PADIN(N__20101),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__20094),
            .DIN(N__20093),
            .DOUT(N__20092),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__20094),
            .PADOUT(N__20093),
            .PADIN(N__20092),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__20085),
            .DIN(N__20084),
            .DOUT(N__20083),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__20085),
            .PADOUT(N__20084),
            .PADIN(N__20083),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__20076),
            .DIN(N__20075),
            .DOUT(N__20074),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__20076),
            .PADOUT(N__20075),
            .PADIN(N__20074),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__20067),
            .DIN(N__20066),
            .DOUT(N__20065),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__20067),
            .PADOUT(N__20066),
            .PADIN(N__20065),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__20058),
            .DIN(N__20057),
            .DOUT(N__20056),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__20058),
            .PADOUT(N__20057),
            .PADIN(N__20056),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7427),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__20049),
            .DIN(N__20048),
            .DOUT(N__20047),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__20049),
            .PADOUT(N__20048),
            .PADIN(N__20047),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7330),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__20040),
            .DIN(N__20039),
            .DOUT(N__20038),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__20040),
            .PADOUT(N__20039),
            .PADIN(N__20038),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__20031),
            .DIN(N__20030),
            .DOUT(N__20029),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__20031),
            .PADOUT(N__20030),
            .PADIN(N__20029),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7910),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_ibuf_iopad (
            .OE(N__20022),
            .DIN(N__20021),
            .DOUT(N__20020),
            .PACKAGEPIN(port_rw));
    defparam port_rw_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_rw_ibuf_preio (
            .PADOEN(N__20022),
            .PADOUT(N__20021),
            .PADIN(N__20020),
            .CLOCKENABLE(),
            .DIN0(port_rw_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__20013),
            .DIN(N__20012),
            .DOUT(N__20011),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__20013),
            .PADOUT(N__20012),
            .PADIN(N__20011),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7469),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__20004),
            .DIN(N__20003),
            .DOUT(N__20002),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__20004),
            .PADOUT(N__20003),
            .PADIN(N__20002),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7439),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__19995),
            .DIN(N__19994),
            .DOUT(N__19993),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__19995),
            .PADOUT(N__19994),
            .PADIN(N__19993),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7526),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__19986),
            .DIN(N__19985),
            .DOUT(N__19984),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__19986),
            .PADOUT(N__19985),
            .PADIN(N__19984),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7580),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__19977),
            .DIN(N__19976),
            .DOUT(N__19975),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__19977),
            .PADOUT(N__19976),
            .PADIN(N__19975),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7481),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__19968),
            .DIN(N__19967),
            .DOUT(N__19966),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__19968),
            .PADOUT(N__19967),
            .PADIN(N__19966),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7517),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__19959),
            .DIN(N__19958),
            .DOUT(N__19957),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__19959),
            .PADOUT(N__19958),
            .PADIN(N__19957),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__19950),
            .DIN(N__19949),
            .DOUT(N__19948),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__19950),
            .PADOUT(N__19949),
            .PADIN(N__19948),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7538),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__19941),
            .DIN(N__19940),
            .DOUT(N__19939),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__19941),
            .PADOUT(N__19940),
            .PADIN(N__19939),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8126),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__4782 (
            .O(N__19922),
            .I(N__19919));
    LocalMux I__4781 (
            .O(N__19919),
            .I(N__19916));
    Span4Mux_v I__4780 (
            .O(N__19916),
            .I(N__19912));
    InMux I__4779 (
            .O(N__19915),
            .I(N__19909));
    Sp12to4 I__4778 (
            .O(N__19912),
            .I(N__19905));
    LocalMux I__4777 (
            .O(N__19909),
            .I(N__19901));
    InMux I__4776 (
            .O(N__19908),
            .I(N__19898));
    Span12Mux_v I__4775 (
            .O(N__19905),
            .I(N__19895));
    InMux I__4774 (
            .O(N__19904),
            .I(N__19892));
    Span4Mux_v I__4773 (
            .O(N__19901),
            .I(N__19887));
    LocalMux I__4772 (
            .O(N__19898),
            .I(N__19887));
    Odrv12 I__4771 (
            .O(N__19895),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    LocalMux I__4770 (
            .O(N__19892),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    Odrv4 I__4769 (
            .O(N__19887),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    InMux I__4768 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__4767 (
            .O(N__19877),
            .I(N__19874));
    Span4Mux_s3_v I__4766 (
            .O(N__19874),
            .I(N__19871));
    Span4Mux_h I__4765 (
            .O(N__19871),
            .I(N__19868));
    Span4Mux_v I__4764 (
            .O(N__19868),
            .I(N__19865));
    Span4Mux_v I__4763 (
            .O(N__19865),
            .I(N__19861));
    InMux I__4762 (
            .O(N__19864),
            .I(N__19858));
    Span4Mux_v I__4761 (
            .O(N__19861),
            .I(N__19853));
    LocalMux I__4760 (
            .O(N__19858),
            .I(N__19853));
    Span4Mux_v I__4759 (
            .O(N__19853),
            .I(N__19846));
    InMux I__4758 (
            .O(N__19852),
            .I(N__19839));
    InMux I__4757 (
            .O(N__19851),
            .I(N__19839));
    InMux I__4756 (
            .O(N__19850),
            .I(N__19839));
    InMux I__4755 (
            .O(N__19849),
            .I(N__19836));
    Odrv4 I__4754 (
            .O(N__19846),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    LocalMux I__4753 (
            .O(N__19839),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    LocalMux I__4752 (
            .O(N__19836),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    CascadeMux I__4751 (
            .O(N__19829),
            .I(N__19826));
    CascadeBuf I__4750 (
            .O(N__19826),
            .I(N__19823));
    CascadeMux I__4749 (
            .O(N__19823),
            .I(N__19820));
    CascadeBuf I__4748 (
            .O(N__19820),
            .I(N__19817));
    CascadeMux I__4747 (
            .O(N__19817),
            .I(N__19814));
    CascadeBuf I__4746 (
            .O(N__19814),
            .I(N__19811));
    CascadeMux I__4745 (
            .O(N__19811),
            .I(N__19808));
    CascadeBuf I__4744 (
            .O(N__19808),
            .I(N__19805));
    CascadeMux I__4743 (
            .O(N__19805),
            .I(N__19802));
    CascadeBuf I__4742 (
            .O(N__19802),
            .I(N__19799));
    CascadeMux I__4741 (
            .O(N__19799),
            .I(N__19796));
    CascadeBuf I__4740 (
            .O(N__19796),
            .I(N__19793));
    CascadeMux I__4739 (
            .O(N__19793),
            .I(N__19790));
    CascadeBuf I__4738 (
            .O(N__19790),
            .I(N__19787));
    CascadeMux I__4737 (
            .O(N__19787),
            .I(N__19784));
    CascadeBuf I__4736 (
            .O(N__19784),
            .I(N__19781));
    CascadeMux I__4735 (
            .O(N__19781),
            .I(N__19778));
    CascadeBuf I__4734 (
            .O(N__19778),
            .I(N__19775));
    CascadeMux I__4733 (
            .O(N__19775),
            .I(N__19772));
    CascadeBuf I__4732 (
            .O(N__19772),
            .I(N__19769));
    CascadeMux I__4731 (
            .O(N__19769),
            .I(N__19766));
    CascadeBuf I__4730 (
            .O(N__19766),
            .I(N__19763));
    CascadeMux I__4729 (
            .O(N__19763),
            .I(N__19760));
    CascadeBuf I__4728 (
            .O(N__19760),
            .I(N__19757));
    CascadeMux I__4727 (
            .O(N__19757),
            .I(N__19754));
    CascadeBuf I__4726 (
            .O(N__19754),
            .I(N__19751));
    CascadeMux I__4725 (
            .O(N__19751),
            .I(N__19748));
    CascadeBuf I__4724 (
            .O(N__19748),
            .I(N__19745));
    CascadeMux I__4723 (
            .O(N__19745),
            .I(N__19742));
    CascadeBuf I__4722 (
            .O(N__19742),
            .I(N__19739));
    CascadeMux I__4721 (
            .O(N__19739),
            .I(N__19736));
    InMux I__4720 (
            .O(N__19736),
            .I(N__19733));
    LocalMux I__4719 (
            .O(N__19733),
            .I(this_vga_signals_un6_address_if_generate_plus_mult1_un61_sum_i_3));
    InMux I__4718 (
            .O(N__19730),
            .I(N__19727));
    LocalMux I__4717 (
            .O(N__19727),
            .I(N__19724));
    Span4Mux_v I__4716 (
            .O(N__19724),
            .I(N__19719));
    InMux I__4715 (
            .O(N__19723),
            .I(N__19716));
    InMux I__4714 (
            .O(N__19722),
            .I(N__19713));
    Sp12to4 I__4713 (
            .O(N__19719),
            .I(N__19708));
    LocalMux I__4712 (
            .O(N__19716),
            .I(N__19708));
    LocalMux I__4711 (
            .O(N__19713),
            .I(N__19705));
    Span12Mux_h I__4710 (
            .O(N__19708),
            .I(N__19700));
    Sp12to4 I__4709 (
            .O(N__19705),
            .I(N__19700));
    Odrv12 I__4708 (
            .O(N__19700),
            .I(port_data_c_2));
    InMux I__4707 (
            .O(N__19697),
            .I(N__19694));
    LocalMux I__4706 (
            .O(N__19694),
            .I(N__19690));
    InMux I__4705 (
            .O(N__19693),
            .I(N__19687));
    Span4Mux_v I__4704 (
            .O(N__19690),
            .I(N__19680));
    LocalMux I__4703 (
            .O(N__19687),
            .I(N__19680));
    InMux I__4702 (
            .O(N__19686),
            .I(N__19677));
    InMux I__4701 (
            .O(N__19685),
            .I(N__19672));
    Span4Mux_v I__4700 (
            .O(N__19680),
            .I(N__19666));
    LocalMux I__4699 (
            .O(N__19677),
            .I(N__19666));
    InMux I__4698 (
            .O(N__19676),
            .I(N__19663));
    InMux I__4697 (
            .O(N__19675),
            .I(N__19660));
    LocalMux I__4696 (
            .O(N__19672),
            .I(N__19657));
    InMux I__4695 (
            .O(N__19671),
            .I(N__19654));
    Span4Mux_v I__4694 (
            .O(N__19666),
            .I(N__19649));
    LocalMux I__4693 (
            .O(N__19663),
            .I(N__19649));
    LocalMux I__4692 (
            .O(N__19660),
            .I(N__19646));
    Span4Mux_v I__4691 (
            .O(N__19657),
            .I(N__19641));
    LocalMux I__4690 (
            .O(N__19654),
            .I(N__19641));
    Sp12to4 I__4689 (
            .O(N__19649),
            .I(N__19636));
    Span4Mux_h I__4688 (
            .O(N__19646),
            .I(N__19633));
    Span4Mux_v I__4687 (
            .O(N__19641),
            .I(N__19630));
    InMux I__4686 (
            .O(N__19640),
            .I(N__19627));
    InMux I__4685 (
            .O(N__19639),
            .I(N__19624));
    Odrv12 I__4684 (
            .O(N__19636),
            .I(M_current_data_qZ0Z_2));
    Odrv4 I__4683 (
            .O(N__19633),
            .I(M_current_data_qZ0Z_2));
    Odrv4 I__4682 (
            .O(N__19630),
            .I(M_current_data_qZ0Z_2));
    LocalMux I__4681 (
            .O(N__19627),
            .I(M_current_data_qZ0Z_2));
    LocalMux I__4680 (
            .O(N__19624),
            .I(M_current_data_qZ0Z_2));
    InMux I__4679 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__4678 (
            .O(N__19610),
            .I(N__19605));
    InMux I__4677 (
            .O(N__19609),
            .I(N__19602));
    InMux I__4676 (
            .O(N__19608),
            .I(N__19598));
    Span4Mux_v I__4675 (
            .O(N__19605),
            .I(N__19593));
    LocalMux I__4674 (
            .O(N__19602),
            .I(N__19593));
    InMux I__4673 (
            .O(N__19601),
            .I(N__19590));
    LocalMux I__4672 (
            .O(N__19598),
            .I(N__19587));
    Span4Mux_h I__4671 (
            .O(N__19593),
            .I(N__19584));
    LocalMux I__4670 (
            .O(N__19590),
            .I(N__19581));
    Span12Mux_s10_h I__4669 (
            .O(N__19587),
            .I(N__19574));
    Sp12to4 I__4668 (
            .O(N__19584),
            .I(N__19574));
    Span12Mux_s5_v I__4667 (
            .O(N__19581),
            .I(N__19574));
    Odrv12 I__4666 (
            .O(N__19574),
            .I(M_current_data_d_0_sqmuxa));
    InMux I__4665 (
            .O(N__19571),
            .I(N__19567));
    CascadeMux I__4664 (
            .O(N__19570),
            .I(N__19563));
    LocalMux I__4663 (
            .O(N__19567),
            .I(N__19560));
    InMux I__4662 (
            .O(N__19566),
            .I(N__19557));
    InMux I__4661 (
            .O(N__19563),
            .I(N__19554));
    Span4Mux_v I__4660 (
            .O(N__19560),
            .I(N__19551));
    LocalMux I__4659 (
            .O(N__19557),
            .I(N__19546));
    LocalMux I__4658 (
            .O(N__19554),
            .I(N__19546));
    Span4Mux_h I__4657 (
            .O(N__19551),
            .I(N__19543));
    Span12Mux_h I__4656 (
            .O(N__19546),
            .I(N__19540));
    Odrv4 I__4655 (
            .O(N__19543),
            .I(port_data_c_3));
    Odrv12 I__4654 (
            .O(N__19540),
            .I(port_data_c_3));
    InMux I__4653 (
            .O(N__19535),
            .I(N__19524));
    InMux I__4652 (
            .O(N__19534),
            .I(N__19524));
    InMux I__4651 (
            .O(N__19533),
            .I(N__19524));
    InMux I__4650 (
            .O(N__19532),
            .I(N__19520));
    InMux I__4649 (
            .O(N__19531),
            .I(N__19515));
    LocalMux I__4648 (
            .O(N__19524),
            .I(N__19512));
    CascadeMux I__4647 (
            .O(N__19523),
            .I(N__19506));
    LocalMux I__4646 (
            .O(N__19520),
            .I(N__19501));
    InMux I__4645 (
            .O(N__19519),
            .I(N__19496));
    InMux I__4644 (
            .O(N__19518),
            .I(N__19496));
    LocalMux I__4643 (
            .O(N__19515),
            .I(N__19491));
    Span4Mux_v I__4642 (
            .O(N__19512),
            .I(N__19491));
    InMux I__4641 (
            .O(N__19511),
            .I(N__19488));
    IoInMux I__4640 (
            .O(N__19510),
            .I(N__19485));
    CascadeMux I__4639 (
            .O(N__19509),
            .I(N__19482));
    InMux I__4638 (
            .O(N__19506),
            .I(N__19465));
    InMux I__4637 (
            .O(N__19505),
            .I(N__19462));
    InMux I__4636 (
            .O(N__19504),
            .I(N__19459));
    Span4Mux_v I__4635 (
            .O(N__19501),
            .I(N__19456));
    LocalMux I__4634 (
            .O(N__19496),
            .I(N__19449));
    Span4Mux_h I__4633 (
            .O(N__19491),
            .I(N__19449));
    LocalMux I__4632 (
            .O(N__19488),
            .I(N__19449));
    LocalMux I__4631 (
            .O(N__19485),
            .I(N__19446));
    InMux I__4630 (
            .O(N__19482),
            .I(N__19442));
    InMux I__4629 (
            .O(N__19481),
            .I(N__19439));
    InMux I__4628 (
            .O(N__19480),
            .I(N__19434));
    InMux I__4627 (
            .O(N__19479),
            .I(N__19434));
    InMux I__4626 (
            .O(N__19478),
            .I(N__19429));
    InMux I__4625 (
            .O(N__19477),
            .I(N__19429));
    InMux I__4624 (
            .O(N__19476),
            .I(N__19426));
    InMux I__4623 (
            .O(N__19475),
            .I(N__19421));
    InMux I__4622 (
            .O(N__19474),
            .I(N__19421));
    InMux I__4621 (
            .O(N__19473),
            .I(N__19418));
    InMux I__4620 (
            .O(N__19472),
            .I(N__19415));
    InMux I__4619 (
            .O(N__19471),
            .I(N__19412));
    InMux I__4618 (
            .O(N__19470),
            .I(N__19407));
    InMux I__4617 (
            .O(N__19469),
            .I(N__19407));
    InMux I__4616 (
            .O(N__19468),
            .I(N__19404));
    LocalMux I__4615 (
            .O(N__19465),
            .I(N__19401));
    LocalMux I__4614 (
            .O(N__19462),
            .I(N__19398));
    LocalMux I__4613 (
            .O(N__19459),
            .I(N__19395));
    Span4Mux_h I__4612 (
            .O(N__19456),
            .I(N__19390));
    Span4Mux_v I__4611 (
            .O(N__19449),
            .I(N__19390));
    Span4Mux_s3_v I__4610 (
            .O(N__19446),
            .I(N__19387));
    InMux I__4609 (
            .O(N__19445),
            .I(N__19384));
    LocalMux I__4608 (
            .O(N__19442),
            .I(N__19379));
    LocalMux I__4607 (
            .O(N__19439),
            .I(N__19379));
    LocalMux I__4606 (
            .O(N__19434),
            .I(N__19370));
    LocalMux I__4605 (
            .O(N__19429),
            .I(N__19370));
    LocalMux I__4604 (
            .O(N__19426),
            .I(N__19363));
    LocalMux I__4603 (
            .O(N__19421),
            .I(N__19363));
    LocalMux I__4602 (
            .O(N__19418),
            .I(N__19363));
    LocalMux I__4601 (
            .O(N__19415),
            .I(N__19358));
    LocalMux I__4600 (
            .O(N__19412),
            .I(N__19358));
    LocalMux I__4599 (
            .O(N__19407),
            .I(N__19353));
    LocalMux I__4598 (
            .O(N__19404),
            .I(N__19353));
    Span4Mux_v I__4597 (
            .O(N__19401),
            .I(N__19346));
    Span4Mux_v I__4596 (
            .O(N__19398),
            .I(N__19346));
    Span4Mux_v I__4595 (
            .O(N__19395),
            .I(N__19346));
    Span4Mux_v I__4594 (
            .O(N__19390),
            .I(N__19341));
    Span4Mux_v I__4593 (
            .O(N__19387),
            .I(N__19341));
    LocalMux I__4592 (
            .O(N__19384),
            .I(N__19336));
    Span4Mux_v I__4591 (
            .O(N__19379),
            .I(N__19336));
    InMux I__4590 (
            .O(N__19378),
            .I(N__19327));
    InMux I__4589 (
            .O(N__19377),
            .I(N__19327));
    InMux I__4588 (
            .O(N__19376),
            .I(N__19327));
    InMux I__4587 (
            .O(N__19375),
            .I(N__19327));
    Span4Mux_h I__4586 (
            .O(N__19370),
            .I(N__19324));
    Span4Mux_h I__4585 (
            .O(N__19363),
            .I(N__19321));
    Span4Mux_h I__4584 (
            .O(N__19358),
            .I(N__19316));
    Span4Mux_h I__4583 (
            .O(N__19353),
            .I(N__19316));
    Sp12to4 I__4582 (
            .O(N__19346),
            .I(N__19311));
    Sp12to4 I__4581 (
            .O(N__19341),
            .I(N__19311));
    Span4Mux_h I__4580 (
            .O(N__19336),
            .I(N__19308));
    LocalMux I__4579 (
            .O(N__19327),
            .I(N__19303));
    Span4Mux_v I__4578 (
            .O(N__19324),
            .I(N__19303));
    Sp12to4 I__4577 (
            .O(N__19321),
            .I(N__19296));
    Sp12to4 I__4576 (
            .O(N__19316),
            .I(N__19296));
    Span12Mux_h I__4575 (
            .O(N__19311),
            .I(N__19296));
    Span4Mux_v I__4574 (
            .O(N__19308),
            .I(N__19293));
    Span4Mux_v I__4573 (
            .O(N__19303),
            .I(N__19290));
    Span12Mux_v I__4572 (
            .O(N__19296),
            .I(N__19287));
    Odrv4 I__4571 (
            .O(N__19293),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__4570 (
            .O(N__19290),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__4569 (
            .O(N__19287),
            .I(M_this_reset_cond_out_0));
    InMux I__4568 (
            .O(N__19280),
            .I(N__19277));
    LocalMux I__4567 (
            .O(N__19277),
            .I(N__19273));
    InMux I__4566 (
            .O(N__19276),
            .I(N__19270));
    Span4Mux_v I__4565 (
            .O(N__19273),
            .I(N__19264));
    LocalMux I__4564 (
            .O(N__19270),
            .I(N__19264));
    InMux I__4563 (
            .O(N__19269),
            .I(N__19261));
    Span4Mux_v I__4562 (
            .O(N__19264),
            .I(N__19255));
    LocalMux I__4561 (
            .O(N__19261),
            .I(N__19255));
    InMux I__4560 (
            .O(N__19260),
            .I(N__19252));
    Span4Mux_v I__4559 (
            .O(N__19255),
            .I(N__19245));
    LocalMux I__4558 (
            .O(N__19252),
            .I(N__19245));
    InMux I__4557 (
            .O(N__19251),
            .I(N__19242));
    InMux I__4556 (
            .O(N__19250),
            .I(N__19238));
    Span4Mux_v I__4555 (
            .O(N__19245),
            .I(N__19233));
    LocalMux I__4554 (
            .O(N__19242),
            .I(N__19233));
    InMux I__4553 (
            .O(N__19241),
            .I(N__19230));
    LocalMux I__4552 (
            .O(N__19238),
            .I(N__19227));
    Span4Mux_v I__4551 (
            .O(N__19233),
            .I(N__19222));
    LocalMux I__4550 (
            .O(N__19230),
            .I(N__19222));
    Span4Mux_s2_v I__4549 (
            .O(N__19227),
            .I(N__19215));
    Span4Mux_v I__4548 (
            .O(N__19222),
            .I(N__19215));
    InMux I__4547 (
            .O(N__19221),
            .I(N__19212));
    InMux I__4546 (
            .O(N__19220),
            .I(N__19209));
    Odrv4 I__4545 (
            .O(N__19215),
            .I(M_current_data_qZ0Z_3));
    LocalMux I__4544 (
            .O(N__19212),
            .I(M_current_data_qZ0Z_3));
    LocalMux I__4543 (
            .O(N__19209),
            .I(M_current_data_qZ0Z_3));
    ClkMux I__4542 (
            .O(N__19202),
            .I(N__18923));
    ClkMux I__4541 (
            .O(N__19201),
            .I(N__18923));
    ClkMux I__4540 (
            .O(N__19200),
            .I(N__18923));
    ClkMux I__4539 (
            .O(N__19199),
            .I(N__18923));
    ClkMux I__4538 (
            .O(N__19198),
            .I(N__18923));
    ClkMux I__4537 (
            .O(N__19197),
            .I(N__18923));
    ClkMux I__4536 (
            .O(N__19196),
            .I(N__18923));
    ClkMux I__4535 (
            .O(N__19195),
            .I(N__18923));
    ClkMux I__4534 (
            .O(N__19194),
            .I(N__18923));
    ClkMux I__4533 (
            .O(N__19193),
            .I(N__18923));
    ClkMux I__4532 (
            .O(N__19192),
            .I(N__18923));
    ClkMux I__4531 (
            .O(N__19191),
            .I(N__18923));
    ClkMux I__4530 (
            .O(N__19190),
            .I(N__18923));
    ClkMux I__4529 (
            .O(N__19189),
            .I(N__18923));
    ClkMux I__4528 (
            .O(N__19188),
            .I(N__18923));
    ClkMux I__4527 (
            .O(N__19187),
            .I(N__18923));
    ClkMux I__4526 (
            .O(N__19186),
            .I(N__18923));
    ClkMux I__4525 (
            .O(N__19185),
            .I(N__18923));
    ClkMux I__4524 (
            .O(N__19184),
            .I(N__18923));
    ClkMux I__4523 (
            .O(N__19183),
            .I(N__18923));
    ClkMux I__4522 (
            .O(N__19182),
            .I(N__18923));
    ClkMux I__4521 (
            .O(N__19181),
            .I(N__18923));
    ClkMux I__4520 (
            .O(N__19180),
            .I(N__18923));
    ClkMux I__4519 (
            .O(N__19179),
            .I(N__18923));
    ClkMux I__4518 (
            .O(N__19178),
            .I(N__18923));
    ClkMux I__4517 (
            .O(N__19177),
            .I(N__18923));
    ClkMux I__4516 (
            .O(N__19176),
            .I(N__18923));
    ClkMux I__4515 (
            .O(N__19175),
            .I(N__18923));
    ClkMux I__4514 (
            .O(N__19174),
            .I(N__18923));
    ClkMux I__4513 (
            .O(N__19173),
            .I(N__18923));
    ClkMux I__4512 (
            .O(N__19172),
            .I(N__18923));
    ClkMux I__4511 (
            .O(N__19171),
            .I(N__18923));
    ClkMux I__4510 (
            .O(N__19170),
            .I(N__18923));
    ClkMux I__4509 (
            .O(N__19169),
            .I(N__18923));
    ClkMux I__4508 (
            .O(N__19168),
            .I(N__18923));
    ClkMux I__4507 (
            .O(N__19167),
            .I(N__18923));
    ClkMux I__4506 (
            .O(N__19166),
            .I(N__18923));
    ClkMux I__4505 (
            .O(N__19165),
            .I(N__18923));
    ClkMux I__4504 (
            .O(N__19164),
            .I(N__18923));
    ClkMux I__4503 (
            .O(N__19163),
            .I(N__18923));
    ClkMux I__4502 (
            .O(N__19162),
            .I(N__18923));
    ClkMux I__4501 (
            .O(N__19161),
            .I(N__18923));
    ClkMux I__4500 (
            .O(N__19160),
            .I(N__18923));
    ClkMux I__4499 (
            .O(N__19159),
            .I(N__18923));
    ClkMux I__4498 (
            .O(N__19158),
            .I(N__18923));
    ClkMux I__4497 (
            .O(N__19157),
            .I(N__18923));
    ClkMux I__4496 (
            .O(N__19156),
            .I(N__18923));
    ClkMux I__4495 (
            .O(N__19155),
            .I(N__18923));
    ClkMux I__4494 (
            .O(N__19154),
            .I(N__18923));
    ClkMux I__4493 (
            .O(N__19153),
            .I(N__18923));
    ClkMux I__4492 (
            .O(N__19152),
            .I(N__18923));
    ClkMux I__4491 (
            .O(N__19151),
            .I(N__18923));
    ClkMux I__4490 (
            .O(N__19150),
            .I(N__18923));
    ClkMux I__4489 (
            .O(N__19149),
            .I(N__18923));
    ClkMux I__4488 (
            .O(N__19148),
            .I(N__18923));
    ClkMux I__4487 (
            .O(N__19147),
            .I(N__18923));
    ClkMux I__4486 (
            .O(N__19146),
            .I(N__18923));
    ClkMux I__4485 (
            .O(N__19145),
            .I(N__18923));
    ClkMux I__4484 (
            .O(N__19144),
            .I(N__18923));
    ClkMux I__4483 (
            .O(N__19143),
            .I(N__18923));
    ClkMux I__4482 (
            .O(N__19142),
            .I(N__18923));
    ClkMux I__4481 (
            .O(N__19141),
            .I(N__18923));
    ClkMux I__4480 (
            .O(N__19140),
            .I(N__18923));
    ClkMux I__4479 (
            .O(N__19139),
            .I(N__18923));
    ClkMux I__4478 (
            .O(N__19138),
            .I(N__18923));
    ClkMux I__4477 (
            .O(N__19137),
            .I(N__18923));
    ClkMux I__4476 (
            .O(N__19136),
            .I(N__18923));
    ClkMux I__4475 (
            .O(N__19135),
            .I(N__18923));
    ClkMux I__4474 (
            .O(N__19134),
            .I(N__18923));
    ClkMux I__4473 (
            .O(N__19133),
            .I(N__18923));
    ClkMux I__4472 (
            .O(N__19132),
            .I(N__18923));
    ClkMux I__4471 (
            .O(N__19131),
            .I(N__18923));
    ClkMux I__4470 (
            .O(N__19130),
            .I(N__18923));
    ClkMux I__4469 (
            .O(N__19129),
            .I(N__18923));
    ClkMux I__4468 (
            .O(N__19128),
            .I(N__18923));
    ClkMux I__4467 (
            .O(N__19127),
            .I(N__18923));
    ClkMux I__4466 (
            .O(N__19126),
            .I(N__18923));
    ClkMux I__4465 (
            .O(N__19125),
            .I(N__18923));
    ClkMux I__4464 (
            .O(N__19124),
            .I(N__18923));
    ClkMux I__4463 (
            .O(N__19123),
            .I(N__18923));
    ClkMux I__4462 (
            .O(N__19122),
            .I(N__18923));
    ClkMux I__4461 (
            .O(N__19121),
            .I(N__18923));
    ClkMux I__4460 (
            .O(N__19120),
            .I(N__18923));
    ClkMux I__4459 (
            .O(N__19119),
            .I(N__18923));
    ClkMux I__4458 (
            .O(N__19118),
            .I(N__18923));
    ClkMux I__4457 (
            .O(N__19117),
            .I(N__18923));
    ClkMux I__4456 (
            .O(N__19116),
            .I(N__18923));
    ClkMux I__4455 (
            .O(N__19115),
            .I(N__18923));
    ClkMux I__4454 (
            .O(N__19114),
            .I(N__18923));
    ClkMux I__4453 (
            .O(N__19113),
            .I(N__18923));
    ClkMux I__4452 (
            .O(N__19112),
            .I(N__18923));
    ClkMux I__4451 (
            .O(N__19111),
            .I(N__18923));
    ClkMux I__4450 (
            .O(N__19110),
            .I(N__18923));
    GlobalMux I__4449 (
            .O(N__18923),
            .I(N__18920));
    gio2CtrlBuf I__4448 (
            .O(N__18920),
            .I(clk_c_g));
    InMux I__4447 (
            .O(N__18917),
            .I(N__18914));
    LocalMux I__4446 (
            .O(N__18914),
            .I(N__18911));
    Span4Mux_v I__4445 (
            .O(N__18911),
            .I(N__18908));
    Odrv4 I__4444 (
            .O(N__18908),
            .I(port_address_c_4));
    InMux I__4443 (
            .O(N__18905),
            .I(N__18902));
    LocalMux I__4442 (
            .O(N__18902),
            .I(N__18899));
    Span4Mux_v I__4441 (
            .O(N__18899),
            .I(N__18896));
    Span4Mux_v I__4440 (
            .O(N__18896),
            .I(N__18893));
    Span4Mux_v I__4439 (
            .O(N__18893),
            .I(N__18890));
    Span4Mux_v I__4438 (
            .O(N__18890),
            .I(N__18887));
    Odrv4 I__4437 (
            .O(N__18887),
            .I(port_address_c_7));
    CascadeMux I__4436 (
            .O(N__18884),
            .I(N__18881));
    InMux I__4435 (
            .O(N__18881),
            .I(N__18878));
    LocalMux I__4434 (
            .O(N__18878),
            .I(N__18875));
    Span12Mux_v I__4433 (
            .O(N__18875),
            .I(N__18872));
    Odrv12 I__4432 (
            .O(N__18872),
            .I(port_address_c_3));
    InMux I__4431 (
            .O(N__18869),
            .I(N__18866));
    LocalMux I__4430 (
            .O(N__18866),
            .I(N__18863));
    Span12Mux_s10_h I__4429 (
            .O(N__18863),
            .I(N__18860));
    Span12Mux_h I__4428 (
            .O(N__18860),
            .I(N__18856));
    InMux I__4427 (
            .O(N__18859),
            .I(N__18853));
    Odrv12 I__4426 (
            .O(N__18856),
            .I(port_rw_c));
    LocalMux I__4425 (
            .O(N__18853),
            .I(port_rw_c));
    CascadeMux I__4424 (
            .O(N__18848),
            .I(N__18845));
    InMux I__4423 (
            .O(N__18845),
            .I(N__18842));
    LocalMux I__4422 (
            .O(N__18842),
            .I(N__18839));
    Span12Mux_v I__4421 (
            .O(N__18839),
            .I(N__18836));
    Span12Mux_h I__4420 (
            .O(N__18836),
            .I(N__18833));
    Odrv12 I__4419 (
            .O(N__18833),
            .I(\this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4Z0Z_0 ));
    CascadeMux I__4418 (
            .O(N__18830),
            .I(N__18827));
    CascadeBuf I__4417 (
            .O(N__18827),
            .I(N__18824));
    CascadeMux I__4416 (
            .O(N__18824),
            .I(N__18821));
    CascadeBuf I__4415 (
            .O(N__18821),
            .I(N__18818));
    CascadeMux I__4414 (
            .O(N__18818),
            .I(N__18815));
    CascadeBuf I__4413 (
            .O(N__18815),
            .I(N__18812));
    CascadeMux I__4412 (
            .O(N__18812),
            .I(N__18809));
    CascadeBuf I__4411 (
            .O(N__18809),
            .I(N__18806));
    CascadeMux I__4410 (
            .O(N__18806),
            .I(N__18803));
    CascadeBuf I__4409 (
            .O(N__18803),
            .I(N__18800));
    CascadeMux I__4408 (
            .O(N__18800),
            .I(N__18797));
    CascadeBuf I__4407 (
            .O(N__18797),
            .I(N__18794));
    CascadeMux I__4406 (
            .O(N__18794),
            .I(N__18791));
    CascadeBuf I__4405 (
            .O(N__18791),
            .I(N__18788));
    CascadeMux I__4404 (
            .O(N__18788),
            .I(N__18785));
    CascadeBuf I__4403 (
            .O(N__18785),
            .I(N__18782));
    CascadeMux I__4402 (
            .O(N__18782),
            .I(N__18779));
    CascadeBuf I__4401 (
            .O(N__18779),
            .I(N__18776));
    CascadeMux I__4400 (
            .O(N__18776),
            .I(N__18773));
    CascadeBuf I__4399 (
            .O(N__18773),
            .I(N__18770));
    CascadeMux I__4398 (
            .O(N__18770),
            .I(N__18767));
    CascadeBuf I__4397 (
            .O(N__18767),
            .I(N__18764));
    CascadeMux I__4396 (
            .O(N__18764),
            .I(N__18761));
    CascadeBuf I__4395 (
            .O(N__18761),
            .I(N__18758));
    CascadeMux I__4394 (
            .O(N__18758),
            .I(N__18755));
    CascadeBuf I__4393 (
            .O(N__18755),
            .I(N__18752));
    CascadeMux I__4392 (
            .O(N__18752),
            .I(N__18749));
    CascadeBuf I__4391 (
            .O(N__18749),
            .I(N__18746));
    CascadeMux I__4390 (
            .O(N__18746),
            .I(N__18743));
    CascadeBuf I__4389 (
            .O(N__18743),
            .I(N__18740));
    CascadeMux I__4388 (
            .O(N__18740),
            .I(N__18737));
    InMux I__4387 (
            .O(N__18737),
            .I(N__18734));
    LocalMux I__4386 (
            .O(N__18734),
            .I(N__18731));
    Span4Mux_s1_v I__4385 (
            .O(N__18731),
            .I(N__18728));
    Span4Mux_v I__4384 (
            .O(N__18728),
            .I(N__18725));
    Odrv4 I__4383 (
            .O(N__18725),
            .I(M_current_address_qZ0Z_2));
    CascadeMux I__4382 (
            .O(N__18722),
            .I(N__18719));
    CascadeBuf I__4381 (
            .O(N__18719),
            .I(N__18716));
    CascadeMux I__4380 (
            .O(N__18716),
            .I(N__18713));
    CascadeBuf I__4379 (
            .O(N__18713),
            .I(N__18710));
    CascadeMux I__4378 (
            .O(N__18710),
            .I(N__18707));
    CascadeBuf I__4377 (
            .O(N__18707),
            .I(N__18704));
    CascadeMux I__4376 (
            .O(N__18704),
            .I(N__18701));
    CascadeBuf I__4375 (
            .O(N__18701),
            .I(N__18698));
    CascadeMux I__4374 (
            .O(N__18698),
            .I(N__18695));
    CascadeBuf I__4373 (
            .O(N__18695),
            .I(N__18692));
    CascadeMux I__4372 (
            .O(N__18692),
            .I(N__18689));
    CascadeBuf I__4371 (
            .O(N__18689),
            .I(N__18686));
    CascadeMux I__4370 (
            .O(N__18686),
            .I(N__18683));
    CascadeBuf I__4369 (
            .O(N__18683),
            .I(N__18680));
    CascadeMux I__4368 (
            .O(N__18680),
            .I(N__18677));
    CascadeBuf I__4367 (
            .O(N__18677),
            .I(N__18674));
    CascadeMux I__4366 (
            .O(N__18674),
            .I(N__18671));
    CascadeBuf I__4365 (
            .O(N__18671),
            .I(N__18668));
    CascadeMux I__4364 (
            .O(N__18668),
            .I(N__18665));
    CascadeBuf I__4363 (
            .O(N__18665),
            .I(N__18662));
    CascadeMux I__4362 (
            .O(N__18662),
            .I(N__18659));
    CascadeBuf I__4361 (
            .O(N__18659),
            .I(N__18656));
    CascadeMux I__4360 (
            .O(N__18656),
            .I(N__18653));
    CascadeBuf I__4359 (
            .O(N__18653),
            .I(N__18650));
    CascadeMux I__4358 (
            .O(N__18650),
            .I(N__18647));
    CascadeBuf I__4357 (
            .O(N__18647),
            .I(N__18644));
    CascadeMux I__4356 (
            .O(N__18644),
            .I(N__18641));
    CascadeBuf I__4355 (
            .O(N__18641),
            .I(N__18638));
    CascadeMux I__4354 (
            .O(N__18638),
            .I(N__18635));
    CascadeBuf I__4353 (
            .O(N__18635),
            .I(N__18632));
    CascadeMux I__4352 (
            .O(N__18632),
            .I(N__18629));
    InMux I__4351 (
            .O(N__18629),
            .I(N__18626));
    LocalMux I__4350 (
            .O(N__18626),
            .I(N__18623));
    Span4Mux_s1_v I__4349 (
            .O(N__18623),
            .I(N__18620));
    Span4Mux_v I__4348 (
            .O(N__18620),
            .I(N__18617));
    Odrv4 I__4347 (
            .O(N__18617),
            .I(M_current_address_qZ0Z_9));
    InMux I__4346 (
            .O(N__18614),
            .I(N__18611));
    LocalMux I__4345 (
            .O(N__18611),
            .I(N__18607));
    InMux I__4344 (
            .O(N__18610),
            .I(N__18604));
    Span4Mux_v I__4343 (
            .O(N__18607),
            .I(N__18598));
    LocalMux I__4342 (
            .O(N__18604),
            .I(N__18598));
    InMux I__4341 (
            .O(N__18603),
            .I(N__18595));
    Span4Mux_v I__4340 (
            .O(N__18598),
            .I(N__18589));
    LocalMux I__4339 (
            .O(N__18595),
            .I(N__18589));
    InMux I__4338 (
            .O(N__18594),
            .I(N__18586));
    Span4Mux_v I__4337 (
            .O(N__18589),
            .I(N__18580));
    LocalMux I__4336 (
            .O(N__18586),
            .I(N__18580));
    InMux I__4335 (
            .O(N__18585),
            .I(N__18577));
    Span4Mux_v I__4334 (
            .O(N__18580),
            .I(N__18570));
    LocalMux I__4333 (
            .O(N__18577),
            .I(N__18570));
    InMux I__4332 (
            .O(N__18576),
            .I(N__18567));
    InMux I__4331 (
            .O(N__18575),
            .I(N__18564));
    Span4Mux_v I__4330 (
            .O(N__18570),
            .I(N__18559));
    LocalMux I__4329 (
            .O(N__18567),
            .I(N__18559));
    LocalMux I__4328 (
            .O(N__18564),
            .I(N__18556));
    Span4Mux_v I__4327 (
            .O(N__18559),
            .I(N__18549));
    Span4Mux_s3_v I__4326 (
            .O(N__18556),
            .I(N__18549));
    InMux I__4325 (
            .O(N__18555),
            .I(N__18546));
    InMux I__4324 (
            .O(N__18554),
            .I(N__18543));
    Odrv4 I__4323 (
            .O(N__18549),
            .I(M_current_data_qZ0Z_0));
    LocalMux I__4322 (
            .O(N__18546),
            .I(M_current_data_qZ0Z_0));
    LocalMux I__4321 (
            .O(N__18543),
            .I(M_current_data_qZ0Z_0));
    CascadeMux I__4320 (
            .O(N__18536),
            .I(N__18533));
    CascadeBuf I__4319 (
            .O(N__18533),
            .I(N__18530));
    CascadeMux I__4318 (
            .O(N__18530),
            .I(N__18527));
    CascadeBuf I__4317 (
            .O(N__18527),
            .I(N__18524));
    CascadeMux I__4316 (
            .O(N__18524),
            .I(N__18521));
    CascadeBuf I__4315 (
            .O(N__18521),
            .I(N__18518));
    CascadeMux I__4314 (
            .O(N__18518),
            .I(N__18515));
    CascadeBuf I__4313 (
            .O(N__18515),
            .I(N__18512));
    CascadeMux I__4312 (
            .O(N__18512),
            .I(N__18509));
    CascadeBuf I__4311 (
            .O(N__18509),
            .I(N__18506));
    CascadeMux I__4310 (
            .O(N__18506),
            .I(N__18503));
    CascadeBuf I__4309 (
            .O(N__18503),
            .I(N__18500));
    CascadeMux I__4308 (
            .O(N__18500),
            .I(N__18497));
    CascadeBuf I__4307 (
            .O(N__18497),
            .I(N__18494));
    CascadeMux I__4306 (
            .O(N__18494),
            .I(N__18491));
    CascadeBuf I__4305 (
            .O(N__18491),
            .I(N__18488));
    CascadeMux I__4304 (
            .O(N__18488),
            .I(N__18485));
    CascadeBuf I__4303 (
            .O(N__18485),
            .I(N__18482));
    CascadeMux I__4302 (
            .O(N__18482),
            .I(N__18479));
    CascadeBuf I__4301 (
            .O(N__18479),
            .I(N__18476));
    CascadeMux I__4300 (
            .O(N__18476),
            .I(N__18473));
    CascadeBuf I__4299 (
            .O(N__18473),
            .I(N__18470));
    CascadeMux I__4298 (
            .O(N__18470),
            .I(N__18467));
    CascadeBuf I__4297 (
            .O(N__18467),
            .I(N__18464));
    CascadeMux I__4296 (
            .O(N__18464),
            .I(N__18461));
    CascadeBuf I__4295 (
            .O(N__18461),
            .I(N__18458));
    CascadeMux I__4294 (
            .O(N__18458),
            .I(N__18455));
    CascadeBuf I__4293 (
            .O(N__18455),
            .I(N__18452));
    CascadeMux I__4292 (
            .O(N__18452),
            .I(N__18449));
    CascadeBuf I__4291 (
            .O(N__18449),
            .I(N__18446));
    CascadeMux I__4290 (
            .O(N__18446),
            .I(N__18443));
    InMux I__4289 (
            .O(N__18443),
            .I(N__18440));
    LocalMux I__4288 (
            .O(N__18440),
            .I(N__18437));
    Span4Mux_s2_v I__4287 (
            .O(N__18437),
            .I(N__18434));
    Odrv4 I__4286 (
            .O(N__18434),
            .I(M_current_address_qZ0Z_1));
    CascadeMux I__4285 (
            .O(N__18431),
            .I(N__18428));
    CascadeBuf I__4284 (
            .O(N__18428),
            .I(N__18425));
    CascadeMux I__4283 (
            .O(N__18425),
            .I(N__18422));
    CascadeBuf I__4282 (
            .O(N__18422),
            .I(N__18419));
    CascadeMux I__4281 (
            .O(N__18419),
            .I(N__18416));
    CascadeBuf I__4280 (
            .O(N__18416),
            .I(N__18413));
    CascadeMux I__4279 (
            .O(N__18413),
            .I(N__18410));
    CascadeBuf I__4278 (
            .O(N__18410),
            .I(N__18407));
    CascadeMux I__4277 (
            .O(N__18407),
            .I(N__18404));
    CascadeBuf I__4276 (
            .O(N__18404),
            .I(N__18401));
    CascadeMux I__4275 (
            .O(N__18401),
            .I(N__18398));
    CascadeBuf I__4274 (
            .O(N__18398),
            .I(N__18395));
    CascadeMux I__4273 (
            .O(N__18395),
            .I(N__18392));
    CascadeBuf I__4272 (
            .O(N__18392),
            .I(N__18389));
    CascadeMux I__4271 (
            .O(N__18389),
            .I(N__18386));
    CascadeBuf I__4270 (
            .O(N__18386),
            .I(N__18383));
    CascadeMux I__4269 (
            .O(N__18383),
            .I(N__18380));
    CascadeBuf I__4268 (
            .O(N__18380),
            .I(N__18377));
    CascadeMux I__4267 (
            .O(N__18377),
            .I(N__18374));
    CascadeBuf I__4266 (
            .O(N__18374),
            .I(N__18371));
    CascadeMux I__4265 (
            .O(N__18371),
            .I(N__18368));
    CascadeBuf I__4264 (
            .O(N__18368),
            .I(N__18365));
    CascadeMux I__4263 (
            .O(N__18365),
            .I(N__18362));
    CascadeBuf I__4262 (
            .O(N__18362),
            .I(N__18359));
    CascadeMux I__4261 (
            .O(N__18359),
            .I(N__18356));
    CascadeBuf I__4260 (
            .O(N__18356),
            .I(N__18353));
    CascadeMux I__4259 (
            .O(N__18353),
            .I(N__18350));
    CascadeBuf I__4258 (
            .O(N__18350),
            .I(N__18347));
    CascadeMux I__4257 (
            .O(N__18347),
            .I(N__18344));
    CascadeBuf I__4256 (
            .O(N__18344),
            .I(N__18341));
    CascadeMux I__4255 (
            .O(N__18341),
            .I(N__18338));
    InMux I__4254 (
            .O(N__18338),
            .I(N__18335));
    LocalMux I__4253 (
            .O(N__18335),
            .I(N__18332));
    Span4Mux_s3_v I__4252 (
            .O(N__18332),
            .I(N__18329));
    Odrv4 I__4251 (
            .O(N__18329),
            .I(M_current_address_qZ0Z_3));
    CEMux I__4250 (
            .O(N__18326),
            .I(N__18322));
    CEMux I__4249 (
            .O(N__18325),
            .I(N__18319));
    LocalMux I__4248 (
            .O(N__18322),
            .I(N__18311));
    LocalMux I__4247 (
            .O(N__18319),
            .I(N__18311));
    CEMux I__4246 (
            .O(N__18318),
            .I(N__18308));
    CEMux I__4245 (
            .O(N__18317),
            .I(N__18305));
    CEMux I__4244 (
            .O(N__18316),
            .I(N__18302));
    Span4Mux_v I__4243 (
            .O(N__18311),
            .I(N__18296));
    LocalMux I__4242 (
            .O(N__18308),
            .I(N__18296));
    LocalMux I__4241 (
            .O(N__18305),
            .I(N__18291));
    LocalMux I__4240 (
            .O(N__18302),
            .I(N__18291));
    CEMux I__4239 (
            .O(N__18301),
            .I(N__18288));
    Span4Mux_v I__4238 (
            .O(N__18296),
            .I(N__18281));
    Span4Mux_v I__4237 (
            .O(N__18291),
            .I(N__18281));
    LocalMux I__4236 (
            .O(N__18288),
            .I(N__18281));
    Odrv4 I__4235 (
            .O(N__18281),
            .I(M_current_address_q_0_0));
    CascadeMux I__4234 (
            .O(N__18278),
            .I(N__18275));
    CascadeBuf I__4233 (
            .O(N__18275),
            .I(N__18272));
    CascadeMux I__4232 (
            .O(N__18272),
            .I(N__18269));
    CascadeBuf I__4231 (
            .O(N__18269),
            .I(N__18266));
    CascadeMux I__4230 (
            .O(N__18266),
            .I(N__18263));
    CascadeBuf I__4229 (
            .O(N__18263),
            .I(N__18260));
    CascadeMux I__4228 (
            .O(N__18260),
            .I(N__18257));
    CascadeBuf I__4227 (
            .O(N__18257),
            .I(N__18254));
    CascadeMux I__4226 (
            .O(N__18254),
            .I(N__18251));
    CascadeBuf I__4225 (
            .O(N__18251),
            .I(N__18248));
    CascadeMux I__4224 (
            .O(N__18248),
            .I(N__18245));
    CascadeBuf I__4223 (
            .O(N__18245),
            .I(N__18242));
    CascadeMux I__4222 (
            .O(N__18242),
            .I(N__18239));
    CascadeBuf I__4221 (
            .O(N__18239),
            .I(N__18236));
    CascadeMux I__4220 (
            .O(N__18236),
            .I(N__18233));
    CascadeBuf I__4219 (
            .O(N__18233),
            .I(N__18230));
    CascadeMux I__4218 (
            .O(N__18230),
            .I(N__18227));
    CascadeBuf I__4217 (
            .O(N__18227),
            .I(N__18224));
    CascadeMux I__4216 (
            .O(N__18224),
            .I(N__18221));
    CascadeBuf I__4215 (
            .O(N__18221),
            .I(N__18218));
    CascadeMux I__4214 (
            .O(N__18218),
            .I(N__18215));
    CascadeBuf I__4213 (
            .O(N__18215),
            .I(N__18212));
    CascadeMux I__4212 (
            .O(N__18212),
            .I(N__18209));
    CascadeBuf I__4211 (
            .O(N__18209),
            .I(N__18206));
    CascadeMux I__4210 (
            .O(N__18206),
            .I(N__18203));
    CascadeBuf I__4209 (
            .O(N__18203),
            .I(N__18200));
    CascadeMux I__4208 (
            .O(N__18200),
            .I(N__18197));
    CascadeBuf I__4207 (
            .O(N__18197),
            .I(N__18194));
    CascadeMux I__4206 (
            .O(N__18194),
            .I(N__18191));
    CascadeBuf I__4205 (
            .O(N__18191),
            .I(N__18188));
    CascadeMux I__4204 (
            .O(N__18188),
            .I(N__18185));
    InMux I__4203 (
            .O(N__18185),
            .I(N__18182));
    LocalMux I__4202 (
            .O(N__18182),
            .I(N__18179));
    Span4Mux_s1_v I__4201 (
            .O(N__18179),
            .I(N__18176));
    Odrv4 I__4200 (
            .O(N__18176),
            .I(M_current_address_qZ0Z_10));
    CascadeMux I__4199 (
            .O(N__18173),
            .I(N__18170));
    InMux I__4198 (
            .O(N__18170),
            .I(N__18166));
    InMux I__4197 (
            .O(N__18169),
            .I(N__18163));
    LocalMux I__4196 (
            .O(N__18166),
            .I(N__18160));
    LocalMux I__4195 (
            .O(N__18163),
            .I(N__18157));
    Span4Mux_v I__4194 (
            .O(N__18160),
            .I(N__18151));
    Span4Mux_v I__4193 (
            .O(N__18157),
            .I(N__18151));
    InMux I__4192 (
            .O(N__18156),
            .I(N__18148));
    Sp12to4 I__4191 (
            .O(N__18151),
            .I(N__18143));
    LocalMux I__4190 (
            .O(N__18148),
            .I(N__18143));
    Span12Mux_h I__4189 (
            .O(N__18143),
            .I(N__18140));
    Odrv12 I__4188 (
            .O(N__18140),
            .I(port_data_c_0));
    CascadeMux I__4187 (
            .O(N__18137),
            .I(N__18134));
    CascadeBuf I__4186 (
            .O(N__18134),
            .I(N__18131));
    CascadeMux I__4185 (
            .O(N__18131),
            .I(N__18128));
    CascadeBuf I__4184 (
            .O(N__18128),
            .I(N__18125));
    CascadeMux I__4183 (
            .O(N__18125),
            .I(N__18122));
    CascadeBuf I__4182 (
            .O(N__18122),
            .I(N__18119));
    CascadeMux I__4181 (
            .O(N__18119),
            .I(N__18116));
    CascadeBuf I__4180 (
            .O(N__18116),
            .I(N__18113));
    CascadeMux I__4179 (
            .O(N__18113),
            .I(N__18110));
    CascadeBuf I__4178 (
            .O(N__18110),
            .I(N__18107));
    CascadeMux I__4177 (
            .O(N__18107),
            .I(N__18104));
    CascadeBuf I__4176 (
            .O(N__18104),
            .I(N__18101));
    CascadeMux I__4175 (
            .O(N__18101),
            .I(N__18098));
    CascadeBuf I__4174 (
            .O(N__18098),
            .I(N__18095));
    CascadeMux I__4173 (
            .O(N__18095),
            .I(N__18092));
    CascadeBuf I__4172 (
            .O(N__18092),
            .I(N__18089));
    CascadeMux I__4171 (
            .O(N__18089),
            .I(N__18086));
    CascadeBuf I__4170 (
            .O(N__18086),
            .I(N__18083));
    CascadeMux I__4169 (
            .O(N__18083),
            .I(N__18080));
    CascadeBuf I__4168 (
            .O(N__18080),
            .I(N__18077));
    CascadeMux I__4167 (
            .O(N__18077),
            .I(N__18074));
    CascadeBuf I__4166 (
            .O(N__18074),
            .I(N__18071));
    CascadeMux I__4165 (
            .O(N__18071),
            .I(N__18068));
    CascadeBuf I__4164 (
            .O(N__18068),
            .I(N__18065));
    CascadeMux I__4163 (
            .O(N__18065),
            .I(N__18062));
    CascadeBuf I__4162 (
            .O(N__18062),
            .I(N__18059));
    CascadeMux I__4161 (
            .O(N__18059),
            .I(N__18056));
    CascadeBuf I__4160 (
            .O(N__18056),
            .I(N__18053));
    CascadeMux I__4159 (
            .O(N__18053),
            .I(N__18050));
    CascadeBuf I__4158 (
            .O(N__18050),
            .I(N__18047));
    CascadeMux I__4157 (
            .O(N__18047),
            .I(N__18044));
    InMux I__4156 (
            .O(N__18044),
            .I(N__18041));
    LocalMux I__4155 (
            .O(N__18041),
            .I(N__18038));
    Span4Mux_s1_v I__4154 (
            .O(N__18038),
            .I(N__18035));
    Odrv4 I__4153 (
            .O(N__18035),
            .I(M_current_address_qZ0Z_7));
    CascadeMux I__4152 (
            .O(N__18032),
            .I(N__18028));
    InMux I__4151 (
            .O(N__18031),
            .I(N__18025));
    InMux I__4150 (
            .O(N__18028),
            .I(N__18022));
    LocalMux I__4149 (
            .O(N__18025),
            .I(N__18018));
    LocalMux I__4148 (
            .O(N__18022),
            .I(N__18015));
    InMux I__4147 (
            .O(N__18021),
            .I(N__18012));
    Span4Mux_v I__4146 (
            .O(N__18018),
            .I(N__18009));
    Span4Mux_v I__4145 (
            .O(N__18015),
            .I(N__18006));
    LocalMux I__4144 (
            .O(N__18012),
            .I(N__18003));
    Sp12to4 I__4143 (
            .O(N__18009),
            .I(N__17998));
    Sp12to4 I__4142 (
            .O(N__18006),
            .I(N__17998));
    Span12Mux_h I__4141 (
            .O(N__18003),
            .I(N__17995));
    Span12Mux_h I__4140 (
            .O(N__17998),
            .I(N__17992));
    Odrv12 I__4139 (
            .O(N__17995),
            .I(port_data_c_1));
    Odrv12 I__4138 (
            .O(N__17992),
            .I(port_data_c_1));
    CascadeMux I__4137 (
            .O(N__17987),
            .I(N__17984));
    CascadeBuf I__4136 (
            .O(N__17984),
            .I(N__17981));
    CascadeMux I__4135 (
            .O(N__17981),
            .I(N__17978));
    CascadeBuf I__4134 (
            .O(N__17978),
            .I(N__17975));
    CascadeMux I__4133 (
            .O(N__17975),
            .I(N__17972));
    CascadeBuf I__4132 (
            .O(N__17972),
            .I(N__17969));
    CascadeMux I__4131 (
            .O(N__17969),
            .I(N__17966));
    CascadeBuf I__4130 (
            .O(N__17966),
            .I(N__17963));
    CascadeMux I__4129 (
            .O(N__17963),
            .I(N__17960));
    CascadeBuf I__4128 (
            .O(N__17960),
            .I(N__17957));
    CascadeMux I__4127 (
            .O(N__17957),
            .I(N__17954));
    CascadeBuf I__4126 (
            .O(N__17954),
            .I(N__17951));
    CascadeMux I__4125 (
            .O(N__17951),
            .I(N__17948));
    CascadeBuf I__4124 (
            .O(N__17948),
            .I(N__17945));
    CascadeMux I__4123 (
            .O(N__17945),
            .I(N__17942));
    CascadeBuf I__4122 (
            .O(N__17942),
            .I(N__17939));
    CascadeMux I__4121 (
            .O(N__17939),
            .I(N__17936));
    CascadeBuf I__4120 (
            .O(N__17936),
            .I(N__17933));
    CascadeMux I__4119 (
            .O(N__17933),
            .I(N__17930));
    CascadeBuf I__4118 (
            .O(N__17930),
            .I(N__17927));
    CascadeMux I__4117 (
            .O(N__17927),
            .I(N__17924));
    CascadeBuf I__4116 (
            .O(N__17924),
            .I(N__17921));
    CascadeMux I__4115 (
            .O(N__17921),
            .I(N__17918));
    CascadeBuf I__4114 (
            .O(N__17918),
            .I(N__17915));
    CascadeMux I__4113 (
            .O(N__17915),
            .I(N__17912));
    CascadeBuf I__4112 (
            .O(N__17912),
            .I(N__17909));
    CascadeMux I__4111 (
            .O(N__17909),
            .I(N__17906));
    CascadeBuf I__4110 (
            .O(N__17906),
            .I(N__17903));
    CascadeMux I__4109 (
            .O(N__17903),
            .I(N__17900));
    CascadeBuf I__4108 (
            .O(N__17900),
            .I(N__17897));
    CascadeMux I__4107 (
            .O(N__17897),
            .I(N__17894));
    InMux I__4106 (
            .O(N__17894),
            .I(N__17891));
    LocalMux I__4105 (
            .O(N__17891),
            .I(N__17888));
    Odrv4 I__4104 (
            .O(N__17888),
            .I(M_current_address_qZ0Z_8));
    CEMux I__4103 (
            .O(N__17885),
            .I(N__17882));
    LocalMux I__4102 (
            .O(N__17882),
            .I(N__17876));
    CEMux I__4101 (
            .O(N__17881),
            .I(N__17873));
    CEMux I__4100 (
            .O(N__17880),
            .I(N__17870));
    CEMux I__4099 (
            .O(N__17879),
            .I(N__17865));
    Span4Mux_v I__4098 (
            .O(N__17876),
            .I(N__17860));
    LocalMux I__4097 (
            .O(N__17873),
            .I(N__17860));
    LocalMux I__4096 (
            .O(N__17870),
            .I(N__17857));
    CEMux I__4095 (
            .O(N__17869),
            .I(N__17854));
    CEMux I__4094 (
            .O(N__17868),
            .I(N__17851));
    LocalMux I__4093 (
            .O(N__17865),
            .I(N__17846));
    Sp12to4 I__4092 (
            .O(N__17860),
            .I(N__17846));
    Span4Mux_h I__4091 (
            .O(N__17857),
            .I(N__17843));
    LocalMux I__4090 (
            .O(N__17854),
            .I(N__17840));
    LocalMux I__4089 (
            .O(N__17851),
            .I(N__17837));
    Span12Mux_v I__4088 (
            .O(N__17846),
            .I(N__17834));
    Span4Mux_v I__4087 (
            .O(N__17843),
            .I(N__17831));
    Span4Mux_h I__4086 (
            .O(N__17840),
            .I(N__17828));
    Span4Mux_h I__4085 (
            .O(N__17837),
            .I(N__17825));
    Odrv12 I__4084 (
            .O(N__17834),
            .I(M_current_address_q_0_6_0));
    Odrv4 I__4083 (
            .O(N__17831),
            .I(M_current_address_q_0_6_0));
    Odrv4 I__4082 (
            .O(N__17828),
            .I(M_current_address_q_0_6_0));
    Odrv4 I__4081 (
            .O(N__17825),
            .I(M_current_address_q_0_6_0));
    InMux I__4080 (
            .O(N__17816),
            .I(N__17812));
    InMux I__4079 (
            .O(N__17815),
            .I(N__17809));
    LocalMux I__4078 (
            .O(N__17812),
            .I(N__17788));
    LocalMux I__4077 (
            .O(N__17809),
            .I(N__17785));
    SRMux I__4076 (
            .O(N__17808),
            .I(N__17744));
    SRMux I__4075 (
            .O(N__17807),
            .I(N__17744));
    SRMux I__4074 (
            .O(N__17806),
            .I(N__17744));
    SRMux I__4073 (
            .O(N__17805),
            .I(N__17744));
    SRMux I__4072 (
            .O(N__17804),
            .I(N__17744));
    SRMux I__4071 (
            .O(N__17803),
            .I(N__17744));
    SRMux I__4070 (
            .O(N__17802),
            .I(N__17744));
    SRMux I__4069 (
            .O(N__17801),
            .I(N__17744));
    SRMux I__4068 (
            .O(N__17800),
            .I(N__17744));
    SRMux I__4067 (
            .O(N__17799),
            .I(N__17744));
    SRMux I__4066 (
            .O(N__17798),
            .I(N__17744));
    SRMux I__4065 (
            .O(N__17797),
            .I(N__17744));
    SRMux I__4064 (
            .O(N__17796),
            .I(N__17744));
    SRMux I__4063 (
            .O(N__17795),
            .I(N__17744));
    SRMux I__4062 (
            .O(N__17794),
            .I(N__17744));
    SRMux I__4061 (
            .O(N__17793),
            .I(N__17744));
    SRMux I__4060 (
            .O(N__17792),
            .I(N__17744));
    SRMux I__4059 (
            .O(N__17791),
            .I(N__17744));
    Glb2LocalMux I__4058 (
            .O(N__17788),
            .I(N__17744));
    Glb2LocalMux I__4057 (
            .O(N__17785),
            .I(N__17744));
    GlobalMux I__4056 (
            .O(N__17744),
            .I(N__17741));
    gio2CtrlBuf I__4055 (
            .O(N__17741),
            .I(N_631_g));
    InMux I__4054 (
            .O(N__17738),
            .I(N__17735));
    LocalMux I__4053 (
            .O(N__17735),
            .I(N__17732));
    Span4Mux_h I__4052 (
            .O(N__17732),
            .I(N__17729));
    Sp12to4 I__4051 (
            .O(N__17729),
            .I(N__17726));
    Span12Mux_s10_v I__4050 (
            .O(N__17726),
            .I(N__17721));
    InMux I__4049 (
            .O(N__17725),
            .I(N__17715));
    InMux I__4048 (
            .O(N__17724),
            .I(N__17715));
    Span12Mux_v I__4047 (
            .O(N__17721),
            .I(N__17712));
    InMux I__4046 (
            .O(N__17720),
            .I(N__17709));
    LocalMux I__4045 (
            .O(N__17715),
            .I(N__17706));
    Odrv12 I__4044 (
            .O(N__17712),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_2 ));
    LocalMux I__4043 (
            .O(N__17709),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_2 ));
    Odrv4 I__4042 (
            .O(N__17706),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_2 ));
    InMux I__4041 (
            .O(N__17699),
            .I(N__17696));
    LocalMux I__4040 (
            .O(N__17696),
            .I(N__17693));
    Span4Mux_v I__4039 (
            .O(N__17693),
            .I(N__17690));
    Sp12to4 I__4038 (
            .O(N__17690),
            .I(N__17687));
    Span12Mux_h I__4037 (
            .O(N__17687),
            .I(N__17684));
    Span12Mux_v I__4036 (
            .O(N__17684),
            .I(N__17680));
    InMux I__4035 (
            .O(N__17683),
            .I(N__17677));
    Odrv12 I__4034 (
            .O(N__17680),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__4033 (
            .O(N__17677),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    InMux I__4032 (
            .O(N__17672),
            .I(N__17669));
    LocalMux I__4031 (
            .O(N__17669),
            .I(N__17666));
    Span4Mux_h I__4030 (
            .O(N__17666),
            .I(N__17663));
    Span4Mux_h I__4029 (
            .O(N__17663),
            .I(N__17659));
    InMux I__4028 (
            .O(N__17662),
            .I(N__17655));
    Sp12to4 I__4027 (
            .O(N__17659),
            .I(N__17651));
    InMux I__4026 (
            .O(N__17658),
            .I(N__17648));
    LocalMux I__4025 (
            .O(N__17655),
            .I(N__17645));
    InMux I__4024 (
            .O(N__17654),
            .I(N__17640));
    Span12Mux_v I__4023 (
            .O(N__17651),
            .I(N__17633));
    LocalMux I__4022 (
            .O(N__17648),
            .I(N__17630));
    Span4Mux_h I__4021 (
            .O(N__17645),
            .I(N__17627));
    InMux I__4020 (
            .O(N__17644),
            .I(N__17622));
    InMux I__4019 (
            .O(N__17643),
            .I(N__17622));
    LocalMux I__4018 (
            .O(N__17640),
            .I(N__17619));
    InMux I__4017 (
            .O(N__17639),
            .I(N__17614));
    InMux I__4016 (
            .O(N__17638),
            .I(N__17614));
    InMux I__4015 (
            .O(N__17637),
            .I(N__17611));
    InMux I__4014 (
            .O(N__17636),
            .I(N__17608));
    Odrv12 I__4013 (
            .O(N__17633),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    Odrv4 I__4012 (
            .O(N__17630),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    Odrv4 I__4011 (
            .O(N__17627),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    LocalMux I__4010 (
            .O(N__17622),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    Odrv4 I__4009 (
            .O(N__17619),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    LocalMux I__4008 (
            .O(N__17614),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    LocalMux I__4007 (
            .O(N__17611),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    LocalMux I__4006 (
            .O(N__17608),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    CascadeMux I__4005 (
            .O(N__17591),
            .I(N__17588));
    CascadeBuf I__4004 (
            .O(N__17588),
            .I(N__17585));
    CascadeMux I__4003 (
            .O(N__17585),
            .I(N__17582));
    CascadeBuf I__4002 (
            .O(N__17582),
            .I(N__17579));
    CascadeMux I__4001 (
            .O(N__17579),
            .I(N__17576));
    CascadeBuf I__4000 (
            .O(N__17576),
            .I(N__17573));
    CascadeMux I__3999 (
            .O(N__17573),
            .I(N__17570));
    CascadeBuf I__3998 (
            .O(N__17570),
            .I(N__17567));
    CascadeMux I__3997 (
            .O(N__17567),
            .I(N__17564));
    CascadeBuf I__3996 (
            .O(N__17564),
            .I(N__17561));
    CascadeMux I__3995 (
            .O(N__17561),
            .I(N__17558));
    CascadeBuf I__3994 (
            .O(N__17558),
            .I(N__17555));
    CascadeMux I__3993 (
            .O(N__17555),
            .I(N__17552));
    CascadeBuf I__3992 (
            .O(N__17552),
            .I(N__17549));
    CascadeMux I__3991 (
            .O(N__17549),
            .I(N__17546));
    CascadeBuf I__3990 (
            .O(N__17546),
            .I(N__17543));
    CascadeMux I__3989 (
            .O(N__17543),
            .I(N__17540));
    CascadeBuf I__3988 (
            .O(N__17540),
            .I(N__17537));
    CascadeMux I__3987 (
            .O(N__17537),
            .I(N__17534));
    CascadeBuf I__3986 (
            .O(N__17534),
            .I(N__17531));
    CascadeMux I__3985 (
            .O(N__17531),
            .I(N__17528));
    CascadeBuf I__3984 (
            .O(N__17528),
            .I(N__17525));
    CascadeMux I__3983 (
            .O(N__17525),
            .I(N__17522));
    CascadeBuf I__3982 (
            .O(N__17522),
            .I(N__17519));
    CascadeMux I__3981 (
            .O(N__17519),
            .I(N__17516));
    CascadeBuf I__3980 (
            .O(N__17516),
            .I(N__17513));
    CascadeMux I__3979 (
            .O(N__17513),
            .I(N__17510));
    CascadeBuf I__3978 (
            .O(N__17510),
            .I(N__17507));
    CascadeMux I__3977 (
            .O(N__17507),
            .I(N__17504));
    CascadeBuf I__3976 (
            .O(N__17504),
            .I(N__17501));
    CascadeMux I__3975 (
            .O(N__17501),
            .I(N__17498));
    InMux I__3974 (
            .O(N__17498),
            .I(N__17495));
    LocalMux I__3973 (
            .O(N__17495),
            .I(this_vga_signals_un14_address_if_generate_plus_mult1_un61_sum_i_3));
    InMux I__3972 (
            .O(N__17492),
            .I(N__17488));
    InMux I__3971 (
            .O(N__17491),
            .I(N__17485));
    LocalMux I__3970 (
            .O(N__17488),
            .I(N__17480));
    LocalMux I__3969 (
            .O(N__17485),
            .I(N__17480));
    Span12Mux_v I__3968 (
            .O(N__17480),
            .I(N__17477));
    Odrv12 I__3967 (
            .O(N__17477),
            .I(port_data_c_6));
    CascadeMux I__3966 (
            .O(N__17474),
            .I(N__17471));
    CascadeBuf I__3965 (
            .O(N__17471),
            .I(N__17468));
    CascadeMux I__3964 (
            .O(N__17468),
            .I(N__17465));
    CascadeBuf I__3963 (
            .O(N__17465),
            .I(N__17462));
    CascadeMux I__3962 (
            .O(N__17462),
            .I(N__17459));
    CascadeBuf I__3961 (
            .O(N__17459),
            .I(N__17456));
    CascadeMux I__3960 (
            .O(N__17456),
            .I(N__17453));
    CascadeBuf I__3959 (
            .O(N__17453),
            .I(N__17450));
    CascadeMux I__3958 (
            .O(N__17450),
            .I(N__17447));
    CascadeBuf I__3957 (
            .O(N__17447),
            .I(N__17444));
    CascadeMux I__3956 (
            .O(N__17444),
            .I(N__17441));
    CascadeBuf I__3955 (
            .O(N__17441),
            .I(N__17438));
    CascadeMux I__3954 (
            .O(N__17438),
            .I(N__17435));
    CascadeBuf I__3953 (
            .O(N__17435),
            .I(N__17432));
    CascadeMux I__3952 (
            .O(N__17432),
            .I(N__17429));
    CascadeBuf I__3951 (
            .O(N__17429),
            .I(N__17426));
    CascadeMux I__3950 (
            .O(N__17426),
            .I(N__17423));
    CascadeBuf I__3949 (
            .O(N__17423),
            .I(N__17420));
    CascadeMux I__3948 (
            .O(N__17420),
            .I(N__17417));
    CascadeBuf I__3947 (
            .O(N__17417),
            .I(N__17414));
    CascadeMux I__3946 (
            .O(N__17414),
            .I(N__17411));
    CascadeBuf I__3945 (
            .O(N__17411),
            .I(N__17408));
    CascadeMux I__3944 (
            .O(N__17408),
            .I(N__17405));
    CascadeBuf I__3943 (
            .O(N__17405),
            .I(N__17402));
    CascadeMux I__3942 (
            .O(N__17402),
            .I(N__17399));
    CascadeBuf I__3941 (
            .O(N__17399),
            .I(N__17396));
    CascadeMux I__3940 (
            .O(N__17396),
            .I(N__17393));
    CascadeBuf I__3939 (
            .O(N__17393),
            .I(N__17390));
    CascadeMux I__3938 (
            .O(N__17390),
            .I(N__17387));
    CascadeBuf I__3937 (
            .O(N__17387),
            .I(N__17384));
    CascadeMux I__3936 (
            .O(N__17384),
            .I(N__17381));
    InMux I__3935 (
            .O(N__17381),
            .I(N__17378));
    LocalMux I__3934 (
            .O(N__17378),
            .I(N__17375));
    Span12Mux_s2_v I__3933 (
            .O(N__17375),
            .I(N__17372));
    Span12Mux_v I__3932 (
            .O(N__17372),
            .I(N__17369));
    Odrv12 I__3931 (
            .O(N__17369),
            .I(M_current_address_qZ0Z_6));
    CEMux I__3930 (
            .O(N__17366),
            .I(N__17363));
    LocalMux I__3929 (
            .O(N__17363),
            .I(N__17359));
    CEMux I__3928 (
            .O(N__17362),
            .I(N__17356));
    Span4Mux_v I__3927 (
            .O(N__17359),
            .I(N__17351));
    LocalMux I__3926 (
            .O(N__17356),
            .I(N__17351));
    Odrv4 I__3925 (
            .O(N__17351),
            .I(\this_vram.mem_WE_4 ));
    InMux I__3924 (
            .O(N__17348),
            .I(N__17341));
    InMux I__3923 (
            .O(N__17347),
            .I(N__17338));
    InMux I__3922 (
            .O(N__17346),
            .I(N__17331));
    InMux I__3921 (
            .O(N__17345),
            .I(N__17331));
    InMux I__3920 (
            .O(N__17344),
            .I(N__17331));
    LocalMux I__3919 (
            .O(N__17341),
            .I(N__17327));
    LocalMux I__3918 (
            .O(N__17338),
            .I(N__17322));
    LocalMux I__3917 (
            .O(N__17331),
            .I(N__17322));
    InMux I__3916 (
            .O(N__17330),
            .I(N__17319));
    Span4Mux_h I__3915 (
            .O(N__17327),
            .I(N__17314));
    Span4Mux_v I__3914 (
            .O(N__17322),
            .I(N__17309));
    LocalMux I__3913 (
            .O(N__17319),
            .I(N__17309));
    InMux I__3912 (
            .O(N__17318),
            .I(N__17304));
    InMux I__3911 (
            .O(N__17317),
            .I(N__17304));
    Odrv4 I__3910 (
            .O(N__17314),
            .I(M_current_address_qZ0Z_12));
    Odrv4 I__3909 (
            .O(N__17309),
            .I(M_current_address_qZ0Z_12));
    LocalMux I__3908 (
            .O(N__17304),
            .I(M_current_address_qZ0Z_12));
    CascadeMux I__3907 (
            .O(N__17297),
            .I(N__17294));
    InMux I__3906 (
            .O(N__17294),
            .I(N__17285));
    CascadeMux I__3905 (
            .O(N__17293),
            .I(N__17281));
    CascadeMux I__3904 (
            .O(N__17292),
            .I(N__17278));
    CascadeMux I__3903 (
            .O(N__17291),
            .I(N__17275));
    CascadeMux I__3902 (
            .O(N__17290),
            .I(N__17272));
    CascadeMux I__3901 (
            .O(N__17289),
            .I(N__17269));
    CascadeMux I__3900 (
            .O(N__17288),
            .I(N__17266));
    LocalMux I__3899 (
            .O(N__17285),
            .I(N__17263));
    CascadeMux I__3898 (
            .O(N__17284),
            .I(N__17260));
    InMux I__3897 (
            .O(N__17281),
            .I(N__17255));
    InMux I__3896 (
            .O(N__17278),
            .I(N__17255));
    InMux I__3895 (
            .O(N__17275),
            .I(N__17252));
    InMux I__3894 (
            .O(N__17272),
            .I(N__17245));
    InMux I__3893 (
            .O(N__17269),
            .I(N__17245));
    InMux I__3892 (
            .O(N__17266),
            .I(N__17245));
    Span4Mux_h I__3891 (
            .O(N__17263),
            .I(N__17242));
    InMux I__3890 (
            .O(N__17260),
            .I(N__17239));
    LocalMux I__3889 (
            .O(N__17255),
            .I(N__17232));
    LocalMux I__3888 (
            .O(N__17252),
            .I(N__17232));
    LocalMux I__3887 (
            .O(N__17245),
            .I(N__17232));
    Odrv4 I__3886 (
            .O(N__17242),
            .I(M_current_address_qZ0Z_13));
    LocalMux I__3885 (
            .O(N__17239),
            .I(M_current_address_qZ0Z_13));
    Odrv12 I__3884 (
            .O(N__17232),
            .I(M_current_address_qZ0Z_13));
    IoInMux I__3883 (
            .O(N__17225),
            .I(N__17222));
    LocalMux I__3882 (
            .O(N__17222),
            .I(N__17219));
    IoSpan4Mux I__3881 (
            .O(N__17219),
            .I(N__17210));
    InMux I__3880 (
            .O(N__17218),
            .I(N__17207));
    InMux I__3879 (
            .O(N__17217),
            .I(N__17202));
    InMux I__3878 (
            .O(N__17216),
            .I(N__17202));
    InMux I__3877 (
            .O(N__17215),
            .I(N__17195));
    InMux I__3876 (
            .O(N__17214),
            .I(N__17195));
    InMux I__3875 (
            .O(N__17213),
            .I(N__17195));
    IoSpan4Mux I__3874 (
            .O(N__17210),
            .I(N__17191));
    LocalMux I__3873 (
            .O(N__17207),
            .I(N__17188));
    LocalMux I__3872 (
            .O(N__17202),
            .I(N__17185));
    LocalMux I__3871 (
            .O(N__17195),
            .I(N__17182));
    InMux I__3870 (
            .O(N__17194),
            .I(N__17179));
    Sp12to4 I__3869 (
            .O(N__17191),
            .I(N__17175));
    Span4Mux_v I__3868 (
            .O(N__17188),
            .I(N__17172));
    Span4Mux_h I__3867 (
            .O(N__17185),
            .I(N__17169));
    Span4Mux_h I__3866 (
            .O(N__17182),
            .I(N__17164));
    LocalMux I__3865 (
            .O(N__17179),
            .I(N__17164));
    InMux I__3864 (
            .O(N__17178),
            .I(N__17161));
    Span12Mux_s9_v I__3863 (
            .O(N__17175),
            .I(N__17157));
    Span4Mux_h I__3862 (
            .O(N__17172),
            .I(N__17154));
    Span4Mux_h I__3861 (
            .O(N__17169),
            .I(N__17151));
    Span4Mux_v I__3860 (
            .O(N__17164),
            .I(N__17146));
    LocalMux I__3859 (
            .O(N__17161),
            .I(N__17146));
    InMux I__3858 (
            .O(N__17160),
            .I(N__17143));
    Odrv12 I__3857 (
            .O(N__17157),
            .I(debug_c));
    Odrv4 I__3856 (
            .O(N__17154),
            .I(debug_c));
    Odrv4 I__3855 (
            .O(N__17151),
            .I(debug_c));
    Odrv4 I__3854 (
            .O(N__17146),
            .I(debug_c));
    LocalMux I__3853 (
            .O(N__17143),
            .I(debug_c));
    CEMux I__3852 (
            .O(N__17132),
            .I(N__17129));
    LocalMux I__3851 (
            .O(N__17129),
            .I(N__17125));
    CEMux I__3850 (
            .O(N__17128),
            .I(N__17122));
    Span4Mux_s2_v I__3849 (
            .O(N__17125),
            .I(N__17117));
    LocalMux I__3848 (
            .O(N__17122),
            .I(N__17117));
    Span4Mux_v I__3847 (
            .O(N__17117),
            .I(N__17114));
    Span4Mux_v I__3846 (
            .O(N__17114),
            .I(N__17111));
    Odrv4 I__3845 (
            .O(N__17111),
            .I(\this_vram.mem_WE_0 ));
    InMux I__3844 (
            .O(N__17108),
            .I(N__17105));
    LocalMux I__3843 (
            .O(N__17105),
            .I(N__17102));
    Span4Mux_v I__3842 (
            .O(N__17102),
            .I(N__17098));
    InMux I__3841 (
            .O(N__17101),
            .I(N__17095));
    Span4Mux_h I__3840 (
            .O(N__17098),
            .I(N__17092));
    LocalMux I__3839 (
            .O(N__17095),
            .I(N__17089));
    Odrv4 I__3838 (
            .O(N__17092),
            .I(port_data_c_5));
    Odrv12 I__3837 (
            .O(N__17089),
            .I(port_data_c_5));
    CascadeMux I__3836 (
            .O(N__17084),
            .I(N__17081));
    CascadeBuf I__3835 (
            .O(N__17081),
            .I(N__17078));
    CascadeMux I__3834 (
            .O(N__17078),
            .I(N__17075));
    CascadeBuf I__3833 (
            .O(N__17075),
            .I(N__17072));
    CascadeMux I__3832 (
            .O(N__17072),
            .I(N__17069));
    CascadeBuf I__3831 (
            .O(N__17069),
            .I(N__17066));
    CascadeMux I__3830 (
            .O(N__17066),
            .I(N__17063));
    CascadeBuf I__3829 (
            .O(N__17063),
            .I(N__17060));
    CascadeMux I__3828 (
            .O(N__17060),
            .I(N__17057));
    CascadeBuf I__3827 (
            .O(N__17057),
            .I(N__17054));
    CascadeMux I__3826 (
            .O(N__17054),
            .I(N__17051));
    CascadeBuf I__3825 (
            .O(N__17051),
            .I(N__17048));
    CascadeMux I__3824 (
            .O(N__17048),
            .I(N__17045));
    CascadeBuf I__3823 (
            .O(N__17045),
            .I(N__17042));
    CascadeMux I__3822 (
            .O(N__17042),
            .I(N__17039));
    CascadeBuf I__3821 (
            .O(N__17039),
            .I(N__17036));
    CascadeMux I__3820 (
            .O(N__17036),
            .I(N__17033));
    CascadeBuf I__3819 (
            .O(N__17033),
            .I(N__17030));
    CascadeMux I__3818 (
            .O(N__17030),
            .I(N__17027));
    CascadeBuf I__3817 (
            .O(N__17027),
            .I(N__17024));
    CascadeMux I__3816 (
            .O(N__17024),
            .I(N__17021));
    CascadeBuf I__3815 (
            .O(N__17021),
            .I(N__17018));
    CascadeMux I__3814 (
            .O(N__17018),
            .I(N__17015));
    CascadeBuf I__3813 (
            .O(N__17015),
            .I(N__17012));
    CascadeMux I__3812 (
            .O(N__17012),
            .I(N__17009));
    CascadeBuf I__3811 (
            .O(N__17009),
            .I(N__17006));
    CascadeMux I__3810 (
            .O(N__17006),
            .I(N__17003));
    CascadeBuf I__3809 (
            .O(N__17003),
            .I(N__17000));
    CascadeMux I__3808 (
            .O(N__17000),
            .I(N__16997));
    CascadeBuf I__3807 (
            .O(N__16997),
            .I(N__16994));
    CascadeMux I__3806 (
            .O(N__16994),
            .I(N__16991));
    InMux I__3805 (
            .O(N__16991),
            .I(N__16988));
    LocalMux I__3804 (
            .O(N__16988),
            .I(N__16985));
    Span4Mux_s1_v I__3803 (
            .O(N__16985),
            .I(N__16982));
    Span4Mux_v I__3802 (
            .O(N__16982),
            .I(N__16979));
    Span4Mux_v I__3801 (
            .O(N__16979),
            .I(N__16976));
    Odrv4 I__3800 (
            .O(N__16976),
            .I(M_current_address_qZ0Z_5));
    InMux I__3799 (
            .O(N__16973),
            .I(N__16969));
    InMux I__3798 (
            .O(N__16972),
            .I(N__16962));
    LocalMux I__3797 (
            .O(N__16969),
            .I(N__16959));
    InMux I__3796 (
            .O(N__16968),
            .I(N__16956));
    InMux I__3795 (
            .O(N__16967),
            .I(N__16947));
    InMux I__3794 (
            .O(N__16966),
            .I(N__16947));
    InMux I__3793 (
            .O(N__16965),
            .I(N__16947));
    LocalMux I__3792 (
            .O(N__16962),
            .I(N__16944));
    Span4Mux_v I__3791 (
            .O(N__16959),
            .I(N__16939));
    LocalMux I__3790 (
            .O(N__16956),
            .I(N__16939));
    InMux I__3789 (
            .O(N__16955),
            .I(N__16934));
    InMux I__3788 (
            .O(N__16954),
            .I(N__16934));
    LocalMux I__3787 (
            .O(N__16947),
            .I(N__16931));
    Span4Mux_h I__3786 (
            .O(N__16944),
            .I(N__16928));
    Span4Mux_v I__3785 (
            .O(N__16939),
            .I(N__16923));
    LocalMux I__3784 (
            .O(N__16934),
            .I(N__16923));
    Odrv12 I__3783 (
            .O(N__16931),
            .I(M_current_address_qZ0Z_11));
    Odrv4 I__3782 (
            .O(N__16928),
            .I(M_current_address_qZ0Z_11));
    Odrv4 I__3781 (
            .O(N__16923),
            .I(M_current_address_qZ0Z_11));
    InMux I__3780 (
            .O(N__16916),
            .I(N__16913));
    LocalMux I__3779 (
            .O(N__16913),
            .I(N__16909));
    InMux I__3778 (
            .O(N__16912),
            .I(N__16906));
    Span4Mux_v I__3777 (
            .O(N__16909),
            .I(N__16901));
    LocalMux I__3776 (
            .O(N__16906),
            .I(N__16901));
    Span4Mux_h I__3775 (
            .O(N__16901),
            .I(N__16898));
    Span4Mux_v I__3774 (
            .O(N__16898),
            .I(N__16895));
    Span4Mux_h I__3773 (
            .O(N__16895),
            .I(N__16892));
    Odrv4 I__3772 (
            .O(N__16892),
            .I(port_data_c_4));
    CascadeMux I__3771 (
            .O(N__16889),
            .I(N__16886));
    CascadeBuf I__3770 (
            .O(N__16886),
            .I(N__16883));
    CascadeMux I__3769 (
            .O(N__16883),
            .I(N__16880));
    CascadeBuf I__3768 (
            .O(N__16880),
            .I(N__16877));
    CascadeMux I__3767 (
            .O(N__16877),
            .I(N__16874));
    CascadeBuf I__3766 (
            .O(N__16874),
            .I(N__16871));
    CascadeMux I__3765 (
            .O(N__16871),
            .I(N__16868));
    CascadeBuf I__3764 (
            .O(N__16868),
            .I(N__16865));
    CascadeMux I__3763 (
            .O(N__16865),
            .I(N__16862));
    CascadeBuf I__3762 (
            .O(N__16862),
            .I(N__16859));
    CascadeMux I__3761 (
            .O(N__16859),
            .I(N__16856));
    CascadeBuf I__3760 (
            .O(N__16856),
            .I(N__16853));
    CascadeMux I__3759 (
            .O(N__16853),
            .I(N__16850));
    CascadeBuf I__3758 (
            .O(N__16850),
            .I(N__16847));
    CascadeMux I__3757 (
            .O(N__16847),
            .I(N__16844));
    CascadeBuf I__3756 (
            .O(N__16844),
            .I(N__16841));
    CascadeMux I__3755 (
            .O(N__16841),
            .I(N__16838));
    CascadeBuf I__3754 (
            .O(N__16838),
            .I(N__16835));
    CascadeMux I__3753 (
            .O(N__16835),
            .I(N__16832));
    CascadeBuf I__3752 (
            .O(N__16832),
            .I(N__16829));
    CascadeMux I__3751 (
            .O(N__16829),
            .I(N__16826));
    CascadeBuf I__3750 (
            .O(N__16826),
            .I(N__16823));
    CascadeMux I__3749 (
            .O(N__16823),
            .I(N__16820));
    CascadeBuf I__3748 (
            .O(N__16820),
            .I(N__16817));
    CascadeMux I__3747 (
            .O(N__16817),
            .I(N__16814));
    CascadeBuf I__3746 (
            .O(N__16814),
            .I(N__16811));
    CascadeMux I__3745 (
            .O(N__16811),
            .I(N__16808));
    CascadeBuf I__3744 (
            .O(N__16808),
            .I(N__16805));
    CascadeMux I__3743 (
            .O(N__16805),
            .I(N__16802));
    CascadeBuf I__3742 (
            .O(N__16802),
            .I(N__16799));
    CascadeMux I__3741 (
            .O(N__16799),
            .I(N__16796));
    InMux I__3740 (
            .O(N__16796),
            .I(N__16793));
    LocalMux I__3739 (
            .O(N__16793),
            .I(N__16790));
    Span4Mux_s2_v I__3738 (
            .O(N__16790),
            .I(N__16787));
    Span4Mux_v I__3737 (
            .O(N__16787),
            .I(N__16784));
    Odrv4 I__3736 (
            .O(N__16784),
            .I(M_current_address_qZ0Z_4));
    CascadeMux I__3735 (
            .O(N__16781),
            .I(\this_vram.mem_mem_1_1_RNIUSK11Z0Z_0_cascade_ ));
    InMux I__3734 (
            .O(N__16778),
            .I(N__16775));
    LocalMux I__3733 (
            .O(N__16775),
            .I(N__16772));
    Span4Mux_h I__3732 (
            .O(N__16772),
            .I(N__16769));
    Odrv4 I__3731 (
            .O(N__16769),
            .I(\this_vram.mem_N_102 ));
    InMux I__3730 (
            .O(N__16766),
            .I(N__16763));
    LocalMux I__3729 (
            .O(N__16763),
            .I(N__16760));
    Span4Mux_v I__3728 (
            .O(N__16760),
            .I(N__16757));
    Span4Mux_v I__3727 (
            .O(N__16757),
            .I(N__16754));
    Odrv4 I__3726 (
            .O(N__16754),
            .I(\this_vram.mem_out_bus1_2 ));
    InMux I__3725 (
            .O(N__16751),
            .I(N__16748));
    LocalMux I__3724 (
            .O(N__16748),
            .I(N__16745));
    Sp12to4 I__3723 (
            .O(N__16745),
            .I(N__16742));
    Span12Mux_v I__3722 (
            .O(N__16742),
            .I(N__16739));
    Odrv12 I__3721 (
            .O(N__16739),
            .I(\this_vram.mem_out_bus5_2 ));
    InMux I__3720 (
            .O(N__16736),
            .I(N__16725));
    InMux I__3719 (
            .O(N__16735),
            .I(N__16725));
    InMux I__3718 (
            .O(N__16734),
            .I(N__16722));
    InMux I__3717 (
            .O(N__16733),
            .I(N__16717));
    InMux I__3716 (
            .O(N__16732),
            .I(N__16717));
    InMux I__3715 (
            .O(N__16731),
            .I(N__16712));
    InMux I__3714 (
            .O(N__16730),
            .I(N__16712));
    LocalMux I__3713 (
            .O(N__16725),
            .I(N__16704));
    LocalMux I__3712 (
            .O(N__16722),
            .I(N__16704));
    LocalMux I__3711 (
            .O(N__16717),
            .I(N__16704));
    LocalMux I__3710 (
            .O(N__16712),
            .I(N__16701));
    InMux I__3709 (
            .O(N__16711),
            .I(N__16698));
    Span4Mux_v I__3708 (
            .O(N__16704),
            .I(N__16691));
    Span4Mux_v I__3707 (
            .O(N__16701),
            .I(N__16691));
    LocalMux I__3706 (
            .O(N__16698),
            .I(N__16691));
    Odrv4 I__3705 (
            .O(N__16691),
            .I(\this_vram.mem_radregZ0Z_12 ));
    CascadeMux I__3704 (
            .O(N__16688),
            .I(\this_vram.mem_mem_1_1_RNIUSKZ0Z11_cascade_ ));
    InMux I__3703 (
            .O(N__16685),
            .I(N__16682));
    LocalMux I__3702 (
            .O(N__16682),
            .I(\this_vram.mem_N_95 ));
    InMux I__3701 (
            .O(N__16679),
            .I(N__16676));
    LocalMux I__3700 (
            .O(N__16676),
            .I(N__16673));
    Span4Mux_h I__3699 (
            .O(N__16673),
            .I(N__16670));
    Odrv4 I__3698 (
            .O(N__16670),
            .I(\this_vram.mem_out_bus3_0 ));
    InMux I__3697 (
            .O(N__16667),
            .I(N__16664));
    LocalMux I__3696 (
            .O(N__16664),
            .I(N__16661));
    Sp12to4 I__3695 (
            .O(N__16661),
            .I(N__16658));
    Span12Mux_v I__3694 (
            .O(N__16658),
            .I(N__16655));
    Odrv12 I__3693 (
            .O(N__16655),
            .I(\this_vram.mem_out_bus7_0 ));
    InMux I__3692 (
            .O(N__16652),
            .I(N__16649));
    LocalMux I__3691 (
            .O(N__16649),
            .I(N__16646));
    Span4Mux_v I__3690 (
            .O(N__16646),
            .I(N__16643));
    Odrv4 I__3689 (
            .O(N__16643),
            .I(\this_vram.mem_mem_3_0_RNI05PZ0Z11 ));
    CEMux I__3688 (
            .O(N__16640),
            .I(N__16637));
    LocalMux I__3687 (
            .O(N__16637),
            .I(N__16633));
    CEMux I__3686 (
            .O(N__16636),
            .I(N__16630));
    Span4Mux_v I__3685 (
            .O(N__16633),
            .I(N__16625));
    LocalMux I__3684 (
            .O(N__16630),
            .I(N__16625));
    Span4Mux_h I__3683 (
            .O(N__16625),
            .I(N__16622));
    Odrv4 I__3682 (
            .O(N__16622),
            .I(\this_vram.mem_WE_10 ));
    CEMux I__3681 (
            .O(N__16619),
            .I(N__16616));
    LocalMux I__3680 (
            .O(N__16616),
            .I(N__16613));
    Span12Mux_s8_h I__3679 (
            .O(N__16613),
            .I(N__16609));
    CEMux I__3678 (
            .O(N__16612),
            .I(N__16606));
    Odrv12 I__3677 (
            .O(N__16609),
            .I(\this_vram.mem_WE_8 ));
    LocalMux I__3676 (
            .O(N__16606),
            .I(\this_vram.mem_WE_8 ));
    CEMux I__3675 (
            .O(N__16601),
            .I(N__16598));
    LocalMux I__3674 (
            .O(N__16598),
            .I(N__16594));
    CEMux I__3673 (
            .O(N__16597),
            .I(N__16591));
    Span4Mux_s1_v I__3672 (
            .O(N__16594),
            .I(N__16586));
    LocalMux I__3671 (
            .O(N__16591),
            .I(N__16586));
    Span4Mux_v I__3670 (
            .O(N__16586),
            .I(N__16583));
    Span4Mux_v I__3669 (
            .O(N__16583),
            .I(N__16580));
    Odrv4 I__3668 (
            .O(N__16580),
            .I(\this_vram.mem_WE_14 ));
    InMux I__3667 (
            .O(N__16577),
            .I(N__16574));
    LocalMux I__3666 (
            .O(N__16574),
            .I(N__16571));
    Span4Mux_v I__3665 (
            .O(N__16571),
            .I(N__16568));
    Span4Mux_v I__3664 (
            .O(N__16568),
            .I(N__16565));
    Sp12to4 I__3663 (
            .O(N__16565),
            .I(N__16562));
    Odrv12 I__3662 (
            .O(N__16562),
            .I(\this_vram.mem_out_bus7_3 ));
    InMux I__3661 (
            .O(N__16559),
            .I(N__16556));
    LocalMux I__3660 (
            .O(N__16556),
            .I(\this_vram.mem_out_bus3_3 ));
    InMux I__3659 (
            .O(N__16553),
            .I(N__16550));
    LocalMux I__3658 (
            .O(N__16550),
            .I(N__16547));
    Odrv4 I__3657 (
            .O(N__16547),
            .I(\this_vram.mem_mem_3_1_RNI25P11Z0Z_0 ));
    InMux I__3656 (
            .O(N__16544),
            .I(N__16541));
    LocalMux I__3655 (
            .O(N__16541),
            .I(\this_vram.mem_out_bus3_2 ));
    InMux I__3654 (
            .O(N__16538),
            .I(N__16535));
    LocalMux I__3653 (
            .O(N__16535),
            .I(N__16532));
    Span4Mux_v I__3652 (
            .O(N__16532),
            .I(N__16529));
    Span4Mux_v I__3651 (
            .O(N__16529),
            .I(N__16526));
    Sp12to4 I__3650 (
            .O(N__16526),
            .I(N__16523));
    Odrv12 I__3649 (
            .O(N__16523),
            .I(\this_vram.mem_out_bus7_2 ));
    InMux I__3648 (
            .O(N__16520),
            .I(N__16516));
    InMux I__3647 (
            .O(N__16519),
            .I(N__16509));
    LocalMux I__3646 (
            .O(N__16516),
            .I(N__16502));
    InMux I__3645 (
            .O(N__16515),
            .I(N__16497));
    InMux I__3644 (
            .O(N__16514),
            .I(N__16497));
    InMux I__3643 (
            .O(N__16513),
            .I(N__16492));
    InMux I__3642 (
            .O(N__16512),
            .I(N__16492));
    LocalMux I__3641 (
            .O(N__16509),
            .I(N__16489));
    InMux I__3640 (
            .O(N__16508),
            .I(N__16480));
    InMux I__3639 (
            .O(N__16507),
            .I(N__16480));
    InMux I__3638 (
            .O(N__16506),
            .I(N__16480));
    InMux I__3637 (
            .O(N__16505),
            .I(N__16480));
    Span4Mux_v I__3636 (
            .O(N__16502),
            .I(N__16469));
    LocalMux I__3635 (
            .O(N__16497),
            .I(N__16469));
    LocalMux I__3634 (
            .O(N__16492),
            .I(N__16466));
    Span4Mux_v I__3633 (
            .O(N__16489),
            .I(N__16461));
    LocalMux I__3632 (
            .O(N__16480),
            .I(N__16461));
    InMux I__3631 (
            .O(N__16479),
            .I(N__16452));
    InMux I__3630 (
            .O(N__16478),
            .I(N__16452));
    InMux I__3629 (
            .O(N__16477),
            .I(N__16452));
    InMux I__3628 (
            .O(N__16476),
            .I(N__16452));
    InMux I__3627 (
            .O(N__16475),
            .I(N__16447));
    InMux I__3626 (
            .O(N__16474),
            .I(N__16447));
    Odrv4 I__3625 (
            .O(N__16469),
            .I(\this_vram.mem_radregZ0Z_13 ));
    Odrv4 I__3624 (
            .O(N__16466),
            .I(\this_vram.mem_radregZ0Z_13 ));
    Odrv4 I__3623 (
            .O(N__16461),
            .I(\this_vram.mem_radregZ0Z_13 ));
    LocalMux I__3622 (
            .O(N__16452),
            .I(\this_vram.mem_radregZ0Z_13 ));
    LocalMux I__3621 (
            .O(N__16447),
            .I(\this_vram.mem_radregZ0Z_13 ));
    InMux I__3620 (
            .O(N__16436),
            .I(N__16433));
    LocalMux I__3619 (
            .O(N__16433),
            .I(N__16430));
    Odrv12 I__3618 (
            .O(N__16430),
            .I(\this_vram.mem_mem_3_1_RNI25PZ0Z11 ));
    CascadeMux I__3617 (
            .O(N__16427),
            .I(\this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_ ));
    InMux I__3616 (
            .O(N__16424),
            .I(N__16421));
    LocalMux I__3615 (
            .O(N__16421),
            .I(\this_vram.mem_mem_2_0_RNIU0N11Z0Z_0 ));
    InMux I__3614 (
            .O(N__16418),
            .I(N__16415));
    LocalMux I__3613 (
            .O(N__16415),
            .I(N__16412));
    Span4Mux_v I__3612 (
            .O(N__16412),
            .I(N__16409));
    Odrv4 I__3611 (
            .O(N__16409),
            .I(\this_vram.mem_N_91 ));
    InMux I__3610 (
            .O(N__16406),
            .I(N__16402));
    InMux I__3609 (
            .O(N__16405),
            .I(N__16398));
    LocalMux I__3608 (
            .O(N__16402),
            .I(N__16395));
    InMux I__3607 (
            .O(N__16401),
            .I(N__16392));
    LocalMux I__3606 (
            .O(N__16398),
            .I(N__16387));
    Span4Mux_h I__3605 (
            .O(N__16395),
            .I(N__16387));
    LocalMux I__3604 (
            .O(N__16392),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKMEZ0 ));
    Odrv4 I__3603 (
            .O(N__16387),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKMEZ0 ));
    CascadeMux I__3602 (
            .O(N__16382),
            .I(N__16379));
    InMux I__3601 (
            .O(N__16379),
            .I(N__16372));
    InMux I__3600 (
            .O(N__16378),
            .I(N__16372));
    CascadeMux I__3599 (
            .O(N__16377),
            .I(N__16366));
    LocalMux I__3598 (
            .O(N__16372),
            .I(N__16360));
    InMux I__3597 (
            .O(N__16371),
            .I(N__16357));
    InMux I__3596 (
            .O(N__16370),
            .I(N__16353));
    InMux I__3595 (
            .O(N__16369),
            .I(N__16350));
    InMux I__3594 (
            .O(N__16366),
            .I(N__16342));
    InMux I__3593 (
            .O(N__16365),
            .I(N__16339));
    InMux I__3592 (
            .O(N__16364),
            .I(N__16334));
    InMux I__3591 (
            .O(N__16363),
            .I(N__16334));
    Span4Mux_v I__3590 (
            .O(N__16360),
            .I(N__16329));
    LocalMux I__3589 (
            .O(N__16357),
            .I(N__16329));
    InMux I__3588 (
            .O(N__16356),
            .I(N__16326));
    LocalMux I__3587 (
            .O(N__16353),
            .I(N__16321));
    LocalMux I__3586 (
            .O(N__16350),
            .I(N__16321));
    InMux I__3585 (
            .O(N__16349),
            .I(N__16314));
    InMux I__3584 (
            .O(N__16348),
            .I(N__16314));
    InMux I__3583 (
            .O(N__16347),
            .I(N__16314));
    InMux I__3582 (
            .O(N__16346),
            .I(N__16311));
    InMux I__3581 (
            .O(N__16345),
            .I(N__16305));
    LocalMux I__3580 (
            .O(N__16342),
            .I(N__16300));
    LocalMux I__3579 (
            .O(N__16339),
            .I(N__16300));
    LocalMux I__3578 (
            .O(N__16334),
            .I(N__16297));
    Span4Mux_h I__3577 (
            .O(N__16329),
            .I(N__16294));
    LocalMux I__3576 (
            .O(N__16326),
            .I(N__16290));
    Span4Mux_v I__3575 (
            .O(N__16321),
            .I(N__16285));
    LocalMux I__3574 (
            .O(N__16314),
            .I(N__16285));
    LocalMux I__3573 (
            .O(N__16311),
            .I(N__16282));
    InMux I__3572 (
            .O(N__16310),
            .I(N__16275));
    InMux I__3571 (
            .O(N__16309),
            .I(N__16275));
    InMux I__3570 (
            .O(N__16308),
            .I(N__16275));
    LocalMux I__3569 (
            .O(N__16305),
            .I(N__16272));
    Span4Mux_v I__3568 (
            .O(N__16300),
            .I(N__16267));
    Span4Mux_v I__3567 (
            .O(N__16297),
            .I(N__16267));
    Span4Mux_h I__3566 (
            .O(N__16294),
            .I(N__16264));
    InMux I__3565 (
            .O(N__16293),
            .I(N__16261));
    Span4Mux_v I__3564 (
            .O(N__16290),
            .I(N__16252));
    Span4Mux_h I__3563 (
            .O(N__16285),
            .I(N__16252));
    Span4Mux_v I__3562 (
            .O(N__16282),
            .I(N__16252));
    LocalMux I__3561 (
            .O(N__16275),
            .I(N__16252));
    Odrv4 I__3560 (
            .O(N__16272),
            .I(\this_vga_signals.M_vaddress_qZ0Z_5 ));
    Odrv4 I__3559 (
            .O(N__16267),
            .I(\this_vga_signals.M_vaddress_qZ0Z_5 ));
    Odrv4 I__3558 (
            .O(N__16264),
            .I(\this_vga_signals.M_vaddress_qZ0Z_5 ));
    LocalMux I__3557 (
            .O(N__16261),
            .I(\this_vga_signals.M_vaddress_qZ0Z_5 ));
    Odrv4 I__3556 (
            .O(N__16252),
            .I(\this_vga_signals.M_vaddress_qZ0Z_5 ));
    SRMux I__3555 (
            .O(N__16241),
            .I(N__16220));
    SRMux I__3554 (
            .O(N__16240),
            .I(N__16220));
    SRMux I__3553 (
            .O(N__16239),
            .I(N__16220));
    SRMux I__3552 (
            .O(N__16238),
            .I(N__16220));
    SRMux I__3551 (
            .O(N__16237),
            .I(N__16220));
    SRMux I__3550 (
            .O(N__16236),
            .I(N__16220));
    SRMux I__3549 (
            .O(N__16235),
            .I(N__16220));
    GlobalMux I__3548 (
            .O(N__16220),
            .I(N__16217));
    gio2CtrlBuf I__3547 (
            .O(N__16217),
            .I(\this_vga_signals.N_583_g ));
    InMux I__3546 (
            .O(N__16214),
            .I(N__16211));
    LocalMux I__3545 (
            .O(N__16211),
            .I(N__16208));
    Sp12to4 I__3544 (
            .O(N__16208),
            .I(N__16205));
    Span12Mux_v I__3543 (
            .O(N__16205),
            .I(N__16202));
    Span12Mux_v I__3542 (
            .O(N__16202),
            .I(N__16199));
    Odrv12 I__3541 (
            .O(N__16199),
            .I(\this_vram.mem_out_bus6_3 ));
    InMux I__3540 (
            .O(N__16196),
            .I(N__16193));
    LocalMux I__3539 (
            .O(N__16193),
            .I(\this_vram.mem_out_bus2_3 ));
    CascadeMux I__3538 (
            .O(N__16190),
            .I(\this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_ ));
    InMux I__3537 (
            .O(N__16187),
            .I(N__16184));
    LocalMux I__3536 (
            .O(N__16184),
            .I(N__16181));
    Span4Mux_h I__3535 (
            .O(N__16181),
            .I(N__16178));
    Odrv4 I__3534 (
            .O(N__16178),
            .I(\this_vram.mem_N_105 ));
    InMux I__3533 (
            .O(N__16175),
            .I(N__16172));
    LocalMux I__3532 (
            .O(N__16172),
            .I(N__16169));
    Span4Mux_v I__3531 (
            .O(N__16169),
            .I(N__16166));
    Span4Mux_v I__3530 (
            .O(N__16166),
            .I(N__16163));
    Odrv4 I__3529 (
            .O(N__16163),
            .I(\this_vram.mem_out_bus0_3 ));
    InMux I__3528 (
            .O(N__16160),
            .I(N__16157));
    LocalMux I__3527 (
            .O(N__16157),
            .I(N__16154));
    Span4Mux_v I__3526 (
            .O(N__16154),
            .I(N__16151));
    Odrv4 I__3525 (
            .O(N__16151),
            .I(\this_vram.mem_out_bus4_3 ));
    InMux I__3524 (
            .O(N__16148),
            .I(N__16145));
    LocalMux I__3523 (
            .O(N__16145),
            .I(\this_vram.mem_mem_0_1_RNISOI11Z0Z_0 ));
    CEMux I__3522 (
            .O(N__16142),
            .I(N__16139));
    LocalMux I__3521 (
            .O(N__16139),
            .I(N__16135));
    CEMux I__3520 (
            .O(N__16138),
            .I(N__16132));
    Span4Mux_v I__3519 (
            .O(N__16135),
            .I(N__16127));
    LocalMux I__3518 (
            .O(N__16132),
            .I(N__16127));
    Span4Mux_v I__3517 (
            .O(N__16127),
            .I(N__16124));
    Odrv4 I__3516 (
            .O(N__16124),
            .I(\this_vram.mem_WE_12 ));
    InMux I__3515 (
            .O(N__16121),
            .I(N__16118));
    LocalMux I__3514 (
            .O(N__16118),
            .I(N__16115));
    Span4Mux_v I__3513 (
            .O(N__16115),
            .I(N__16112));
    Span4Mux_v I__3512 (
            .O(N__16112),
            .I(N__16109));
    Sp12to4 I__3511 (
            .O(N__16109),
            .I(N__16106));
    Odrv12 I__3510 (
            .O(N__16106),
            .I(\this_vram.mem_out_bus7_1 ));
    InMux I__3509 (
            .O(N__16103),
            .I(N__16100));
    LocalMux I__3508 (
            .O(N__16100),
            .I(\this_vram.mem_out_bus3_1 ));
    InMux I__3507 (
            .O(N__16097),
            .I(N__16094));
    LocalMux I__3506 (
            .O(N__16094),
            .I(N__16091));
    Odrv12 I__3505 (
            .O(N__16091),
            .I(\this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ));
    InMux I__3504 (
            .O(N__16088),
            .I(N__16085));
    LocalMux I__3503 (
            .O(N__16085),
            .I(N__16082));
    Sp12to4 I__3502 (
            .O(N__16082),
            .I(N__16079));
    Span12Mux_v I__3501 (
            .O(N__16079),
            .I(N__16076));
    Odrv12 I__3500 (
            .O(N__16076),
            .I(\this_vram.mem_out_bus5_3 ));
    InMux I__3499 (
            .O(N__16073),
            .I(N__16070));
    LocalMux I__3498 (
            .O(N__16070),
            .I(N__16067));
    Span4Mux_v I__3497 (
            .O(N__16067),
            .I(N__16064));
    Odrv4 I__3496 (
            .O(N__16064),
            .I(\this_vram.mem_out_bus1_3 ));
    CascadeMux I__3495 (
            .O(N__16061),
            .I(N__16058));
    InMux I__3494 (
            .O(N__16058),
            .I(N__16055));
    LocalMux I__3493 (
            .O(N__16055),
            .I(\this_vram.mem_out_bus2_0 ));
    InMux I__3492 (
            .O(N__16052),
            .I(N__16049));
    LocalMux I__3491 (
            .O(N__16049),
            .I(N__16046));
    Span4Mux_v I__3490 (
            .O(N__16046),
            .I(N__16043));
    Span4Mux_v I__3489 (
            .O(N__16043),
            .I(N__16040));
    Sp12to4 I__3488 (
            .O(N__16040),
            .I(N__16037));
    Odrv12 I__3487 (
            .O(N__16037),
            .I(\this_vram.mem_out_bus6_0 ));
    InMux I__3486 (
            .O(N__16034),
            .I(N__16031));
    LocalMux I__3485 (
            .O(N__16031),
            .I(\this_vram.mem_mem_2_0_RNIU0NZ0Z11 ));
    InMux I__3484 (
            .O(N__16028),
            .I(N__16025));
    LocalMux I__3483 (
            .O(N__16025),
            .I(N__16022));
    Span4Mux_v I__3482 (
            .O(N__16022),
            .I(N__16019));
    Odrv4 I__3481 (
            .O(N__16019),
            .I(\this_vram.mem_out_bus1_1 ));
    InMux I__3480 (
            .O(N__16016),
            .I(N__16013));
    LocalMux I__3479 (
            .O(N__16013),
            .I(N__16010));
    Sp12to4 I__3478 (
            .O(N__16010),
            .I(N__16007));
    Span12Mux_v I__3477 (
            .O(N__16007),
            .I(N__16004));
    Odrv12 I__3476 (
            .O(N__16004),
            .I(\this_vram.mem_out_bus5_1 ));
    CascadeMux I__3475 (
            .O(N__16001),
            .I(\this_vram.mem_mem_1_0_RNISSK11Z0Z_0_cascade_ ));
    InMux I__3474 (
            .O(N__15998),
            .I(N__15995));
    LocalMux I__3473 (
            .O(N__15995),
            .I(N__15992));
    Odrv4 I__3472 (
            .O(N__15992),
            .I(\this_vram.mem_N_88 ));
    InMux I__3471 (
            .O(N__15989),
            .I(N__15986));
    LocalMux I__3470 (
            .O(N__15986),
            .I(N__15983));
    Sp12to4 I__3469 (
            .O(N__15983),
            .I(N__15980));
    Span12Mux_v I__3468 (
            .O(N__15980),
            .I(N__15977));
    Odrv12 I__3467 (
            .O(N__15977),
            .I(\this_vram.mem_out_bus4_2 ));
    InMux I__3466 (
            .O(N__15974),
            .I(N__15971));
    LocalMux I__3465 (
            .O(N__15971),
            .I(N__15968));
    Span4Mux_v I__3464 (
            .O(N__15968),
            .I(N__15965));
    Odrv4 I__3463 (
            .O(N__15965),
            .I(\this_vram.mem_out_bus0_2 ));
    InMux I__3462 (
            .O(N__15962),
            .I(N__15959));
    LocalMux I__3461 (
            .O(N__15959),
            .I(N__15956));
    Sp12to4 I__3460 (
            .O(N__15956),
            .I(N__15953));
    Span12Mux_v I__3459 (
            .O(N__15953),
            .I(N__15950));
    Span12Mux_v I__3458 (
            .O(N__15950),
            .I(N__15947));
    Odrv12 I__3457 (
            .O(N__15947),
            .I(\this_vram.mem_out_bus6_2 ));
    InMux I__3456 (
            .O(N__15944),
            .I(N__15941));
    LocalMux I__3455 (
            .O(N__15941),
            .I(N__15938));
    Odrv4 I__3454 (
            .O(N__15938),
            .I(\this_vram.mem_out_bus2_2 ));
    InMux I__3453 (
            .O(N__15935),
            .I(N__15932));
    LocalMux I__3452 (
            .O(N__15932),
            .I(\this_vram.mem_mem_0_1_RNISOIZ0Z11 ));
    CascadeMux I__3451 (
            .O(N__15929),
            .I(\this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_ ));
    InMux I__3450 (
            .O(N__15926),
            .I(N__15923));
    LocalMux I__3449 (
            .O(N__15923),
            .I(N__15920));
    Odrv4 I__3448 (
            .O(N__15920),
            .I(\this_vram.mem_N_98 ));
    InMux I__3447 (
            .O(N__15917),
            .I(N__15914));
    LocalMux I__3446 (
            .O(N__15914),
            .I(N__15911));
    Sp12to4 I__3445 (
            .O(N__15911),
            .I(N__15908));
    Span12Mux_v I__3444 (
            .O(N__15908),
            .I(N__15905));
    Odrv12 I__3443 (
            .O(N__15905),
            .I(\this_vram.mem_out_bus6_1 ));
    InMux I__3442 (
            .O(N__15902),
            .I(N__15899));
    LocalMux I__3441 (
            .O(N__15899),
            .I(\this_vram.mem_out_bus2_1 ));
    InMux I__3440 (
            .O(N__15896),
            .I(N__15893));
    LocalMux I__3439 (
            .O(N__15893),
            .I(N__15890));
    Span4Mux_v I__3438 (
            .O(N__15890),
            .I(N__15887));
    Odrv4 I__3437 (
            .O(N__15887),
            .I(\this_vram.mem_out_bus4_1 ));
    InMux I__3436 (
            .O(N__15884),
            .I(N__15881));
    LocalMux I__3435 (
            .O(N__15881),
            .I(N__15878));
    Span4Mux_v I__3434 (
            .O(N__15878),
            .I(N__15875));
    Span4Mux_v I__3433 (
            .O(N__15875),
            .I(N__15872));
    Odrv4 I__3432 (
            .O(N__15872),
            .I(\this_vram.mem_out_bus0_1 ));
    CascadeMux I__3431 (
            .O(N__15869),
            .I(N__15866));
    InMux I__3430 (
            .O(N__15866),
            .I(N__15860));
    InMux I__3429 (
            .O(N__15865),
            .I(N__15857));
    InMux I__3428 (
            .O(N__15864),
            .I(N__15852));
    CascadeMux I__3427 (
            .O(N__15863),
            .I(N__15849));
    LocalMux I__3426 (
            .O(N__15860),
            .I(N__15844));
    LocalMux I__3425 (
            .O(N__15857),
            .I(N__15844));
    InMux I__3424 (
            .O(N__15856),
            .I(N__15841));
    CascadeMux I__3423 (
            .O(N__15855),
            .I(N__15838));
    LocalMux I__3422 (
            .O(N__15852),
            .I(N__15835));
    InMux I__3421 (
            .O(N__15849),
            .I(N__15832));
    Span4Mux_v I__3420 (
            .O(N__15844),
            .I(N__15827));
    LocalMux I__3419 (
            .O(N__15841),
            .I(N__15827));
    InMux I__3418 (
            .O(N__15838),
            .I(N__15824));
    Span4Mux_v I__3417 (
            .O(N__15835),
            .I(N__15821));
    LocalMux I__3416 (
            .O(N__15832),
            .I(N__15814));
    Sp12to4 I__3415 (
            .O(N__15827),
            .I(N__15814));
    LocalMux I__3414 (
            .O(N__15824),
            .I(N__15814));
    Sp12to4 I__3413 (
            .O(N__15821),
            .I(N__15811));
    Span12Mux_v I__3412 (
            .O(N__15814),
            .I(N__15808));
    Span12Mux_h I__3411 (
            .O(N__15811),
            .I(N__15803));
    Span12Mux_h I__3410 (
            .O(N__15808),
            .I(N__15803));
    Odrv12 I__3409 (
            .O(N__15803),
            .I(M_this_vram_read_data_2));
    CEMux I__3408 (
            .O(N__15800),
            .I(N__15796));
    CEMux I__3407 (
            .O(N__15799),
            .I(N__15793));
    LocalMux I__3406 (
            .O(N__15796),
            .I(N__15788));
    LocalMux I__3405 (
            .O(N__15793),
            .I(N__15788));
    Span4Mux_v I__3404 (
            .O(N__15788),
            .I(N__15785));
    Span4Mux_h I__3403 (
            .O(N__15785),
            .I(N__15782));
    Odrv4 I__3402 (
            .O(N__15782),
            .I(\this_vram.mem_WE_6 ));
    InMux I__3401 (
            .O(N__15779),
            .I(N__15776));
    LocalMux I__3400 (
            .O(N__15776),
            .I(N__15773));
    Odrv4 I__3399 (
            .O(N__15773),
            .I(M_current_address_qZ1Z_0));
    CascadeMux I__3398 (
            .O(N__15770),
            .I(N__15767));
    CascadeBuf I__3397 (
            .O(N__15767),
            .I(N__15764));
    CascadeMux I__3396 (
            .O(N__15764),
            .I(N__15761));
    CascadeBuf I__3395 (
            .O(N__15761),
            .I(N__15758));
    CascadeMux I__3394 (
            .O(N__15758),
            .I(N__15755));
    CascadeBuf I__3393 (
            .O(N__15755),
            .I(N__15752));
    CascadeMux I__3392 (
            .O(N__15752),
            .I(N__15749));
    CascadeBuf I__3391 (
            .O(N__15749),
            .I(N__15746));
    CascadeMux I__3390 (
            .O(N__15746),
            .I(N__15743));
    CascadeBuf I__3389 (
            .O(N__15743),
            .I(N__15740));
    CascadeMux I__3388 (
            .O(N__15740),
            .I(N__15737));
    CascadeBuf I__3387 (
            .O(N__15737),
            .I(N__15734));
    CascadeMux I__3386 (
            .O(N__15734),
            .I(N__15731));
    CascadeBuf I__3385 (
            .O(N__15731),
            .I(N__15728));
    CascadeMux I__3384 (
            .O(N__15728),
            .I(N__15725));
    CascadeBuf I__3383 (
            .O(N__15725),
            .I(N__15722));
    CascadeMux I__3382 (
            .O(N__15722),
            .I(N__15719));
    CascadeBuf I__3381 (
            .O(N__15719),
            .I(N__15716));
    CascadeMux I__3380 (
            .O(N__15716),
            .I(N__15713));
    CascadeBuf I__3379 (
            .O(N__15713),
            .I(N__15710));
    CascadeMux I__3378 (
            .O(N__15710),
            .I(N__15707));
    CascadeBuf I__3377 (
            .O(N__15707),
            .I(N__15704));
    CascadeMux I__3376 (
            .O(N__15704),
            .I(N__15701));
    CascadeBuf I__3375 (
            .O(N__15701),
            .I(N__15698));
    CascadeMux I__3374 (
            .O(N__15698),
            .I(N__15695));
    CascadeBuf I__3373 (
            .O(N__15695),
            .I(N__15692));
    CascadeMux I__3372 (
            .O(N__15692),
            .I(N__15689));
    CascadeBuf I__3371 (
            .O(N__15689),
            .I(N__15686));
    CascadeMux I__3370 (
            .O(N__15686),
            .I(N__15683));
    CascadeBuf I__3369 (
            .O(N__15683),
            .I(N__15680));
    CascadeMux I__3368 (
            .O(N__15680),
            .I(N__15677));
    InMux I__3367 (
            .O(N__15677),
            .I(N__15674));
    LocalMux I__3366 (
            .O(N__15674),
            .I(N__15671));
    Span4Mux_s1_v I__3365 (
            .O(N__15671),
            .I(N__15668));
    Span4Mux_v I__3364 (
            .O(N__15668),
            .I(N__15665));
    Odrv4 I__3363 (
            .O(N__15665),
            .I(M_current_address_qZ0Z_0));
    InMux I__3362 (
            .O(N__15662),
            .I(N__15659));
    LocalMux I__3361 (
            .O(N__15659),
            .I(N__15656));
    Span4Mux_v I__3360 (
            .O(N__15656),
            .I(N__15653));
    Span4Mux_v I__3359 (
            .O(N__15653),
            .I(N__15650));
    Span4Mux_v I__3358 (
            .O(N__15650),
            .I(N__15647));
    Odrv4 I__3357 (
            .O(N__15647),
            .I(\this_vram.mem_out_bus5_0 ));
    InMux I__3356 (
            .O(N__15644),
            .I(N__15641));
    LocalMux I__3355 (
            .O(N__15641),
            .I(\this_vram.mem_out_bus1_0 ));
    InMux I__3354 (
            .O(N__15638),
            .I(N__15635));
    LocalMux I__3353 (
            .O(N__15635),
            .I(\this_vram.mem_mem_1_0_RNISSKZ0Z11 ));
    InMux I__3352 (
            .O(N__15632),
            .I(N__15629));
    LocalMux I__3351 (
            .O(N__15629),
            .I(N__15625));
    InMux I__3350 (
            .O(N__15628),
            .I(N__15622));
    Span4Mux_v I__3349 (
            .O(N__15625),
            .I(N__15618));
    LocalMux I__3348 (
            .O(N__15622),
            .I(N__15615));
    InMux I__3347 (
            .O(N__15621),
            .I(N__15612));
    Span4Mux_h I__3346 (
            .O(N__15618),
            .I(N__15606));
    Span4Mux_v I__3345 (
            .O(N__15615),
            .I(N__15606));
    LocalMux I__3344 (
            .O(N__15612),
            .I(N__15603));
    InMux I__3343 (
            .O(N__15611),
            .I(N__15600));
    Odrv4 I__3342 (
            .O(N__15606),
            .I(\this_vram.mem_radregZ0Z_11 ));
    Odrv12 I__3341 (
            .O(N__15603),
            .I(\this_vram.mem_radregZ0Z_11 ));
    LocalMux I__3340 (
            .O(N__15600),
            .I(\this_vram.mem_radregZ0Z_11 ));
    CascadeMux I__3339 (
            .O(N__15593),
            .I(\this_vram.mem_N_109_cascade_ ));
    InMux I__3338 (
            .O(N__15590),
            .I(N__15585));
    InMux I__3337 (
            .O(N__15589),
            .I(N__15581));
    InMux I__3336 (
            .O(N__15588),
            .I(N__15578));
    LocalMux I__3335 (
            .O(N__15585),
            .I(N__15575));
    InMux I__3334 (
            .O(N__15584),
            .I(N__15572));
    LocalMux I__3333 (
            .O(N__15581),
            .I(N__15567));
    LocalMux I__3332 (
            .O(N__15578),
            .I(N__15567));
    Span4Mux_v I__3331 (
            .O(N__15575),
            .I(N__15558));
    LocalMux I__3330 (
            .O(N__15572),
            .I(N__15558));
    Span4Mux_v I__3329 (
            .O(N__15567),
            .I(N__15558));
    InMux I__3328 (
            .O(N__15566),
            .I(N__15555));
    InMux I__3327 (
            .O(N__15565),
            .I(N__15552));
    Span4Mux_v I__3326 (
            .O(N__15558),
            .I(N__15547));
    LocalMux I__3325 (
            .O(N__15555),
            .I(N__15547));
    LocalMux I__3324 (
            .O(N__15552),
            .I(N__15544));
    Span4Mux_v I__3323 (
            .O(N__15547),
            .I(N__15541));
    Span12Mux_v I__3322 (
            .O(N__15544),
            .I(N__15538));
    Sp12to4 I__3321 (
            .O(N__15541),
            .I(N__15535));
    Span12Mux_h I__3320 (
            .O(N__15538),
            .I(N__15532));
    Span12Mux_h I__3319 (
            .O(N__15535),
            .I(N__15529));
    Odrv12 I__3318 (
            .O(N__15532),
            .I(M_this_vram_read_data_0));
    Odrv12 I__3317 (
            .O(N__15529),
            .I(M_this_vram_read_data_0));
    InMux I__3316 (
            .O(N__15524),
            .I(N__15521));
    LocalMux I__3315 (
            .O(N__15521),
            .I(N__15518));
    Span4Mux_v I__3314 (
            .O(N__15518),
            .I(N__15515));
    Odrv4 I__3313 (
            .O(N__15515),
            .I(\this_vram.mem_out_bus0_0 ));
    InMux I__3312 (
            .O(N__15512),
            .I(N__15509));
    LocalMux I__3311 (
            .O(N__15509),
            .I(N__15506));
    Sp12to4 I__3310 (
            .O(N__15506),
            .I(N__15503));
    Span12Mux_v I__3309 (
            .O(N__15503),
            .I(N__15500));
    Odrv12 I__3308 (
            .O(N__15500),
            .I(\this_vram.mem_out_bus4_0 ));
    CascadeMux I__3307 (
            .O(N__15497),
            .I(\this_vram.mem_mem_0_0_RNIQOIZ0Z11_cascade_ ));
    InMux I__3306 (
            .O(N__15494),
            .I(N__15491));
    LocalMux I__3305 (
            .O(N__15491),
            .I(\this_vram.mem_N_112 ));
    CascadeMux I__3304 (
            .O(N__15488),
            .I(\this_vga_signals.g1_1_cascade_ ));
    InMux I__3303 (
            .O(N__15485),
            .I(N__15482));
    LocalMux I__3302 (
            .O(N__15482),
            .I(\this_vga_signals.N_15_0_0 ));
    InMux I__3301 (
            .O(N__15479),
            .I(N__15476));
    LocalMux I__3300 (
            .O(N__15476),
            .I(\this_vga_signals.N_353_0 ));
    CascadeMux I__3299 (
            .O(N__15473),
            .I(\this_vga_signals.N_3520_0_cascade_ ));
    InMux I__3298 (
            .O(N__15470),
            .I(N__15463));
    InMux I__3297 (
            .O(N__15469),
            .I(N__15460));
    InMux I__3296 (
            .O(N__15468),
            .I(N__15447));
    InMux I__3295 (
            .O(N__15467),
            .I(N__15447));
    InMux I__3294 (
            .O(N__15466),
            .I(N__15444));
    LocalMux I__3293 (
            .O(N__15463),
            .I(N__15439));
    LocalMux I__3292 (
            .O(N__15460),
            .I(N__15439));
    InMux I__3291 (
            .O(N__15459),
            .I(N__15434));
    InMux I__3290 (
            .O(N__15458),
            .I(N__15434));
    InMux I__3289 (
            .O(N__15457),
            .I(N__15429));
    InMux I__3288 (
            .O(N__15456),
            .I(N__15429));
    InMux I__3287 (
            .O(N__15455),
            .I(N__15424));
    InMux I__3286 (
            .O(N__15454),
            .I(N__15424));
    InMux I__3285 (
            .O(N__15453),
            .I(N__15419));
    InMux I__3284 (
            .O(N__15452),
            .I(N__15419));
    LocalMux I__3283 (
            .O(N__15447),
            .I(\this_vga_signals.CO1_2_1 ));
    LocalMux I__3282 (
            .O(N__15444),
            .I(\this_vga_signals.CO1_2_1 ));
    Odrv4 I__3281 (
            .O(N__15439),
            .I(\this_vga_signals.CO1_2_1 ));
    LocalMux I__3280 (
            .O(N__15434),
            .I(\this_vga_signals.CO1_2_1 ));
    LocalMux I__3279 (
            .O(N__15429),
            .I(\this_vga_signals.CO1_2_1 ));
    LocalMux I__3278 (
            .O(N__15424),
            .I(\this_vga_signals.CO1_2_1 ));
    LocalMux I__3277 (
            .O(N__15419),
            .I(\this_vga_signals.CO1_2_1 ));
    InMux I__3276 (
            .O(N__15404),
            .I(N__15401));
    LocalMux I__3275 (
            .O(N__15401),
            .I(\this_vga_signals.mult1_un40_sum_0_2 ));
    InMux I__3274 (
            .O(N__15398),
            .I(N__15392));
    InMux I__3273 (
            .O(N__15397),
            .I(N__15392));
    LocalMux I__3272 (
            .O(N__15392),
            .I(\this_vga_signals.g0_1_N_2L1 ));
    CascadeMux I__3271 (
            .O(N__15389),
            .I(N__15386));
    InMux I__3270 (
            .O(N__15386),
            .I(N__15383));
    LocalMux I__3269 (
            .O(N__15383),
            .I(N__15380));
    Span4Mux_h I__3268 (
            .O(N__15380),
            .I(N__15377));
    Span4Mux_h I__3267 (
            .O(N__15377),
            .I(N__15373));
    InMux I__3266 (
            .O(N__15376),
            .I(N__15370));
    Odrv4 I__3265 (
            .O(N__15373),
            .I(\this_vga_signals.N_1253_0 ));
    LocalMux I__3264 (
            .O(N__15370),
            .I(\this_vga_signals.N_1253_0 ));
    CascadeMux I__3263 (
            .O(N__15365),
            .I(\this_vga_signals.mult1_un40_sum_0_2_cascade_ ));
    InMux I__3262 (
            .O(N__15362),
            .I(N__15356));
    InMux I__3261 (
            .O(N__15361),
            .I(N__15356));
    LocalMux I__3260 (
            .O(N__15356),
            .I(\this_vga_signals.N_3_0 ));
    InMux I__3259 (
            .O(N__15353),
            .I(N__15340));
    InMux I__3258 (
            .O(N__15352),
            .I(N__15340));
    InMux I__3257 (
            .O(N__15351),
            .I(N__15335));
    InMux I__3256 (
            .O(N__15350),
            .I(N__15335));
    InMux I__3255 (
            .O(N__15349),
            .I(N__15330));
    InMux I__3254 (
            .O(N__15348),
            .I(N__15323));
    InMux I__3253 (
            .O(N__15347),
            .I(N__15323));
    InMux I__3252 (
            .O(N__15346),
            .I(N__15318));
    InMux I__3251 (
            .O(N__15345),
            .I(N__15315));
    LocalMux I__3250 (
            .O(N__15340),
            .I(N__15311));
    LocalMux I__3249 (
            .O(N__15335),
            .I(N__15308));
    InMux I__3248 (
            .O(N__15334),
            .I(N__15305));
    CascadeMux I__3247 (
            .O(N__15333),
            .I(N__15302));
    LocalMux I__3246 (
            .O(N__15330),
            .I(N__15294));
    InMux I__3245 (
            .O(N__15329),
            .I(N__15289));
    InMux I__3244 (
            .O(N__15328),
            .I(N__15289));
    LocalMux I__3243 (
            .O(N__15323),
            .I(N__15286));
    InMux I__3242 (
            .O(N__15322),
            .I(N__15283));
    InMux I__3241 (
            .O(N__15321),
            .I(N__15280));
    LocalMux I__3240 (
            .O(N__15318),
            .I(N__15275));
    LocalMux I__3239 (
            .O(N__15315),
            .I(N__15275));
    InMux I__3238 (
            .O(N__15314),
            .I(N__15272));
    Span4Mux_h I__3237 (
            .O(N__15311),
            .I(N__15269));
    Span4Mux_h I__3236 (
            .O(N__15308),
            .I(N__15264));
    LocalMux I__3235 (
            .O(N__15305),
            .I(N__15264));
    InMux I__3234 (
            .O(N__15302),
            .I(N__15255));
    InMux I__3233 (
            .O(N__15301),
            .I(N__15255));
    InMux I__3232 (
            .O(N__15300),
            .I(N__15255));
    InMux I__3231 (
            .O(N__15299),
            .I(N__15255));
    InMux I__3230 (
            .O(N__15298),
            .I(N__15250));
    InMux I__3229 (
            .O(N__15297),
            .I(N__15250));
    Span4Mux_v I__3228 (
            .O(N__15294),
            .I(N__15241));
    LocalMux I__3227 (
            .O(N__15289),
            .I(N__15241));
    Span4Mux_v I__3226 (
            .O(N__15286),
            .I(N__15241));
    LocalMux I__3225 (
            .O(N__15283),
            .I(N__15241));
    LocalMux I__3224 (
            .O(N__15280),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_0 ));
    Odrv4 I__3223 (
            .O(N__15275),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_0 ));
    LocalMux I__3222 (
            .O(N__15272),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_0 ));
    Odrv4 I__3221 (
            .O(N__15269),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_0 ));
    Odrv4 I__3220 (
            .O(N__15264),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_0 ));
    LocalMux I__3219 (
            .O(N__15255),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_0 ));
    LocalMux I__3218 (
            .O(N__15250),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_0 ));
    Odrv4 I__3217 (
            .O(N__15241),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_0 ));
    CascadeMux I__3216 (
            .O(N__15224),
            .I(\this_vga_signals.g0_1_N_5L7_x0_cascade_ ));
    InMux I__3215 (
            .O(N__15221),
            .I(N__15218));
    LocalMux I__3214 (
            .O(N__15218),
            .I(\this_vga_signals.g0_1_N_5L7_x1 ));
    InMux I__3213 (
            .O(N__15215),
            .I(N__15211));
    InMux I__3212 (
            .O(N__15214),
            .I(N__15208));
    LocalMux I__3211 (
            .O(N__15211),
            .I(N__15201));
    LocalMux I__3210 (
            .O(N__15208),
            .I(N__15197));
    InMux I__3209 (
            .O(N__15207),
            .I(N__15192));
    InMux I__3208 (
            .O(N__15206),
            .I(N__15192));
    InMux I__3207 (
            .O(N__15205),
            .I(N__15180));
    InMux I__3206 (
            .O(N__15204),
            .I(N__15180));
    Span4Mux_h I__3205 (
            .O(N__15201),
            .I(N__15176));
    InMux I__3204 (
            .O(N__15200),
            .I(N__15173));
    Span4Mux_h I__3203 (
            .O(N__15197),
            .I(N__15170));
    LocalMux I__3202 (
            .O(N__15192),
            .I(N__15167));
    InMux I__3201 (
            .O(N__15191),
            .I(N__15164));
    InMux I__3200 (
            .O(N__15190),
            .I(N__15159));
    InMux I__3199 (
            .O(N__15189),
            .I(N__15159));
    InMux I__3198 (
            .O(N__15188),
            .I(N__15150));
    InMux I__3197 (
            .O(N__15187),
            .I(N__15150));
    InMux I__3196 (
            .O(N__15186),
            .I(N__15150));
    InMux I__3195 (
            .O(N__15185),
            .I(N__15150));
    LocalMux I__3194 (
            .O(N__15180),
            .I(N__15147));
    InMux I__3193 (
            .O(N__15179),
            .I(N__15144));
    Odrv4 I__3192 (
            .O(N__15176),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    LocalMux I__3191 (
            .O(N__15173),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    Odrv4 I__3190 (
            .O(N__15170),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    Odrv4 I__3189 (
            .O(N__15167),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    LocalMux I__3188 (
            .O(N__15164),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    LocalMux I__3187 (
            .O(N__15159),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    LocalMux I__3186 (
            .O(N__15150),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    Odrv4 I__3185 (
            .O(N__15147),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    LocalMux I__3184 (
            .O(N__15144),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    CascadeMux I__3183 (
            .O(N__15125),
            .I(N__15114));
    InMux I__3182 (
            .O(N__15124),
            .I(N__15106));
    InMux I__3181 (
            .O(N__15123),
            .I(N__15106));
    CascadeMux I__3180 (
            .O(N__15122),
            .I(N__15102));
    CascadeMux I__3179 (
            .O(N__15121),
            .I(N__15097));
    CascadeMux I__3178 (
            .O(N__15120),
            .I(N__15094));
    CascadeMux I__3177 (
            .O(N__15119),
            .I(N__15086));
    CascadeMux I__3176 (
            .O(N__15118),
            .I(N__15079));
    InMux I__3175 (
            .O(N__15117),
            .I(N__15074));
    InMux I__3174 (
            .O(N__15114),
            .I(N__15074));
    CascadeMux I__3173 (
            .O(N__15113),
            .I(N__15071));
    InMux I__3172 (
            .O(N__15112),
            .I(N__15068));
    InMux I__3171 (
            .O(N__15111),
            .I(N__15065));
    LocalMux I__3170 (
            .O(N__15106),
            .I(N__15061));
    InMux I__3169 (
            .O(N__15105),
            .I(N__15058));
    InMux I__3168 (
            .O(N__15102),
            .I(N__15055));
    InMux I__3167 (
            .O(N__15101),
            .I(N__15050));
    InMux I__3166 (
            .O(N__15100),
            .I(N__15050));
    InMux I__3165 (
            .O(N__15097),
            .I(N__15047));
    InMux I__3164 (
            .O(N__15094),
            .I(N__15041));
    InMux I__3163 (
            .O(N__15093),
            .I(N__15038));
    InMux I__3162 (
            .O(N__15092),
            .I(N__15033));
    InMux I__3161 (
            .O(N__15091),
            .I(N__15033));
    InMux I__3160 (
            .O(N__15090),
            .I(N__15026));
    InMux I__3159 (
            .O(N__15089),
            .I(N__15026));
    InMux I__3158 (
            .O(N__15086),
            .I(N__15026));
    InMux I__3157 (
            .O(N__15085),
            .I(N__15019));
    InMux I__3156 (
            .O(N__15084),
            .I(N__15019));
    InMux I__3155 (
            .O(N__15083),
            .I(N__15019));
    InMux I__3154 (
            .O(N__15082),
            .I(N__15014));
    InMux I__3153 (
            .O(N__15079),
            .I(N__15014));
    LocalMux I__3152 (
            .O(N__15074),
            .I(N__15011));
    InMux I__3151 (
            .O(N__15071),
            .I(N__15008));
    LocalMux I__3150 (
            .O(N__15068),
            .I(N__15005));
    LocalMux I__3149 (
            .O(N__15065),
            .I(N__15002));
    InMux I__3148 (
            .O(N__15064),
            .I(N__14996));
    Span4Mux_v I__3147 (
            .O(N__15061),
            .I(N__14991));
    LocalMux I__3146 (
            .O(N__15058),
            .I(N__14991));
    LocalMux I__3145 (
            .O(N__15055),
            .I(N__14984));
    LocalMux I__3144 (
            .O(N__15050),
            .I(N__14984));
    LocalMux I__3143 (
            .O(N__15047),
            .I(N__14984));
    InMux I__3142 (
            .O(N__15046),
            .I(N__14977));
    InMux I__3141 (
            .O(N__15045),
            .I(N__14977));
    InMux I__3140 (
            .O(N__15044),
            .I(N__14977));
    LocalMux I__3139 (
            .O(N__15041),
            .I(N__14964));
    LocalMux I__3138 (
            .O(N__15038),
            .I(N__14964));
    LocalMux I__3137 (
            .O(N__15033),
            .I(N__14964));
    LocalMux I__3136 (
            .O(N__15026),
            .I(N__14964));
    LocalMux I__3135 (
            .O(N__15019),
            .I(N__14964));
    LocalMux I__3134 (
            .O(N__15014),
            .I(N__14964));
    Span4Mux_v I__3133 (
            .O(N__15011),
            .I(N__14961));
    LocalMux I__3132 (
            .O(N__15008),
            .I(N__14958));
    Span4Mux_v I__3131 (
            .O(N__15005),
            .I(N__14953));
    Span4Mux_v I__3130 (
            .O(N__15002),
            .I(N__14953));
    InMux I__3129 (
            .O(N__15001),
            .I(N__14950));
    InMux I__3128 (
            .O(N__15000),
            .I(N__14947));
    InMux I__3127 (
            .O(N__14999),
            .I(N__14944));
    LocalMux I__3126 (
            .O(N__14996),
            .I(N__14941));
    Span4Mux_h I__3125 (
            .O(N__14991),
            .I(N__14936));
    Span4Mux_v I__3124 (
            .O(N__14984),
            .I(N__14936));
    LocalMux I__3123 (
            .O(N__14977),
            .I(N__14931));
    Span4Mux_v I__3122 (
            .O(N__14964),
            .I(N__14931));
    Span4Mux_h I__3121 (
            .O(N__14961),
            .I(N__14920));
    Span4Mux_h I__3120 (
            .O(N__14958),
            .I(N__14920));
    Span4Mux_h I__3119 (
            .O(N__14953),
            .I(N__14920));
    LocalMux I__3118 (
            .O(N__14950),
            .I(N__14920));
    LocalMux I__3117 (
            .O(N__14947),
            .I(N__14920));
    LocalMux I__3116 (
            .O(N__14944),
            .I(\this_vga_signals.M_vaddress_qZ0Z_4 ));
    Odrv4 I__3115 (
            .O(N__14941),
            .I(\this_vga_signals.M_vaddress_qZ0Z_4 ));
    Odrv4 I__3114 (
            .O(N__14936),
            .I(\this_vga_signals.M_vaddress_qZ0Z_4 ));
    Odrv4 I__3113 (
            .O(N__14931),
            .I(\this_vga_signals.M_vaddress_qZ0Z_4 ));
    Odrv4 I__3112 (
            .O(N__14920),
            .I(\this_vga_signals.M_vaddress_qZ0Z_4 ));
    CascadeMux I__3111 (
            .O(N__14909),
            .I(\this_vga_signals.g0_1_N_5L7_ns_cascade_ ));
    InMux I__3110 (
            .O(N__14906),
            .I(N__14903));
    LocalMux I__3109 (
            .O(N__14903),
            .I(N__14900));
    Span4Mux_h I__3108 (
            .O(N__14900),
            .I(N__14897));
    Odrv4 I__3107 (
            .O(N__14897),
            .I(\this_vga_signals.g0_1_1_0 ));
    InMux I__3106 (
            .O(N__14894),
            .I(N__14890));
    InMux I__3105 (
            .O(N__14893),
            .I(N__14887));
    LocalMux I__3104 (
            .O(N__14890),
            .I(\this_vga_signals.N_355_0 ));
    LocalMux I__3103 (
            .O(N__14887),
            .I(\this_vga_signals.N_355_0 ));
    InMux I__3102 (
            .O(N__14882),
            .I(N__14879));
    LocalMux I__3101 (
            .O(N__14879),
            .I(\this_vga_signals.g1_4 ));
    InMux I__3100 (
            .O(N__14876),
            .I(N__14867));
    InMux I__3099 (
            .O(N__14875),
            .I(N__14862));
    InMux I__3098 (
            .O(N__14874),
            .I(N__14862));
    InMux I__3097 (
            .O(N__14873),
            .I(N__14857));
    InMux I__3096 (
            .O(N__14872),
            .I(N__14857));
    InMux I__3095 (
            .O(N__14871),
            .I(N__14854));
    InMux I__3094 (
            .O(N__14870),
            .I(N__14851));
    LocalMux I__3093 (
            .O(N__14867),
            .I(N__14846));
    LocalMux I__3092 (
            .O(N__14862),
            .I(N__14846));
    LocalMux I__3091 (
            .O(N__14857),
            .I(N__14843));
    LocalMux I__3090 (
            .O(N__14854),
            .I(N__14840));
    LocalMux I__3089 (
            .O(N__14851),
            .I(\this_vga_signals.M_vaddress_qZ0Z_7 ));
    Odrv4 I__3088 (
            .O(N__14846),
            .I(\this_vga_signals.M_vaddress_qZ0Z_7 ));
    Odrv4 I__3087 (
            .O(N__14843),
            .I(\this_vga_signals.M_vaddress_qZ0Z_7 ));
    Odrv12 I__3086 (
            .O(N__14840),
            .I(\this_vga_signals.M_vaddress_qZ0Z_7 ));
    InMux I__3085 (
            .O(N__14831),
            .I(N__14819));
    InMux I__3084 (
            .O(N__14830),
            .I(N__14816));
    InMux I__3083 (
            .O(N__14829),
            .I(N__14813));
    InMux I__3082 (
            .O(N__14828),
            .I(N__14810));
    InMux I__3081 (
            .O(N__14827),
            .I(N__14801));
    InMux I__3080 (
            .O(N__14826),
            .I(N__14801));
    InMux I__3079 (
            .O(N__14825),
            .I(N__14801));
    InMux I__3078 (
            .O(N__14824),
            .I(N__14801));
    InMux I__3077 (
            .O(N__14823),
            .I(N__14797));
    InMux I__3076 (
            .O(N__14822),
            .I(N__14794));
    LocalMux I__3075 (
            .O(N__14819),
            .I(N__14791));
    LocalMux I__3074 (
            .O(N__14816),
            .I(N__14782));
    LocalMux I__3073 (
            .O(N__14813),
            .I(N__14782));
    LocalMux I__3072 (
            .O(N__14810),
            .I(N__14782));
    LocalMux I__3071 (
            .O(N__14801),
            .I(N__14782));
    InMux I__3070 (
            .O(N__14800),
            .I(N__14779));
    LocalMux I__3069 (
            .O(N__14797),
            .I(\this_vga_signals.M_vaddress_qZ0Z_8 ));
    LocalMux I__3068 (
            .O(N__14794),
            .I(\this_vga_signals.M_vaddress_qZ0Z_8 ));
    Odrv4 I__3067 (
            .O(N__14791),
            .I(\this_vga_signals.M_vaddress_qZ0Z_8 ));
    Odrv4 I__3066 (
            .O(N__14782),
            .I(\this_vga_signals.M_vaddress_qZ0Z_8 ));
    LocalMux I__3065 (
            .O(N__14779),
            .I(\this_vga_signals.M_vaddress_qZ0Z_8 ));
    CascadeMux I__3064 (
            .O(N__14768),
            .I(N__14762));
    CascadeMux I__3063 (
            .O(N__14767),
            .I(N__14759));
    InMux I__3062 (
            .O(N__14766),
            .I(N__14750));
    InMux I__3061 (
            .O(N__14765),
            .I(N__14746));
    InMux I__3060 (
            .O(N__14762),
            .I(N__14743));
    InMux I__3059 (
            .O(N__14759),
            .I(N__14738));
    InMux I__3058 (
            .O(N__14758),
            .I(N__14738));
    InMux I__3057 (
            .O(N__14757),
            .I(N__14735));
    CascadeMux I__3056 (
            .O(N__14756),
            .I(N__14732));
    CascadeMux I__3055 (
            .O(N__14755),
            .I(N__14729));
    InMux I__3054 (
            .O(N__14754),
            .I(N__14724));
    InMux I__3053 (
            .O(N__14753),
            .I(N__14724));
    LocalMux I__3052 (
            .O(N__14750),
            .I(N__14720));
    InMux I__3051 (
            .O(N__14749),
            .I(N__14717));
    LocalMux I__3050 (
            .O(N__14746),
            .I(N__14708));
    LocalMux I__3049 (
            .O(N__14743),
            .I(N__14708));
    LocalMux I__3048 (
            .O(N__14738),
            .I(N__14708));
    LocalMux I__3047 (
            .O(N__14735),
            .I(N__14708));
    InMux I__3046 (
            .O(N__14732),
            .I(N__14702));
    InMux I__3045 (
            .O(N__14729),
            .I(N__14702));
    LocalMux I__3044 (
            .O(N__14724),
            .I(N__14699));
    InMux I__3043 (
            .O(N__14723),
            .I(N__14696));
    Span4Mux_v I__3042 (
            .O(N__14720),
            .I(N__14689));
    LocalMux I__3041 (
            .O(N__14717),
            .I(N__14689));
    Span4Mux_v I__3040 (
            .O(N__14708),
            .I(N__14689));
    InMux I__3039 (
            .O(N__14707),
            .I(N__14686));
    LocalMux I__3038 (
            .O(N__14702),
            .I(N__14683));
    Odrv4 I__3037 (
            .O(N__14699),
            .I(\this_vga_signals.M_vaddress_qZ0Z_6 ));
    LocalMux I__3036 (
            .O(N__14696),
            .I(\this_vga_signals.M_vaddress_qZ0Z_6 ));
    Odrv4 I__3035 (
            .O(N__14689),
            .I(\this_vga_signals.M_vaddress_qZ0Z_6 ));
    LocalMux I__3034 (
            .O(N__14686),
            .I(\this_vga_signals.M_vaddress_qZ0Z_6 ));
    Odrv4 I__3033 (
            .O(N__14683),
            .I(\this_vga_signals.M_vaddress_qZ0Z_6 ));
    InMux I__3032 (
            .O(N__14672),
            .I(N__14661));
    CascadeMux I__3031 (
            .O(N__14671),
            .I(N__14657));
    InMux I__3030 (
            .O(N__14670),
            .I(N__14653));
    InMux I__3029 (
            .O(N__14669),
            .I(N__14650));
    InMux I__3028 (
            .O(N__14668),
            .I(N__14645));
    InMux I__3027 (
            .O(N__14667),
            .I(N__14645));
    InMux I__3026 (
            .O(N__14666),
            .I(N__14640));
    InMux I__3025 (
            .O(N__14665),
            .I(N__14640));
    InMux I__3024 (
            .O(N__14664),
            .I(N__14637));
    LocalMux I__3023 (
            .O(N__14661),
            .I(N__14634));
    InMux I__3022 (
            .O(N__14660),
            .I(N__14629));
    InMux I__3021 (
            .O(N__14657),
            .I(N__14629));
    InMux I__3020 (
            .O(N__14656),
            .I(N__14626));
    LocalMux I__3019 (
            .O(N__14653),
            .I(\this_vga_signals.CO0 ));
    LocalMux I__3018 (
            .O(N__14650),
            .I(\this_vga_signals.CO0 ));
    LocalMux I__3017 (
            .O(N__14645),
            .I(\this_vga_signals.CO0 ));
    LocalMux I__3016 (
            .O(N__14640),
            .I(\this_vga_signals.CO0 ));
    LocalMux I__3015 (
            .O(N__14637),
            .I(\this_vga_signals.CO0 ));
    Odrv4 I__3014 (
            .O(N__14634),
            .I(\this_vga_signals.CO0 ));
    LocalMux I__3013 (
            .O(N__14629),
            .I(\this_vga_signals.CO0 ));
    LocalMux I__3012 (
            .O(N__14626),
            .I(\this_vga_signals.CO0 ));
    InMux I__3011 (
            .O(N__14609),
            .I(N__14606));
    LocalMux I__3010 (
            .O(N__14606),
            .I(N__14603));
    Span4Mux_h I__3009 (
            .O(N__14603),
            .I(N__14600));
    Odrv4 I__3008 (
            .O(N__14600),
            .I(\this_vga_signals.if_i2_mux ));
    InMux I__3007 (
            .O(N__14597),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_4 ));
    InMux I__3006 (
            .O(N__14594),
            .I(N__14587));
    InMux I__3005 (
            .O(N__14593),
            .I(N__14587));
    InMux I__3004 (
            .O(N__14592),
            .I(N__14584));
    LocalMux I__3003 (
            .O(N__14587),
            .I(N__14581));
    LocalMux I__3002 (
            .O(N__14584),
            .I(N__14578));
    Span4Mux_h I__3001 (
            .O(N__14581),
            .I(N__14575));
    Odrv4 I__3000 (
            .O(N__14578),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNEZ0 ));
    Odrv4 I__2999 (
            .O(N__14575),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNEZ0 ));
    InMux I__2998 (
            .O(N__14570),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_5 ));
    InMux I__2997 (
            .O(N__14567),
            .I(N__14558));
    InMux I__2996 (
            .O(N__14566),
            .I(N__14558));
    InMux I__2995 (
            .O(N__14565),
            .I(N__14558));
    LocalMux I__2994 (
            .O(N__14558),
            .I(N__14555));
    Odrv4 I__2993 (
            .O(N__14555),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOEZ0 ));
    InMux I__2992 (
            .O(N__14552),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_6 ));
    InMux I__2991 (
            .O(N__14549),
            .I(bfn_23_10_0_));
    InMux I__2990 (
            .O(N__14546),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_8 ));
    InMux I__2989 (
            .O(N__14543),
            .I(N__14540));
    LocalMux I__2988 (
            .O(N__14540),
            .I(N__14536));
    InMux I__2987 (
            .O(N__14539),
            .I(N__14533));
    Odrv4 I__2986 (
            .O(N__14536),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01REZ0 ));
    LocalMux I__2985 (
            .O(N__14533),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01REZ0 ));
    InMux I__2984 (
            .O(N__14528),
            .I(N__14524));
    InMux I__2983 (
            .O(N__14527),
            .I(N__14521));
    LocalMux I__2982 (
            .O(N__14524),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPEZ0 ));
    LocalMux I__2981 (
            .O(N__14521),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPEZ0 ));
    CascadeMux I__2980 (
            .O(N__14516),
            .I(N__14512));
    CascadeMux I__2979 (
            .O(N__14515),
            .I(N__14489));
    InMux I__2978 (
            .O(N__14512),
            .I(N__14486));
    CascadeMux I__2977 (
            .O(N__14511),
            .I(N__14483));
    CascadeMux I__2976 (
            .O(N__14510),
            .I(N__14478));
    CascadeMux I__2975 (
            .O(N__14509),
            .I(N__14472));
    CascadeMux I__2974 (
            .O(N__14508),
            .I(N__14468));
    InMux I__2973 (
            .O(N__14507),
            .I(N__14465));
    InMux I__2972 (
            .O(N__14506),
            .I(N__14462));
    InMux I__2971 (
            .O(N__14505),
            .I(N__14459));
    InMux I__2970 (
            .O(N__14504),
            .I(N__14454));
    InMux I__2969 (
            .O(N__14503),
            .I(N__14454));
    InMux I__2968 (
            .O(N__14502),
            .I(N__14449));
    InMux I__2967 (
            .O(N__14501),
            .I(N__14449));
    InMux I__2966 (
            .O(N__14500),
            .I(N__14445));
    InMux I__2965 (
            .O(N__14499),
            .I(N__14442));
    InMux I__2964 (
            .O(N__14498),
            .I(N__14437));
    InMux I__2963 (
            .O(N__14497),
            .I(N__14437));
    InMux I__2962 (
            .O(N__14496),
            .I(N__14427));
    InMux I__2961 (
            .O(N__14495),
            .I(N__14427));
    InMux I__2960 (
            .O(N__14494),
            .I(N__14427));
    InMux I__2959 (
            .O(N__14493),
            .I(N__14427));
    InMux I__2958 (
            .O(N__14492),
            .I(N__14422));
    InMux I__2957 (
            .O(N__14489),
            .I(N__14422));
    LocalMux I__2956 (
            .O(N__14486),
            .I(N__14419));
    InMux I__2955 (
            .O(N__14483),
            .I(N__14416));
    InMux I__2954 (
            .O(N__14482),
            .I(N__14413));
    InMux I__2953 (
            .O(N__14481),
            .I(N__14406));
    InMux I__2952 (
            .O(N__14478),
            .I(N__14406));
    InMux I__2951 (
            .O(N__14477),
            .I(N__14406));
    InMux I__2950 (
            .O(N__14476),
            .I(N__14403));
    InMux I__2949 (
            .O(N__14475),
            .I(N__14400));
    InMux I__2948 (
            .O(N__14472),
            .I(N__14397));
    InMux I__2947 (
            .O(N__14471),
            .I(N__14394));
    InMux I__2946 (
            .O(N__14468),
            .I(N__14391));
    LocalMux I__2945 (
            .O(N__14465),
            .I(N__14388));
    LocalMux I__2944 (
            .O(N__14462),
            .I(N__14385));
    LocalMux I__2943 (
            .O(N__14459),
            .I(N__14382));
    LocalMux I__2942 (
            .O(N__14454),
            .I(N__14377));
    LocalMux I__2941 (
            .O(N__14449),
            .I(N__14377));
    InMux I__2940 (
            .O(N__14448),
            .I(N__14374));
    LocalMux I__2939 (
            .O(N__14445),
            .I(N__14367));
    LocalMux I__2938 (
            .O(N__14442),
            .I(N__14367));
    LocalMux I__2937 (
            .O(N__14437),
            .I(N__14367));
    CascadeMux I__2936 (
            .O(N__14436),
            .I(N__14364));
    LocalMux I__2935 (
            .O(N__14427),
            .I(N__14351));
    LocalMux I__2934 (
            .O(N__14422),
            .I(N__14351));
    Span4Mux_h I__2933 (
            .O(N__14419),
            .I(N__14351));
    LocalMux I__2932 (
            .O(N__14416),
            .I(N__14351));
    LocalMux I__2931 (
            .O(N__14413),
            .I(N__14351));
    LocalMux I__2930 (
            .O(N__14406),
            .I(N__14351));
    LocalMux I__2929 (
            .O(N__14403),
            .I(N__14340));
    LocalMux I__2928 (
            .O(N__14400),
            .I(N__14340));
    LocalMux I__2927 (
            .O(N__14397),
            .I(N__14340));
    LocalMux I__2926 (
            .O(N__14394),
            .I(N__14340));
    LocalMux I__2925 (
            .O(N__14391),
            .I(N__14340));
    Span4Mux_v I__2924 (
            .O(N__14388),
            .I(N__14336));
    Span4Mux_v I__2923 (
            .O(N__14385),
            .I(N__14329));
    Span4Mux_v I__2922 (
            .O(N__14382),
            .I(N__14329));
    Span4Mux_h I__2921 (
            .O(N__14377),
            .I(N__14329));
    LocalMux I__2920 (
            .O(N__14374),
            .I(N__14324));
    Span4Mux_v I__2919 (
            .O(N__14367),
            .I(N__14324));
    InMux I__2918 (
            .O(N__14364),
            .I(N__14321));
    Span4Mux_v I__2917 (
            .O(N__14351),
            .I(N__14316));
    Span4Mux_v I__2916 (
            .O(N__14340),
            .I(N__14316));
    InMux I__2915 (
            .O(N__14339),
            .I(N__14313));
    Span4Mux_h I__2914 (
            .O(N__14336),
            .I(N__14310));
    Span4Mux_h I__2913 (
            .O(N__14329),
            .I(N__14307));
    Span4Mux_h I__2912 (
            .O(N__14324),
            .I(N__14302));
    LocalMux I__2911 (
            .O(N__14321),
            .I(N__14302));
    Span4Mux_h I__2910 (
            .O(N__14316),
            .I(N__14299));
    LocalMux I__2909 (
            .O(N__14313),
            .I(\this_vga_signals.M_vaddress_qZ0Z_3 ));
    Odrv4 I__2908 (
            .O(N__14310),
            .I(\this_vga_signals.M_vaddress_qZ0Z_3 ));
    Odrv4 I__2907 (
            .O(N__14307),
            .I(\this_vga_signals.M_vaddress_qZ0Z_3 ));
    Odrv4 I__2906 (
            .O(N__14302),
            .I(\this_vga_signals.M_vaddress_qZ0Z_3 ));
    Odrv4 I__2905 (
            .O(N__14299),
            .I(\this_vga_signals.M_vaddress_qZ0Z_3 ));
    CascadeMux I__2904 (
            .O(N__14288),
            .I(\this_vga_signals.N_1253_0_cascade_ ));
    CEMux I__2903 (
            .O(N__14285),
            .I(N__14282));
    LocalMux I__2902 (
            .O(N__14282),
            .I(N__14278));
    CEMux I__2901 (
            .O(N__14281),
            .I(N__14275));
    Span4Mux_v I__2900 (
            .O(N__14278),
            .I(N__14270));
    LocalMux I__2899 (
            .O(N__14275),
            .I(N__14270));
    Span4Mux_v I__2898 (
            .O(N__14270),
            .I(N__14267));
    Span4Mux_v I__2897 (
            .O(N__14267),
            .I(N__14264));
    Odrv4 I__2896 (
            .O(N__14264),
            .I(\this_vram.mem_WE_2 ));
    InMux I__2895 (
            .O(N__14261),
            .I(N__14258));
    LocalMux I__2894 (
            .O(N__14258),
            .I(N__14255));
    Span12Mux_h I__2893 (
            .O(N__14255),
            .I(N__14252));
    Odrv12 I__2892 (
            .O(N__14252),
            .I(port_address_c_5));
    InMux I__2891 (
            .O(N__14249),
            .I(N__14246));
    LocalMux I__2890 (
            .O(N__14246),
            .I(N__14243));
    Span12Mux_v I__2889 (
            .O(N__14243),
            .I(N__14240));
    Odrv12 I__2888 (
            .O(N__14240),
            .I(port_address_c_2));
    InMux I__2887 (
            .O(N__14237),
            .I(N__14234));
    LocalMux I__2886 (
            .O(N__14234),
            .I(N__14231));
    Span4Mux_v I__2885 (
            .O(N__14231),
            .I(N__14228));
    Sp12to4 I__2884 (
            .O(N__14228),
            .I(N__14225));
    Odrv12 I__2883 (
            .O(N__14225),
            .I(port_address_c_6));
    InMux I__2882 (
            .O(N__14222),
            .I(N__14219));
    LocalMux I__2881 (
            .O(N__14219),
            .I(N__14216));
    Span4Mux_v I__2880 (
            .O(N__14216),
            .I(N__14213));
    Odrv4 I__2879 (
            .O(N__14213),
            .I(\this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3Z0Z_0 ));
    InMux I__2878 (
            .O(N__14210),
            .I(N__14207));
    LocalMux I__2877 (
            .O(N__14207),
            .I(N__14203));
    InMux I__2876 (
            .O(N__14206),
            .I(N__14200));
    Span4Mux_h I__2875 (
            .O(N__14203),
            .I(N__14196));
    LocalMux I__2874 (
            .O(N__14200),
            .I(N__14193));
    InMux I__2873 (
            .O(N__14199),
            .I(N__14190));
    Span4Mux_v I__2872 (
            .O(N__14196),
            .I(N__14184));
    Span4Mux_h I__2871 (
            .O(N__14193),
            .I(N__14184));
    LocalMux I__2870 (
            .O(N__14190),
            .I(N__14181));
    InMux I__2869 (
            .O(N__14189),
            .I(N__14178));
    Span4Mux_v I__2868 (
            .O(N__14184),
            .I(N__14172));
    Span4Mux_h I__2867 (
            .O(N__14181),
            .I(N__14172));
    LocalMux I__2866 (
            .O(N__14178),
            .I(N__14169));
    InMux I__2865 (
            .O(N__14177),
            .I(N__14166));
    Span4Mux_v I__2864 (
            .O(N__14172),
            .I(N__14160));
    Span4Mux_h I__2863 (
            .O(N__14169),
            .I(N__14160));
    LocalMux I__2862 (
            .O(N__14166),
            .I(N__14157));
    InMux I__2861 (
            .O(N__14165),
            .I(N__14154));
    Span4Mux_v I__2860 (
            .O(N__14160),
            .I(N__14147));
    Span4Mux_h I__2859 (
            .O(N__14157),
            .I(N__14147));
    LocalMux I__2858 (
            .O(N__14154),
            .I(N__14144));
    InMux I__2857 (
            .O(N__14153),
            .I(N__14141));
    InMux I__2856 (
            .O(N__14152),
            .I(N__14138));
    Span4Mux_v I__2855 (
            .O(N__14147),
            .I(N__14133));
    Span4Mux_h I__2854 (
            .O(N__14144),
            .I(N__14133));
    LocalMux I__2853 (
            .O(N__14141),
            .I(N__14130));
    LocalMux I__2852 (
            .O(N__14138),
            .I(N__14127));
    Span4Mux_v I__2851 (
            .O(N__14133),
            .I(N__14119));
    Span4Mux_h I__2850 (
            .O(N__14130),
            .I(N__14119));
    Span4Mux_h I__2849 (
            .O(N__14127),
            .I(N__14119));
    InMux I__2848 (
            .O(N__14126),
            .I(N__14116));
    Odrv4 I__2847 (
            .O(N__14119),
            .I(M_current_data_qZ0Z_1));
    LocalMux I__2846 (
            .O(N__14116),
            .I(M_current_data_qZ0Z_1));
    CascadeMux I__2845 (
            .O(N__14111),
            .I(N__14107));
    InMux I__2844 (
            .O(N__14110),
            .I(N__14104));
    InMux I__2843 (
            .O(N__14107),
            .I(N__14101));
    LocalMux I__2842 (
            .O(N__14104),
            .I(N__14094));
    LocalMux I__2841 (
            .O(N__14101),
            .I(N__14094));
    InMux I__2840 (
            .O(N__14100),
            .I(N__14089));
    InMux I__2839 (
            .O(N__14099),
            .I(N__14086));
    Span4Mux_h I__2838 (
            .O(N__14094),
            .I(N__14083));
    InMux I__2837 (
            .O(N__14093),
            .I(N__14077));
    InMux I__2836 (
            .O(N__14092),
            .I(N__14077));
    LocalMux I__2835 (
            .O(N__14089),
            .I(N__14072));
    LocalMux I__2834 (
            .O(N__14086),
            .I(N__14072));
    Span4Mux_v I__2833 (
            .O(N__14083),
            .I(N__14069));
    InMux I__2832 (
            .O(N__14082),
            .I(N__14066));
    LocalMux I__2831 (
            .O(N__14077),
            .I(N__14063));
    Span4Mux_h I__2830 (
            .O(N__14072),
            .I(N__14058));
    Span4Mux_h I__2829 (
            .O(N__14069),
            .I(N__14058));
    LocalMux I__2828 (
            .O(N__14066),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    Odrv4 I__2827 (
            .O(N__14063),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    Odrv4 I__2826 (
            .O(N__14058),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    InMux I__2825 (
            .O(N__14051),
            .I(N__14047));
    InMux I__2824 (
            .O(N__14050),
            .I(N__14044));
    LocalMux I__2823 (
            .O(N__14047),
            .I(N__14041));
    LocalMux I__2822 (
            .O(N__14044),
            .I(\this_vga_signals.M_vaddress_qZ0Z_0 ));
    Odrv4 I__2821 (
            .O(N__14041),
            .I(\this_vga_signals.M_vaddress_qZ0Z_0 ));
    InMux I__2820 (
            .O(N__14036),
            .I(N__14033));
    LocalMux I__2819 (
            .O(N__14033),
            .I(N__14024));
    InMux I__2818 (
            .O(N__14032),
            .I(N__14021));
    InMux I__2817 (
            .O(N__14031),
            .I(N__14017));
    InMux I__2816 (
            .O(N__14030),
            .I(N__14010));
    InMux I__2815 (
            .O(N__14029),
            .I(N__14010));
    InMux I__2814 (
            .O(N__14028),
            .I(N__14010));
    InMux I__2813 (
            .O(N__14027),
            .I(N__14007));
    Span4Mux_v I__2812 (
            .O(N__14024),
            .I(N__14004));
    LocalMux I__2811 (
            .O(N__14021),
            .I(N__14001));
    InMux I__2810 (
            .O(N__14020),
            .I(N__13998));
    LocalMux I__2809 (
            .O(N__14017),
            .I(N__13991));
    LocalMux I__2808 (
            .O(N__14010),
            .I(N__13991));
    LocalMux I__2807 (
            .O(N__14007),
            .I(N__13991));
    Span4Mux_h I__2806 (
            .O(N__14004),
            .I(N__13986));
    Span4Mux_h I__2805 (
            .O(N__14001),
            .I(N__13986));
    LocalMux I__2804 (
            .O(N__13998),
            .I(\this_vga_signals.M_vaddress_qZ0Z_1 ));
    Odrv12 I__2803 (
            .O(N__13991),
            .I(\this_vga_signals.M_vaddress_qZ0Z_1 ));
    Odrv4 I__2802 (
            .O(N__13986),
            .I(\this_vga_signals.M_vaddress_qZ0Z_1 ));
    InMux I__2801 (
            .O(N__13979),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_0 ));
    CascadeMux I__2800 (
            .O(N__13976),
            .I(N__13969));
    InMux I__2799 (
            .O(N__13975),
            .I(N__13966));
    CascadeMux I__2798 (
            .O(N__13974),
            .I(N__13955));
    CascadeMux I__2797 (
            .O(N__13973),
            .I(N__13952));
    CascadeMux I__2796 (
            .O(N__13972),
            .I(N__13949));
    InMux I__2795 (
            .O(N__13969),
            .I(N__13945));
    LocalMux I__2794 (
            .O(N__13966),
            .I(N__13941));
    InMux I__2793 (
            .O(N__13965),
            .I(N__13936));
    InMux I__2792 (
            .O(N__13964),
            .I(N__13936));
    InMux I__2791 (
            .O(N__13963),
            .I(N__13933));
    InMux I__2790 (
            .O(N__13962),
            .I(N__13929));
    InMux I__2789 (
            .O(N__13961),
            .I(N__13926));
    InMux I__2788 (
            .O(N__13960),
            .I(N__13915));
    InMux I__2787 (
            .O(N__13959),
            .I(N__13915));
    InMux I__2786 (
            .O(N__13958),
            .I(N__13915));
    InMux I__2785 (
            .O(N__13955),
            .I(N__13915));
    InMux I__2784 (
            .O(N__13952),
            .I(N__13915));
    InMux I__2783 (
            .O(N__13949),
            .I(N__13910));
    InMux I__2782 (
            .O(N__13948),
            .I(N__13910));
    LocalMux I__2781 (
            .O(N__13945),
            .I(N__13907));
    InMux I__2780 (
            .O(N__13944),
            .I(N__13904));
    Span4Mux_v I__2779 (
            .O(N__13941),
            .I(N__13901));
    LocalMux I__2778 (
            .O(N__13936),
            .I(N__13896));
    LocalMux I__2777 (
            .O(N__13933),
            .I(N__13896));
    InMux I__2776 (
            .O(N__13932),
            .I(N__13891));
    LocalMux I__2775 (
            .O(N__13929),
            .I(N__13882));
    LocalMux I__2774 (
            .O(N__13926),
            .I(N__13882));
    LocalMux I__2773 (
            .O(N__13915),
            .I(N__13882));
    LocalMux I__2772 (
            .O(N__13910),
            .I(N__13882));
    Span12Mux_h I__2771 (
            .O(N__13907),
            .I(N__13879));
    LocalMux I__2770 (
            .O(N__13904),
            .I(N__13871));
    Span4Mux_h I__2769 (
            .O(N__13901),
            .I(N__13871));
    Span4Mux_v I__2768 (
            .O(N__13896),
            .I(N__13871));
    InMux I__2767 (
            .O(N__13895),
            .I(N__13866));
    InMux I__2766 (
            .O(N__13894),
            .I(N__13866));
    LocalMux I__2765 (
            .O(N__13891),
            .I(N__13861));
    Span4Mux_v I__2764 (
            .O(N__13882),
            .I(N__13861));
    Span12Mux_v I__2763 (
            .O(N__13879),
            .I(N__13858));
    InMux I__2762 (
            .O(N__13878),
            .I(N__13855));
    Sp12to4 I__2761 (
            .O(N__13871),
            .I(N__13850));
    LocalMux I__2760 (
            .O(N__13866),
            .I(N__13850));
    Span4Mux_h I__2759 (
            .O(N__13861),
            .I(N__13847));
    Odrv12 I__2758 (
            .O(N__13858),
            .I(\this_vga_signals.M_vaddress_qZ0Z_2 ));
    LocalMux I__2757 (
            .O(N__13855),
            .I(\this_vga_signals.M_vaddress_qZ0Z_2 ));
    Odrv12 I__2756 (
            .O(N__13850),
            .I(\this_vga_signals.M_vaddress_qZ0Z_2 ));
    Odrv4 I__2755 (
            .O(N__13847),
            .I(\this_vga_signals.M_vaddress_qZ0Z_2 ));
    InMux I__2754 (
            .O(N__13838),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_1 ));
    InMux I__2753 (
            .O(N__13835),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_2 ));
    InMux I__2752 (
            .O(N__13832),
            .I(\this_vga_signals.un1_M_vaddress_q_cry_3 ));
    CascadeMux I__2751 (
            .O(N__13829),
            .I(N__13825));
    InMux I__2750 (
            .O(N__13828),
            .I(N__13820));
    InMux I__2749 (
            .O(N__13825),
            .I(N__13820));
    LocalMux I__2748 (
            .O(N__13820),
            .I(\this_vga_signals.N_9_0 ));
    CascadeMux I__2747 (
            .O(N__13817),
            .I(N__13812));
    InMux I__2746 (
            .O(N__13816),
            .I(N__13806));
    CascadeMux I__2745 (
            .O(N__13815),
            .I(N__13801));
    InMux I__2744 (
            .O(N__13812),
            .I(N__13798));
    InMux I__2743 (
            .O(N__13811),
            .I(N__13795));
    InMux I__2742 (
            .O(N__13810),
            .I(N__13792));
    InMux I__2741 (
            .O(N__13809),
            .I(N__13789));
    LocalMux I__2740 (
            .O(N__13806),
            .I(N__13786));
    InMux I__2739 (
            .O(N__13805),
            .I(N__13783));
    InMux I__2738 (
            .O(N__13804),
            .I(N__13778));
    InMux I__2737 (
            .O(N__13801),
            .I(N__13778));
    LocalMux I__2736 (
            .O(N__13798),
            .I(\this_vga_signals.M_vaddress_q_6_repZ0Z1 ));
    LocalMux I__2735 (
            .O(N__13795),
            .I(\this_vga_signals.M_vaddress_q_6_repZ0Z1 ));
    LocalMux I__2734 (
            .O(N__13792),
            .I(\this_vga_signals.M_vaddress_q_6_repZ0Z1 ));
    LocalMux I__2733 (
            .O(N__13789),
            .I(\this_vga_signals.M_vaddress_q_6_repZ0Z1 ));
    Odrv4 I__2732 (
            .O(N__13786),
            .I(\this_vga_signals.M_vaddress_q_6_repZ0Z1 ));
    LocalMux I__2731 (
            .O(N__13783),
            .I(\this_vga_signals.M_vaddress_q_6_repZ0Z1 ));
    LocalMux I__2730 (
            .O(N__13778),
            .I(\this_vga_signals.M_vaddress_q_6_repZ0Z1 ));
    CascadeMux I__2729 (
            .O(N__13763),
            .I(N__13756));
    CascadeMux I__2728 (
            .O(N__13762),
            .I(N__13753));
    CascadeMux I__2727 (
            .O(N__13761),
            .I(N__13749));
    InMux I__2726 (
            .O(N__13760),
            .I(N__13744));
    InMux I__2725 (
            .O(N__13759),
            .I(N__13741));
    InMux I__2724 (
            .O(N__13756),
            .I(N__13734));
    InMux I__2723 (
            .O(N__13753),
            .I(N__13734));
    InMux I__2722 (
            .O(N__13752),
            .I(N__13734));
    InMux I__2721 (
            .O(N__13749),
            .I(N__13731));
    InMux I__2720 (
            .O(N__13748),
            .I(N__13728));
    InMux I__2719 (
            .O(N__13747),
            .I(N__13725));
    LocalMux I__2718 (
            .O(N__13744),
            .I(N__13720));
    LocalMux I__2717 (
            .O(N__13741),
            .I(N__13720));
    LocalMux I__2716 (
            .O(N__13734),
            .I(N__13717));
    LocalMux I__2715 (
            .O(N__13731),
            .I(\this_vga_signals.M_vaddress_q_7_repZ0Z1 ));
    LocalMux I__2714 (
            .O(N__13728),
            .I(\this_vga_signals.M_vaddress_q_7_repZ0Z1 ));
    LocalMux I__2713 (
            .O(N__13725),
            .I(\this_vga_signals.M_vaddress_q_7_repZ0Z1 ));
    Odrv12 I__2712 (
            .O(N__13720),
            .I(\this_vga_signals.M_vaddress_q_7_repZ0Z1 ));
    Odrv4 I__2711 (
            .O(N__13717),
            .I(\this_vga_signals.M_vaddress_q_7_repZ0Z1 ));
    InMux I__2710 (
            .O(N__13706),
            .I(N__13696));
    InMux I__2709 (
            .O(N__13705),
            .I(N__13696));
    InMux I__2708 (
            .O(N__13704),
            .I(N__13696));
    InMux I__2707 (
            .O(N__13703),
            .I(N__13693));
    LocalMux I__2706 (
            .O(N__13696),
            .I(N__13688));
    LocalMux I__2705 (
            .O(N__13693),
            .I(N__13688));
    Odrv4 I__2704 (
            .O(N__13688),
            .I(\this_vga_signals.N_15_0 ));
    CascadeMux I__2703 (
            .O(N__13685),
            .I(\this_vga_signals.N_15_0_0_cascade_ ));
    InMux I__2702 (
            .O(N__13682),
            .I(N__13679));
    LocalMux I__2701 (
            .O(N__13679),
            .I(N__13674));
    InMux I__2700 (
            .O(N__13678),
            .I(N__13670));
    InMux I__2699 (
            .O(N__13677),
            .I(N__13666));
    Span4Mux_h I__2698 (
            .O(N__13674),
            .I(N__13663));
    InMux I__2697 (
            .O(N__13673),
            .I(N__13660));
    LocalMux I__2696 (
            .O(N__13670),
            .I(N__13648));
    InMux I__2695 (
            .O(N__13669),
            .I(N__13645));
    LocalMux I__2694 (
            .O(N__13666),
            .I(N__13640));
    Span4Mux_v I__2693 (
            .O(N__13663),
            .I(N__13640));
    LocalMux I__2692 (
            .O(N__13660),
            .I(N__13637));
    InMux I__2691 (
            .O(N__13659),
            .I(N__13628));
    InMux I__2690 (
            .O(N__13658),
            .I(N__13628));
    InMux I__2689 (
            .O(N__13657),
            .I(N__13628));
    InMux I__2688 (
            .O(N__13656),
            .I(N__13628));
    InMux I__2687 (
            .O(N__13655),
            .I(N__13617));
    InMux I__2686 (
            .O(N__13654),
            .I(N__13617));
    InMux I__2685 (
            .O(N__13653),
            .I(N__13617));
    InMux I__2684 (
            .O(N__13652),
            .I(N__13617));
    InMux I__2683 (
            .O(N__13651),
            .I(N__13617));
    Odrv12 I__2682 (
            .O(N__13648),
            .I(\this_vga_signals.M_haddress_qZ0Z_9 ));
    LocalMux I__2681 (
            .O(N__13645),
            .I(\this_vga_signals.M_haddress_qZ0Z_9 ));
    Odrv4 I__2680 (
            .O(N__13640),
            .I(\this_vga_signals.M_haddress_qZ0Z_9 ));
    Odrv4 I__2679 (
            .O(N__13637),
            .I(\this_vga_signals.M_haddress_qZ0Z_9 ));
    LocalMux I__2678 (
            .O(N__13628),
            .I(\this_vga_signals.M_haddress_qZ0Z_9 ));
    LocalMux I__2677 (
            .O(N__13617),
            .I(\this_vga_signals.M_haddress_qZ0Z_9 ));
    InMux I__2676 (
            .O(N__13604),
            .I(N__13601));
    LocalMux I__2675 (
            .O(N__13601),
            .I(N__13596));
    InMux I__2674 (
            .O(N__13600),
            .I(N__13592));
    InMux I__2673 (
            .O(N__13599),
            .I(N__13588));
    Span4Mux_h I__2672 (
            .O(N__13596),
            .I(N__13585));
    InMux I__2671 (
            .O(N__13595),
            .I(N__13582));
    LocalMux I__2670 (
            .O(N__13592),
            .I(N__13570));
    InMux I__2669 (
            .O(N__13591),
            .I(N__13567));
    LocalMux I__2668 (
            .O(N__13588),
            .I(N__13562));
    Span4Mux_v I__2667 (
            .O(N__13585),
            .I(N__13562));
    LocalMux I__2666 (
            .O(N__13582),
            .I(N__13559));
    InMux I__2665 (
            .O(N__13581),
            .I(N__13552));
    InMux I__2664 (
            .O(N__13580),
            .I(N__13552));
    InMux I__2663 (
            .O(N__13579),
            .I(N__13552));
    InMux I__2662 (
            .O(N__13578),
            .I(N__13547));
    InMux I__2661 (
            .O(N__13577),
            .I(N__13547));
    InMux I__2660 (
            .O(N__13576),
            .I(N__13542));
    InMux I__2659 (
            .O(N__13575),
            .I(N__13542));
    InMux I__2658 (
            .O(N__13574),
            .I(N__13537));
    InMux I__2657 (
            .O(N__13573),
            .I(N__13537));
    Odrv12 I__2656 (
            .O(N__13570),
            .I(\this_vga_signals.M_haddress_qZ0Z_8 ));
    LocalMux I__2655 (
            .O(N__13567),
            .I(\this_vga_signals.M_haddress_qZ0Z_8 ));
    Odrv4 I__2654 (
            .O(N__13562),
            .I(\this_vga_signals.M_haddress_qZ0Z_8 ));
    Odrv4 I__2653 (
            .O(N__13559),
            .I(\this_vga_signals.M_haddress_qZ0Z_8 ));
    LocalMux I__2652 (
            .O(N__13552),
            .I(\this_vga_signals.M_haddress_qZ0Z_8 ));
    LocalMux I__2651 (
            .O(N__13547),
            .I(\this_vga_signals.M_haddress_qZ0Z_8 ));
    LocalMux I__2650 (
            .O(N__13542),
            .I(\this_vga_signals.M_haddress_qZ0Z_8 ));
    LocalMux I__2649 (
            .O(N__13537),
            .I(\this_vga_signals.M_haddress_qZ0Z_8 ));
    CascadeMux I__2648 (
            .O(N__13520),
            .I(N__13517));
    InMux I__2647 (
            .O(N__13517),
            .I(N__13511));
    CascadeMux I__2646 (
            .O(N__13516),
            .I(N__13508));
    CascadeMux I__2645 (
            .O(N__13515),
            .I(N__13504));
    CascadeMux I__2644 (
            .O(N__13514),
            .I(N__13498));
    LocalMux I__2643 (
            .O(N__13511),
            .I(N__13494));
    InMux I__2642 (
            .O(N__13508),
            .I(N__13490));
    CascadeMux I__2641 (
            .O(N__13507),
            .I(N__13487));
    InMux I__2640 (
            .O(N__13504),
            .I(N__13484));
    CascadeMux I__2639 (
            .O(N__13503),
            .I(N__13480));
    CascadeMux I__2638 (
            .O(N__13502),
            .I(N__13477));
    CascadeMux I__2637 (
            .O(N__13501),
            .I(N__13472));
    InMux I__2636 (
            .O(N__13498),
            .I(N__13465));
    InMux I__2635 (
            .O(N__13497),
            .I(N__13465));
    Span4Mux_h I__2634 (
            .O(N__13494),
            .I(N__13462));
    InMux I__2633 (
            .O(N__13493),
            .I(N__13459));
    LocalMux I__2632 (
            .O(N__13490),
            .I(N__13456));
    InMux I__2631 (
            .O(N__13487),
            .I(N__13453));
    LocalMux I__2630 (
            .O(N__13484),
            .I(N__13450));
    InMux I__2629 (
            .O(N__13483),
            .I(N__13445));
    InMux I__2628 (
            .O(N__13480),
            .I(N__13445));
    InMux I__2627 (
            .O(N__13477),
            .I(N__13436));
    InMux I__2626 (
            .O(N__13476),
            .I(N__13436));
    InMux I__2625 (
            .O(N__13475),
            .I(N__13436));
    InMux I__2624 (
            .O(N__13472),
            .I(N__13436));
    InMux I__2623 (
            .O(N__13471),
            .I(N__13431));
    InMux I__2622 (
            .O(N__13470),
            .I(N__13431));
    LocalMux I__2621 (
            .O(N__13465),
            .I(N__13426));
    Span4Mux_v I__2620 (
            .O(N__13462),
            .I(N__13426));
    LocalMux I__2619 (
            .O(N__13459),
            .I(\this_vga_signals.M_haddress_qZ0Z_10 ));
    Odrv12 I__2618 (
            .O(N__13456),
            .I(\this_vga_signals.M_haddress_qZ0Z_10 ));
    LocalMux I__2617 (
            .O(N__13453),
            .I(\this_vga_signals.M_haddress_qZ0Z_10 ));
    Odrv4 I__2616 (
            .O(N__13450),
            .I(\this_vga_signals.M_haddress_qZ0Z_10 ));
    LocalMux I__2615 (
            .O(N__13445),
            .I(\this_vga_signals.M_haddress_qZ0Z_10 ));
    LocalMux I__2614 (
            .O(N__13436),
            .I(\this_vga_signals.M_haddress_qZ0Z_10 ));
    LocalMux I__2613 (
            .O(N__13431),
            .I(\this_vga_signals.M_haddress_qZ0Z_10 ));
    Odrv4 I__2612 (
            .O(N__13426),
            .I(\this_vga_signals.M_haddress_qZ0Z_10 ));
    InMux I__2611 (
            .O(N__13409),
            .I(N__13406));
    LocalMux I__2610 (
            .O(N__13406),
            .I(N__13399));
    InMux I__2609 (
            .O(N__13405),
            .I(N__13395));
    InMux I__2608 (
            .O(N__13404),
            .I(N__13392));
    InMux I__2607 (
            .O(N__13403),
            .I(N__13387));
    InMux I__2606 (
            .O(N__13402),
            .I(N__13387));
    Span4Mux_v I__2605 (
            .O(N__13399),
            .I(N__13376));
    InMux I__2604 (
            .O(N__13398),
            .I(N__13373));
    LocalMux I__2603 (
            .O(N__13395),
            .I(N__13370));
    LocalMux I__2602 (
            .O(N__13392),
            .I(N__13365));
    LocalMux I__2601 (
            .O(N__13387),
            .I(N__13365));
    InMux I__2600 (
            .O(N__13386),
            .I(N__13354));
    InMux I__2599 (
            .O(N__13385),
            .I(N__13354));
    InMux I__2598 (
            .O(N__13384),
            .I(N__13354));
    InMux I__2597 (
            .O(N__13383),
            .I(N__13354));
    InMux I__2596 (
            .O(N__13382),
            .I(N__13354));
    InMux I__2595 (
            .O(N__13381),
            .I(N__13347));
    InMux I__2594 (
            .O(N__13380),
            .I(N__13347));
    InMux I__2593 (
            .O(N__13379),
            .I(N__13347));
    Span4Mux_h I__2592 (
            .O(N__13376),
            .I(N__13344));
    LocalMux I__2591 (
            .O(N__13373),
            .I(\this_vga_signals.CO0_0 ));
    Odrv12 I__2590 (
            .O(N__13370),
            .I(\this_vga_signals.CO0_0 ));
    Odrv4 I__2589 (
            .O(N__13365),
            .I(\this_vga_signals.CO0_0 ));
    LocalMux I__2588 (
            .O(N__13354),
            .I(\this_vga_signals.CO0_0 ));
    LocalMux I__2587 (
            .O(N__13347),
            .I(\this_vga_signals.CO0_0 ));
    Odrv4 I__2586 (
            .O(N__13344),
            .I(\this_vga_signals.CO0_0 ));
    CascadeMux I__2585 (
            .O(N__13331),
            .I(N__13328));
    CascadeBuf I__2584 (
            .O(N__13328),
            .I(N__13325));
    CascadeMux I__2583 (
            .O(N__13325),
            .I(N__13322));
    CascadeBuf I__2582 (
            .O(N__13322),
            .I(N__13319));
    CascadeMux I__2581 (
            .O(N__13319),
            .I(N__13316));
    CascadeBuf I__2580 (
            .O(N__13316),
            .I(N__13313));
    CascadeMux I__2579 (
            .O(N__13313),
            .I(N__13310));
    CascadeBuf I__2578 (
            .O(N__13310),
            .I(N__13307));
    CascadeMux I__2577 (
            .O(N__13307),
            .I(N__13304));
    CascadeBuf I__2576 (
            .O(N__13304),
            .I(N__13301));
    CascadeMux I__2575 (
            .O(N__13301),
            .I(N__13298));
    CascadeBuf I__2574 (
            .O(N__13298),
            .I(N__13295));
    CascadeMux I__2573 (
            .O(N__13295),
            .I(N__13292));
    CascadeBuf I__2572 (
            .O(N__13292),
            .I(N__13289));
    CascadeMux I__2571 (
            .O(N__13289),
            .I(N__13286));
    CascadeBuf I__2570 (
            .O(N__13286),
            .I(N__13283));
    CascadeMux I__2569 (
            .O(N__13283),
            .I(N__13280));
    CascadeBuf I__2568 (
            .O(N__13280),
            .I(N__13277));
    CascadeMux I__2567 (
            .O(N__13277),
            .I(N__13274));
    CascadeBuf I__2566 (
            .O(N__13274),
            .I(N__13271));
    CascadeMux I__2565 (
            .O(N__13271),
            .I(N__13268));
    CascadeBuf I__2564 (
            .O(N__13268),
            .I(N__13265));
    CascadeMux I__2563 (
            .O(N__13265),
            .I(N__13262));
    CascadeBuf I__2562 (
            .O(N__13262),
            .I(N__13259));
    CascadeMux I__2561 (
            .O(N__13259),
            .I(N__13256));
    CascadeBuf I__2560 (
            .O(N__13256),
            .I(N__13253));
    CascadeMux I__2559 (
            .O(N__13253),
            .I(N__13250));
    CascadeBuf I__2558 (
            .O(N__13250),
            .I(N__13247));
    CascadeMux I__2557 (
            .O(N__13247),
            .I(N__13244));
    CascadeBuf I__2556 (
            .O(N__13244),
            .I(N__13241));
    CascadeMux I__2555 (
            .O(N__13241),
            .I(N__13238));
    InMux I__2554 (
            .O(N__13238),
            .I(N__13235));
    LocalMux I__2553 (
            .O(N__13235),
            .I(N__13232));
    Span4Mux_v I__2552 (
            .O(N__13232),
            .I(N__13229));
    Span4Mux_v I__2551 (
            .O(N__13229),
            .I(N__13226));
    Span4Mux_v I__2550 (
            .O(N__13226),
            .I(N__13223));
    Span4Mux_v I__2549 (
            .O(N__13223),
            .I(N__13220));
    Odrv4 I__2548 (
            .O(N__13220),
            .I(M_haddress_q_RNI8ARU_11));
    InMux I__2547 (
            .O(N__13217),
            .I(N__13214));
    LocalMux I__2546 (
            .O(N__13214),
            .I(N__13210));
    InMux I__2545 (
            .O(N__13213),
            .I(N__13205));
    Span4Mux_h I__2544 (
            .O(N__13210),
            .I(N__13202));
    InMux I__2543 (
            .O(N__13209),
            .I(N__13199));
    InMux I__2542 (
            .O(N__13208),
            .I(N__13196));
    LocalMux I__2541 (
            .O(N__13205),
            .I(M_state_qZ0Z_1));
    Odrv4 I__2540 (
            .O(N__13202),
            .I(M_state_qZ0Z_1));
    LocalMux I__2539 (
            .O(N__13199),
            .I(M_state_qZ0Z_1));
    LocalMux I__2538 (
            .O(N__13196),
            .I(M_state_qZ0Z_1));
    CascadeMux I__2537 (
            .O(N__13187),
            .I(N__13181));
    CascadeMux I__2536 (
            .O(N__13186),
            .I(N__13177));
    InMux I__2535 (
            .O(N__13185),
            .I(N__13174));
    InMux I__2534 (
            .O(N__13184),
            .I(N__13169));
    InMux I__2533 (
            .O(N__13181),
            .I(N__13169));
    CascadeMux I__2532 (
            .O(N__13180),
            .I(N__13162));
    InMux I__2531 (
            .O(N__13177),
            .I(N__13159));
    LocalMux I__2530 (
            .O(N__13174),
            .I(N__13154));
    LocalMux I__2529 (
            .O(N__13169),
            .I(N__13154));
    InMux I__2528 (
            .O(N__13168),
            .I(N__13149));
    InMux I__2527 (
            .O(N__13167),
            .I(N__13149));
    InMux I__2526 (
            .O(N__13166),
            .I(N__13146));
    InMux I__2525 (
            .O(N__13165),
            .I(N__13143));
    InMux I__2524 (
            .O(N__13162),
            .I(N__13140));
    LocalMux I__2523 (
            .O(N__13159),
            .I(N__13137));
    Span4Mux_v I__2522 (
            .O(N__13154),
            .I(N__13134));
    LocalMux I__2521 (
            .O(N__13149),
            .I(N__13129));
    LocalMux I__2520 (
            .O(N__13146),
            .I(N__13129));
    LocalMux I__2519 (
            .O(N__13143),
            .I(N__13124));
    LocalMux I__2518 (
            .O(N__13140),
            .I(N__13124));
    Span4Mux_v I__2517 (
            .O(N__13137),
            .I(N__13121));
    Span4Mux_h I__2516 (
            .O(N__13134),
            .I(N__13118));
    Span4Mux_v I__2515 (
            .O(N__13129),
            .I(N__13115));
    Span12Mux_v I__2514 (
            .O(N__13124),
            .I(N__13110));
    Sp12to4 I__2513 (
            .O(N__13121),
            .I(N__13110));
    Sp12to4 I__2512 (
            .O(N__13118),
            .I(N__13105));
    Sp12to4 I__2511 (
            .O(N__13115),
            .I(N__13105));
    Span12Mux_h I__2510 (
            .O(N__13110),
            .I(N__13102));
    Span12Mux_h I__2509 (
            .O(N__13105),
            .I(N__13099));
    Odrv12 I__2508 (
            .O(N__13102),
            .I(port_enb_c));
    Odrv12 I__2507 (
            .O(N__13099),
            .I(port_enb_c));
    InMux I__2506 (
            .O(N__13094),
            .I(N__13088));
    InMux I__2505 (
            .O(N__13093),
            .I(N__13085));
    InMux I__2504 (
            .O(N__13092),
            .I(N__13082));
    InMux I__2503 (
            .O(N__13091),
            .I(N__13079));
    LocalMux I__2502 (
            .O(N__13088),
            .I(N__13074));
    LocalMux I__2501 (
            .O(N__13085),
            .I(N__13074));
    LocalMux I__2500 (
            .O(N__13082),
            .I(M_state_qZ0Z_3));
    LocalMux I__2499 (
            .O(N__13079),
            .I(M_state_qZ0Z_3));
    Odrv4 I__2498 (
            .O(N__13074),
            .I(M_state_qZ0Z_3));
    InMux I__2497 (
            .O(N__13067),
            .I(N__13059));
    InMux I__2496 (
            .O(N__13066),
            .I(N__13056));
    InMux I__2495 (
            .O(N__13065),
            .I(N__13053));
    InMux I__2494 (
            .O(N__13064),
            .I(N__13047));
    InMux I__2493 (
            .O(N__13063),
            .I(N__13047));
    InMux I__2492 (
            .O(N__13062),
            .I(N__13042));
    LocalMux I__2491 (
            .O(N__13059),
            .I(N__13039));
    LocalMux I__2490 (
            .O(N__13056),
            .I(N__13034));
    LocalMux I__2489 (
            .O(N__13053),
            .I(N__13034));
    InMux I__2488 (
            .O(N__13052),
            .I(N__13031));
    LocalMux I__2487 (
            .O(N__13047),
            .I(N__13028));
    InMux I__2486 (
            .O(N__13046),
            .I(N__13023));
    InMux I__2485 (
            .O(N__13045),
            .I(N__13023));
    LocalMux I__2484 (
            .O(N__13042),
            .I(N__13018));
    Span4Mux_h I__2483 (
            .O(N__13039),
            .I(N__13018));
    Span4Mux_h I__2482 (
            .O(N__13034),
            .I(N__13015));
    LocalMux I__2481 (
            .O(N__13031),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__2480 (
            .O(N__13028),
            .I(M_this_start_data_delay_out_0));
    LocalMux I__2479 (
            .O(N__13023),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__2478 (
            .O(N__13018),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__2477 (
            .O(N__13015),
            .I(M_this_start_data_delay_out_0));
    InMux I__2476 (
            .O(N__13004),
            .I(N__12998));
    InMux I__2475 (
            .O(N__13003),
            .I(N__12998));
    LocalMux I__2474 (
            .O(N__12998),
            .I(\this_vga_signals.M_vaddress_q_fastZ0Z_5 ));
    InMux I__2473 (
            .O(N__12995),
            .I(N__12991));
    CascadeMux I__2472 (
            .O(N__12994),
            .I(N__12985));
    LocalMux I__2471 (
            .O(N__12991),
            .I(N__12982));
    InMux I__2470 (
            .O(N__12990),
            .I(N__12975));
    InMux I__2469 (
            .O(N__12989),
            .I(N__12975));
    InMux I__2468 (
            .O(N__12988),
            .I(N__12975));
    InMux I__2467 (
            .O(N__12985),
            .I(N__12972));
    Odrv4 I__2466 (
            .O(N__12982),
            .I(\this_vga_signals.M_vaddress_q_fastZ0Z_9 ));
    LocalMux I__2465 (
            .O(N__12975),
            .I(\this_vga_signals.M_vaddress_q_fastZ0Z_9 ));
    LocalMux I__2464 (
            .O(N__12972),
            .I(\this_vga_signals.M_vaddress_q_fastZ0Z_9 ));
    CascadeMux I__2463 (
            .O(N__12965),
            .I(N__12958));
    CascadeMux I__2462 (
            .O(N__12964),
            .I(N__12955));
    CascadeMux I__2461 (
            .O(N__12963),
            .I(N__12952));
    InMux I__2460 (
            .O(N__12962),
            .I(N__12949));
    InMux I__2459 (
            .O(N__12961),
            .I(N__12940));
    InMux I__2458 (
            .O(N__12958),
            .I(N__12940));
    InMux I__2457 (
            .O(N__12955),
            .I(N__12940));
    InMux I__2456 (
            .O(N__12952),
            .I(N__12940));
    LocalMux I__2455 (
            .O(N__12949),
            .I(\this_vga_signals.M_vaddress_q_fastZ0Z_8 ));
    LocalMux I__2454 (
            .O(N__12940),
            .I(\this_vga_signals.M_vaddress_q_fastZ0Z_8 ));
    InMux I__2453 (
            .O(N__12935),
            .I(N__12931));
    InMux I__2452 (
            .O(N__12934),
            .I(N__12928));
    LocalMux I__2451 (
            .O(N__12931),
            .I(\this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8 ));
    LocalMux I__2450 (
            .O(N__12928),
            .I(\this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8 ));
    CascadeMux I__2449 (
            .O(N__12923),
            .I(\this_vga_signals.N_353_0_cascade_ ));
    InMux I__2448 (
            .O(N__12920),
            .I(N__12912));
    InMux I__2447 (
            .O(N__12919),
            .I(N__12912));
    InMux I__2446 (
            .O(N__12918),
            .I(N__12907));
    InMux I__2445 (
            .O(N__12917),
            .I(N__12907));
    LocalMux I__2444 (
            .O(N__12912),
            .I(\this_vga_signals.mult1_un40_sum_m_bm_2 ));
    LocalMux I__2443 (
            .O(N__12907),
            .I(\this_vga_signals.mult1_un40_sum_m_bm_2 ));
    CascadeMux I__2442 (
            .O(N__12902),
            .I(\this_vga_signals.mult1_un40_sum_0_axbxc3_5_1_0_cascade_ ));
    InMux I__2441 (
            .O(N__12899),
            .I(N__12896));
    LocalMux I__2440 (
            .O(N__12896),
            .I(\this_vga_signals.mult1_un40_sum_0_axbxc3_5_3 ));
    InMux I__2439 (
            .O(N__12893),
            .I(N__12887));
    InMux I__2438 (
            .O(N__12892),
            .I(N__12887));
    LocalMux I__2437 (
            .O(N__12887),
            .I(N__12883));
    InMux I__2436 (
            .O(N__12886),
            .I(N__12878));
    Span4Mux_h I__2435 (
            .O(N__12883),
            .I(N__12875));
    InMux I__2434 (
            .O(N__12882),
            .I(N__12870));
    InMux I__2433 (
            .O(N__12881),
            .I(N__12870));
    LocalMux I__2432 (
            .O(N__12878),
            .I(\this_vga_signals.mult1_un40_sum0_3 ));
    Odrv4 I__2431 (
            .O(N__12875),
            .I(\this_vga_signals.mult1_un40_sum0_3 ));
    LocalMux I__2430 (
            .O(N__12870),
            .I(\this_vga_signals.mult1_un40_sum0_3 ));
    InMux I__2429 (
            .O(N__12863),
            .I(N__12852));
    InMux I__2428 (
            .O(N__12862),
            .I(N__12852));
    InMux I__2427 (
            .O(N__12861),
            .I(N__12845));
    InMux I__2426 (
            .O(N__12860),
            .I(N__12845));
    InMux I__2425 (
            .O(N__12859),
            .I(N__12845));
    InMux I__2424 (
            .O(N__12858),
            .I(N__12840));
    InMux I__2423 (
            .O(N__12857),
            .I(N__12840));
    LocalMux I__2422 (
            .O(N__12852),
            .I(\this_vga_signals.M_vaddress_q_5_repZ0Z1 ));
    LocalMux I__2421 (
            .O(N__12845),
            .I(\this_vga_signals.M_vaddress_q_5_repZ0Z1 ));
    LocalMux I__2420 (
            .O(N__12840),
            .I(\this_vga_signals.M_vaddress_q_5_repZ0Z1 ));
    CascadeMux I__2419 (
            .O(N__12833),
            .I(N__12830));
    InMux I__2418 (
            .O(N__12830),
            .I(N__12827));
    LocalMux I__2417 (
            .O(N__12827),
            .I(N__12824));
    Span4Mux_v I__2416 (
            .O(N__12824),
            .I(N__12821));
    Odrv4 I__2415 (
            .O(N__12821),
            .I(\this_vga_signals.mult1_un40_sum_0_axb1 ));
    InMux I__2414 (
            .O(N__12818),
            .I(N__12815));
    LocalMux I__2413 (
            .O(N__12815),
            .I(\this_vga_signals.mult1_un40_sum_m_1_1 ));
    CascadeMux I__2412 (
            .O(N__12812),
            .I(\this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8_cascade_ ));
    InMux I__2411 (
            .O(N__12809),
            .I(N__12805));
    CascadeMux I__2410 (
            .O(N__12808),
            .I(N__12801));
    LocalMux I__2409 (
            .O(N__12805),
            .I(N__12798));
    InMux I__2408 (
            .O(N__12804),
            .I(N__12795));
    InMux I__2407 (
            .O(N__12801),
            .I(N__12792));
    Span4Mux_v I__2406 (
            .O(N__12798),
            .I(N__12787));
    LocalMux I__2405 (
            .O(N__12795),
            .I(N__12787));
    LocalMux I__2404 (
            .O(N__12792),
            .I(\this_vga_signals.mult1_un40_sum_m_0_1 ));
    Odrv4 I__2403 (
            .O(N__12787),
            .I(\this_vga_signals.mult1_un40_sum_m_0_1 ));
    CascadeMux I__2402 (
            .O(N__12782),
            .I(N__12779));
    InMux I__2401 (
            .O(N__12779),
            .I(N__12775));
    InMux I__2400 (
            .O(N__12778),
            .I(N__12772));
    LocalMux I__2399 (
            .O(N__12775),
            .I(\this_vga_signals.M_vaddress_q_fastZ0Z_6 ));
    LocalMux I__2398 (
            .O(N__12772),
            .I(\this_vga_signals.M_vaddress_q_fastZ0Z_6 ));
    CascadeMux I__2397 (
            .O(N__12767),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_2_0_cascade_ ));
    CascadeMux I__2396 (
            .O(N__12764),
            .I(N__12760));
    InMux I__2395 (
            .O(N__12763),
            .I(N__12757));
    InMux I__2394 (
            .O(N__12760),
            .I(N__12754));
    LocalMux I__2393 (
            .O(N__12757),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_2 ));
    LocalMux I__2392 (
            .O(N__12754),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_2 ));
    CascadeMux I__2391 (
            .O(N__12749),
            .I(N__12746));
    InMux I__2390 (
            .O(N__12746),
            .I(N__12743));
    LocalMux I__2389 (
            .O(N__12743),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_a4_1_0 ));
    InMux I__2388 (
            .O(N__12740),
            .I(N__12734));
    InMux I__2387 (
            .O(N__12739),
            .I(N__12731));
    InMux I__2386 (
            .O(N__12738),
            .I(N__12726));
    InMux I__2385 (
            .O(N__12737),
            .I(N__12726));
    LocalMux I__2384 (
            .O(N__12734),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_2_0 ));
    LocalMux I__2383 (
            .O(N__12731),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_2_0 ));
    LocalMux I__2382 (
            .O(N__12726),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_2_0 ));
    InMux I__2381 (
            .O(N__12719),
            .I(N__12714));
    InMux I__2380 (
            .O(N__12718),
            .I(N__12711));
    InMux I__2379 (
            .O(N__12717),
            .I(N__12708));
    LocalMux I__2378 (
            .O(N__12714),
            .I(\this_vga_signals.if_m5_0_s ));
    LocalMux I__2377 (
            .O(N__12711),
            .I(\this_vga_signals.if_m5_0_s ));
    LocalMux I__2376 (
            .O(N__12708),
            .I(\this_vga_signals.if_m5_0_s ));
    InMux I__2375 (
            .O(N__12701),
            .I(N__12696));
    InMux I__2374 (
            .O(N__12700),
            .I(N__12693));
    InMux I__2373 (
            .O(N__12699),
            .I(N__12690));
    LocalMux I__2372 (
            .O(N__12696),
            .I(\this_vga_signals.if_m1_0 ));
    LocalMux I__2371 (
            .O(N__12693),
            .I(\this_vga_signals.if_m1_0 ));
    LocalMux I__2370 (
            .O(N__12690),
            .I(\this_vga_signals.if_m1_0 ));
    CascadeMux I__2369 (
            .O(N__12683),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ));
    CascadeMux I__2368 (
            .O(N__12680),
            .I(\this_vga_signals.if_N_2_2_cascade_ ));
    InMux I__2367 (
            .O(N__12677),
            .I(N__12674));
    LocalMux I__2366 (
            .O(N__12674),
            .I(N__12670));
    InMux I__2365 (
            .O(N__12673),
            .I(N__12667));
    Span4Mux_v I__2364 (
            .O(N__12670),
            .I(N__12664));
    LocalMux I__2363 (
            .O(N__12667),
            .I(\this_vga_signals.mult1_un54_sum_axb1_3 ));
    Odrv4 I__2362 (
            .O(N__12664),
            .I(\this_vga_signals.mult1_un54_sum_axb1_3 ));
    InMux I__2361 (
            .O(N__12659),
            .I(N__12656));
    LocalMux I__2360 (
            .O(N__12656),
            .I(N__12653));
    Span4Mux_h I__2359 (
            .O(N__12653),
            .I(N__12650));
    Odrv4 I__2358 (
            .O(N__12650),
            .I(\this_vga_signals.mult1_un61_sum_c3_1_0 ));
    InMux I__2357 (
            .O(N__12647),
            .I(N__12642));
    InMux I__2356 (
            .O(N__12646),
            .I(N__12637));
    InMux I__2355 (
            .O(N__12645),
            .I(N__12637));
    LocalMux I__2354 (
            .O(N__12642),
            .I(M_state_qZ0Z_2));
    LocalMux I__2353 (
            .O(N__12637),
            .I(M_state_qZ0Z_2));
    InMux I__2352 (
            .O(N__12632),
            .I(N__12624));
    InMux I__2351 (
            .O(N__12631),
            .I(N__12615));
    InMux I__2350 (
            .O(N__12630),
            .I(N__12615));
    InMux I__2349 (
            .O(N__12629),
            .I(N__12612));
    InMux I__2348 (
            .O(N__12628),
            .I(N__12609));
    InMux I__2347 (
            .O(N__12627),
            .I(N__12602));
    LocalMux I__2346 (
            .O(N__12624),
            .I(N__12599));
    CascadeMux I__2345 (
            .O(N__12623),
            .I(N__12595));
    InMux I__2344 (
            .O(N__12622),
            .I(N__12588));
    InMux I__2343 (
            .O(N__12621),
            .I(N__12588));
    InMux I__2342 (
            .O(N__12620),
            .I(N__12581));
    LocalMux I__2341 (
            .O(N__12615),
            .I(N__12576));
    LocalMux I__2340 (
            .O(N__12612),
            .I(N__12576));
    LocalMux I__2339 (
            .O(N__12609),
            .I(N__12573));
    InMux I__2338 (
            .O(N__12608),
            .I(N__12568));
    InMux I__2337 (
            .O(N__12607),
            .I(N__12568));
    InMux I__2336 (
            .O(N__12606),
            .I(N__12565));
    CascadeMux I__2335 (
            .O(N__12605),
            .I(N__12560));
    LocalMux I__2334 (
            .O(N__12602),
            .I(N__12549));
    Span12Mux_h I__2333 (
            .O(N__12599),
            .I(N__12549));
    InMux I__2332 (
            .O(N__12598),
            .I(N__12546));
    InMux I__2331 (
            .O(N__12595),
            .I(N__12541));
    InMux I__2330 (
            .O(N__12594),
            .I(N__12541));
    InMux I__2329 (
            .O(N__12593),
            .I(N__12538));
    LocalMux I__2328 (
            .O(N__12588),
            .I(N__12535));
    InMux I__2327 (
            .O(N__12587),
            .I(N__12526));
    InMux I__2326 (
            .O(N__12586),
            .I(N__12526));
    InMux I__2325 (
            .O(N__12585),
            .I(N__12526));
    InMux I__2324 (
            .O(N__12584),
            .I(N__12526));
    LocalMux I__2323 (
            .O(N__12581),
            .I(N__12519));
    Span4Mux_v I__2322 (
            .O(N__12576),
            .I(N__12519));
    Span4Mux_v I__2321 (
            .O(N__12573),
            .I(N__12519));
    LocalMux I__2320 (
            .O(N__12568),
            .I(N__12514));
    LocalMux I__2319 (
            .O(N__12565),
            .I(N__12514));
    InMux I__2318 (
            .O(N__12564),
            .I(N__12509));
    InMux I__2317 (
            .O(N__12563),
            .I(N__12509));
    InMux I__2316 (
            .O(N__12560),
            .I(N__12502));
    InMux I__2315 (
            .O(N__12559),
            .I(N__12502));
    InMux I__2314 (
            .O(N__12558),
            .I(N__12502));
    InMux I__2313 (
            .O(N__12557),
            .I(N__12495));
    InMux I__2312 (
            .O(N__12556),
            .I(N__12495));
    InMux I__2311 (
            .O(N__12555),
            .I(N__12495));
    InMux I__2310 (
            .O(N__12554),
            .I(N__12492));
    Odrv12 I__2309 (
            .O(N__12549),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2308 (
            .O(N__12546),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2307 (
            .O(N__12541),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2306 (
            .O(N__12538),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    Odrv4 I__2305 (
            .O(N__12535),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2304 (
            .O(N__12526),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    Odrv4 I__2303 (
            .O(N__12519),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    Odrv4 I__2302 (
            .O(N__12514),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2301 (
            .O(N__12509),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2300 (
            .O(N__12502),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2299 (
            .O(N__12495),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2298 (
            .O(N__12492),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    InMux I__2297 (
            .O(N__12467),
            .I(N__12464));
    LocalMux I__2296 (
            .O(N__12464),
            .I(N__12461));
    Sp12to4 I__2295 (
            .O(N__12461),
            .I(N__12458));
    Span12Mux_v I__2294 (
            .O(N__12458),
            .I(N__12451));
    InMux I__2293 (
            .O(N__12457),
            .I(N__12446));
    InMux I__2292 (
            .O(N__12456),
            .I(N__12446));
    InMux I__2291 (
            .O(N__12455),
            .I(N__12443));
    InMux I__2290 (
            .O(N__12454),
            .I(N__12440));
    Odrv12 I__2289 (
            .O(N__12451),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__2288 (
            .O(N__12446),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__2287 (
            .O(N__12443),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__2286 (
            .O(N__12440),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    CascadeMux I__2285 (
            .O(N__12431),
            .I(N__12428));
    InMux I__2284 (
            .O(N__12428),
            .I(N__12424));
    CascadeMux I__2283 (
            .O(N__12427),
            .I(N__12421));
    LocalMux I__2282 (
            .O(N__12424),
            .I(N__12417));
    InMux I__2281 (
            .O(N__12421),
            .I(N__12413));
    CascadeMux I__2280 (
            .O(N__12420),
            .I(N__12409));
    Span4Mux_v I__2279 (
            .O(N__12417),
            .I(N__12406));
    InMux I__2278 (
            .O(N__12416),
            .I(N__12403));
    LocalMux I__2277 (
            .O(N__12413),
            .I(N__12400));
    InMux I__2276 (
            .O(N__12412),
            .I(N__12393));
    InMux I__2275 (
            .O(N__12409),
            .I(N__12393));
    Span4Mux_v I__2274 (
            .O(N__12406),
            .I(N__12388));
    LocalMux I__2273 (
            .O(N__12403),
            .I(N__12388));
    Span4Mux_v I__2272 (
            .O(N__12400),
            .I(N__12385));
    InMux I__2271 (
            .O(N__12399),
            .I(N__12380));
    InMux I__2270 (
            .O(N__12398),
            .I(N__12380));
    LocalMux I__2269 (
            .O(N__12393),
            .I(N__12377));
    Odrv4 I__2268 (
            .O(N__12388),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1 ));
    Odrv4 I__2267 (
            .O(N__12385),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1 ));
    LocalMux I__2266 (
            .O(N__12380),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1 ));
    Odrv4 I__2265 (
            .O(N__12377),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1 ));
    InMux I__2264 (
            .O(N__12368),
            .I(N__12364));
    InMux I__2263 (
            .O(N__12367),
            .I(N__12359));
    LocalMux I__2262 (
            .O(N__12364),
            .I(N__12349));
    InMux I__2261 (
            .O(N__12363),
            .I(N__12343));
    InMux I__2260 (
            .O(N__12362),
            .I(N__12343));
    LocalMux I__2259 (
            .O(N__12359),
            .I(N__12340));
    InMux I__2258 (
            .O(N__12358),
            .I(N__12337));
    InMux I__2257 (
            .O(N__12357),
            .I(N__12332));
    InMux I__2256 (
            .O(N__12356),
            .I(N__12332));
    InMux I__2255 (
            .O(N__12355),
            .I(N__12329));
    InMux I__2254 (
            .O(N__12354),
            .I(N__12324));
    InMux I__2253 (
            .O(N__12353),
            .I(N__12324));
    InMux I__2252 (
            .O(N__12352),
            .I(N__12319));
    Span4Mux_v I__2251 (
            .O(N__12349),
            .I(N__12306));
    InMux I__2250 (
            .O(N__12348),
            .I(N__12303));
    LocalMux I__2249 (
            .O(N__12343),
            .I(N__12298));
    Span4Mux_v I__2248 (
            .O(N__12340),
            .I(N__12298));
    LocalMux I__2247 (
            .O(N__12337),
            .I(N__12295));
    LocalMux I__2246 (
            .O(N__12332),
            .I(N__12292));
    LocalMux I__2245 (
            .O(N__12329),
            .I(N__12279));
    LocalMux I__2244 (
            .O(N__12324),
            .I(N__12279));
    InMux I__2243 (
            .O(N__12323),
            .I(N__12274));
    InMux I__2242 (
            .O(N__12322),
            .I(N__12274));
    LocalMux I__2241 (
            .O(N__12319),
            .I(N__12271));
    InMux I__2240 (
            .O(N__12318),
            .I(N__12266));
    InMux I__2239 (
            .O(N__12317),
            .I(N__12266));
    InMux I__2238 (
            .O(N__12316),
            .I(N__12259));
    InMux I__2237 (
            .O(N__12315),
            .I(N__12259));
    InMux I__2236 (
            .O(N__12314),
            .I(N__12259));
    InMux I__2235 (
            .O(N__12313),
            .I(N__12256));
    InMux I__2234 (
            .O(N__12312),
            .I(N__12247));
    InMux I__2233 (
            .O(N__12311),
            .I(N__12247));
    InMux I__2232 (
            .O(N__12310),
            .I(N__12247));
    InMux I__2231 (
            .O(N__12309),
            .I(N__12247));
    Span4Mux_v I__2230 (
            .O(N__12306),
            .I(N__12236));
    LocalMux I__2229 (
            .O(N__12303),
            .I(N__12236));
    Span4Mux_h I__2228 (
            .O(N__12298),
            .I(N__12236));
    Span4Mux_v I__2227 (
            .O(N__12295),
            .I(N__12236));
    Span4Mux_v I__2226 (
            .O(N__12292),
            .I(N__12236));
    InMux I__2225 (
            .O(N__12291),
            .I(N__12229));
    InMux I__2224 (
            .O(N__12290),
            .I(N__12229));
    InMux I__2223 (
            .O(N__12289),
            .I(N__12229));
    InMux I__2222 (
            .O(N__12288),
            .I(N__12226));
    InMux I__2221 (
            .O(N__12287),
            .I(N__12217));
    InMux I__2220 (
            .O(N__12286),
            .I(N__12217));
    InMux I__2219 (
            .O(N__12285),
            .I(N__12217));
    InMux I__2218 (
            .O(N__12284),
            .I(N__12217));
    Odrv4 I__2217 (
            .O(N__12279),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2216 (
            .O(N__12274),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    Odrv4 I__2215 (
            .O(N__12271),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2214 (
            .O(N__12266),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2213 (
            .O(N__12259),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2212 (
            .O(N__12256),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2211 (
            .O(N__12247),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    Odrv4 I__2210 (
            .O(N__12236),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2209 (
            .O(N__12229),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2208 (
            .O(N__12226),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2207 (
            .O(N__12217),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    CascadeMux I__2206 (
            .O(N__12194),
            .I(N__12191));
    CascadeBuf I__2205 (
            .O(N__12191),
            .I(N__12188));
    CascadeMux I__2204 (
            .O(N__12188),
            .I(N__12185));
    CascadeBuf I__2203 (
            .O(N__12185),
            .I(N__12182));
    CascadeMux I__2202 (
            .O(N__12182),
            .I(N__12179));
    CascadeBuf I__2201 (
            .O(N__12179),
            .I(N__12176));
    CascadeMux I__2200 (
            .O(N__12176),
            .I(N__12173));
    CascadeBuf I__2199 (
            .O(N__12173),
            .I(N__12170));
    CascadeMux I__2198 (
            .O(N__12170),
            .I(N__12167));
    CascadeBuf I__2197 (
            .O(N__12167),
            .I(N__12164));
    CascadeMux I__2196 (
            .O(N__12164),
            .I(N__12161));
    CascadeBuf I__2195 (
            .O(N__12161),
            .I(N__12158));
    CascadeMux I__2194 (
            .O(N__12158),
            .I(N__12155));
    CascadeBuf I__2193 (
            .O(N__12155),
            .I(N__12152));
    CascadeMux I__2192 (
            .O(N__12152),
            .I(N__12149));
    CascadeBuf I__2191 (
            .O(N__12149),
            .I(N__12146));
    CascadeMux I__2190 (
            .O(N__12146),
            .I(N__12143));
    CascadeBuf I__2189 (
            .O(N__12143),
            .I(N__12140));
    CascadeMux I__2188 (
            .O(N__12140),
            .I(N__12137));
    CascadeBuf I__2187 (
            .O(N__12137),
            .I(N__12134));
    CascadeMux I__2186 (
            .O(N__12134),
            .I(N__12131));
    CascadeBuf I__2185 (
            .O(N__12131),
            .I(N__12128));
    CascadeMux I__2184 (
            .O(N__12128),
            .I(N__12125));
    CascadeBuf I__2183 (
            .O(N__12125),
            .I(N__12122));
    CascadeMux I__2182 (
            .O(N__12122),
            .I(N__12119));
    CascadeBuf I__2181 (
            .O(N__12119),
            .I(N__12116));
    CascadeMux I__2180 (
            .O(N__12116),
            .I(N__12113));
    CascadeBuf I__2179 (
            .O(N__12113),
            .I(N__12110));
    CascadeMux I__2178 (
            .O(N__12110),
            .I(N__12107));
    CascadeBuf I__2177 (
            .O(N__12107),
            .I(N__12104));
    CascadeMux I__2176 (
            .O(N__12104),
            .I(N__12101));
    InMux I__2175 (
            .O(N__12101),
            .I(N__12098));
    LocalMux I__2174 (
            .O(N__12098),
            .I(N__12095));
    Span4Mux_v I__2173 (
            .O(N__12095),
            .I(N__12092));
    Span4Mux_h I__2172 (
            .O(N__12092),
            .I(N__12089));
    Sp12to4 I__2171 (
            .O(N__12089),
            .I(N__12086));
    Odrv12 I__2170 (
            .O(N__12086),
            .I(this_vga_signals_un14_address_if_generate_plus_mult1_un54_sum_i_3));
    InMux I__2169 (
            .O(N__12083),
            .I(N__12079));
    InMux I__2168 (
            .O(N__12082),
            .I(N__12076));
    LocalMux I__2167 (
            .O(N__12079),
            .I(N__12073));
    LocalMux I__2166 (
            .O(N__12076),
            .I(N__12068));
    Span4Mux_v I__2165 (
            .O(N__12073),
            .I(N__12068));
    Odrv4 I__2164 (
            .O(N__12068),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_4 ));
    InMux I__2163 (
            .O(N__12065),
            .I(N__12062));
    LocalMux I__2162 (
            .O(N__12062),
            .I(\this_vga_signals.M_vaddress_q_fastZ0Z_7 ));
    CascadeMux I__2161 (
            .O(N__12059),
            .I(\this_vga_signals.mult1_un40_sum_m_am_x_2_cascade_ ));
    InMux I__2160 (
            .O(N__12056),
            .I(N__12052));
    InMux I__2159 (
            .O(N__12055),
            .I(N__12049));
    LocalMux I__2158 (
            .O(N__12052),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_2 ));
    LocalMux I__2157 (
            .O(N__12049),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_2 ));
    InMux I__2156 (
            .O(N__12044),
            .I(N__12040));
    InMux I__2155 (
            .O(N__12043),
            .I(N__12037));
    LocalMux I__2154 (
            .O(N__12040),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_3 ));
    LocalMux I__2153 (
            .O(N__12037),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_3 ));
    CascadeMux I__2152 (
            .O(N__12032),
            .I(\this_vga_signals.mult1_un40_sum_m_x1_3_cascade_ ));
    CascadeMux I__2151 (
            .O(N__12029),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3_cascade_ ));
    InMux I__2150 (
            .O(N__12026),
            .I(N__12023));
    LocalMux I__2149 (
            .O(N__12023),
            .I(\this_vga_signals.N_6_i ));
    CascadeMux I__2148 (
            .O(N__12020),
            .I(N__12016));
    InMux I__2147 (
            .O(N__12019),
            .I(N__12012));
    InMux I__2146 (
            .O(N__12016),
            .I(N__12007));
    InMux I__2145 (
            .O(N__12015),
            .I(N__12007));
    LocalMux I__2144 (
            .O(N__12012),
            .I(N__12004));
    LocalMux I__2143 (
            .O(N__12007),
            .I(\this_vga_signals.mult1_un40_sum_m_am_2 ));
    Odrv4 I__2142 (
            .O(N__12004),
            .I(\this_vga_signals.mult1_un40_sum_m_am_2 ));
    InMux I__2141 (
            .O(N__11999),
            .I(N__11996));
    LocalMux I__2140 (
            .O(N__11996),
            .I(N__11992));
    InMux I__2139 (
            .O(N__11995),
            .I(N__11989));
    Span4Mux_h I__2138 (
            .O(N__11992),
            .I(N__11986));
    LocalMux I__2137 (
            .O(N__11989),
            .I(\this_vga_signals.mult1_un40_sum1_3 ));
    Odrv4 I__2136 (
            .O(N__11986),
            .I(\this_vga_signals.mult1_un40_sum1_3 ));
    InMux I__2135 (
            .O(N__11981),
            .I(N__11978));
    LocalMux I__2134 (
            .O(N__11978),
            .I(\this_vga_signals.N_6_i_0 ));
    CascadeMux I__2133 (
            .O(N__11975),
            .I(\this_vga_signals.mult1_un40_sum1_3_cascade_ ));
    InMux I__2132 (
            .O(N__11972),
            .I(N__11969));
    LocalMux I__2131 (
            .O(N__11969),
            .I(\this_vga_signals.g0_4_0 ));
    CascadeMux I__2130 (
            .O(N__11966),
            .I(N__11963));
    InMux I__2129 (
            .O(N__11963),
            .I(N__11959));
    InMux I__2128 (
            .O(N__11962),
            .I(N__11955));
    LocalMux I__2127 (
            .O(N__11959),
            .I(N__11952));
    InMux I__2126 (
            .O(N__11958),
            .I(N__11949));
    LocalMux I__2125 (
            .O(N__11955),
            .I(N__11942));
    Span4Mux_h I__2124 (
            .O(N__11952),
            .I(N__11942));
    LocalMux I__2123 (
            .O(N__11949),
            .I(N__11942));
    Span4Mux_v I__2122 (
            .O(N__11942),
            .I(N__11936));
    InMux I__2121 (
            .O(N__11941),
            .I(N__11933));
    InMux I__2120 (
            .O(N__11940),
            .I(N__11930));
    InMux I__2119 (
            .O(N__11939),
            .I(N__11927));
    Sp12to4 I__2118 (
            .O(N__11936),
            .I(N__11924));
    LocalMux I__2117 (
            .O(N__11933),
            .I(N__11917));
    LocalMux I__2116 (
            .O(N__11930),
            .I(N__11917));
    LocalMux I__2115 (
            .O(N__11927),
            .I(N__11917));
    Span12Mux_h I__2114 (
            .O(N__11924),
            .I(N__11914));
    Span12Mux_v I__2113 (
            .O(N__11917),
            .I(N__11911));
    Odrv12 I__2112 (
            .O(N__11914),
            .I(M_this_vram_read_data_1));
    Odrv12 I__2111 (
            .O(N__11911),
            .I(M_this_vram_read_data_1));
    CascadeMux I__2110 (
            .O(N__11906),
            .I(\this_vga_signals.g0_1_1_1_cascade_ ));
    InMux I__2109 (
            .O(N__11903),
            .I(N__11900));
    LocalMux I__2108 (
            .O(N__11900),
            .I(\this_vga_signals.g0_3_0_0 ));
    InMux I__2107 (
            .O(N__11897),
            .I(N__11893));
    CascadeMux I__2106 (
            .O(N__11896),
            .I(N__11890));
    LocalMux I__2105 (
            .O(N__11893),
            .I(N__11887));
    InMux I__2104 (
            .O(N__11890),
            .I(N__11884));
    Odrv4 I__2103 (
            .O(N__11887),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_1 ));
    LocalMux I__2102 (
            .O(N__11884),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_1 ));
    InMux I__2101 (
            .O(N__11879),
            .I(N__11876));
    LocalMux I__2100 (
            .O(N__11876),
            .I(\this_vga_signals.N_2_1_0 ));
    InMux I__2099 (
            .O(N__11873),
            .I(N__11870));
    LocalMux I__2098 (
            .O(N__11870),
            .I(\this_vga_signals.g0_3_2_1 ));
    CascadeMux I__2097 (
            .O(N__11867),
            .I(\this_start_data_delay.this_edge_detector.N_263_cascade_ ));
    InMux I__2096 (
            .O(N__11864),
            .I(N__11857));
    InMux I__2095 (
            .O(N__11863),
            .I(N__11857));
    InMux I__2094 (
            .O(N__11862),
            .I(N__11854));
    LocalMux I__2093 (
            .O(N__11857),
            .I(M_state_qZ0Z_0));
    LocalMux I__2092 (
            .O(N__11854),
            .I(M_state_qZ0Z_0));
    InMux I__2091 (
            .O(N__11849),
            .I(N__11843));
    InMux I__2090 (
            .O(N__11848),
            .I(N__11843));
    LocalMux I__2089 (
            .O(N__11843),
            .I(N__11838));
    InMux I__2088 (
            .O(N__11842),
            .I(N__11833));
    InMux I__2087 (
            .O(N__11841),
            .I(N__11833));
    Span4Mux_h I__2086 (
            .O(N__11838),
            .I(N__11828));
    LocalMux I__2085 (
            .O(N__11833),
            .I(N__11828));
    Span4Mux_v I__2084 (
            .O(N__11828),
            .I(N__11825));
    Span4Mux_v I__2083 (
            .O(N__11825),
            .I(N__11822));
    Span4Mux_v I__2082 (
            .O(N__11822),
            .I(N__11819));
    IoSpan4Mux I__2081 (
            .O(N__11819),
            .I(N__11816));
    Odrv4 I__2080 (
            .O(N__11816),
            .I(port_address_c_0));
    CascadeMux I__2079 (
            .O(N__11813),
            .I(N__11808));
    CascadeMux I__2078 (
            .O(N__11812),
            .I(N__11804));
    CascadeMux I__2077 (
            .O(N__11811),
            .I(N__11801));
    InMux I__2076 (
            .O(N__11808),
            .I(N__11796));
    InMux I__2075 (
            .O(N__11807),
            .I(N__11796));
    InMux I__2074 (
            .O(N__11804),
            .I(N__11791));
    InMux I__2073 (
            .O(N__11801),
            .I(N__11791));
    LocalMux I__2072 (
            .O(N__11796),
            .I(N__11788));
    LocalMux I__2071 (
            .O(N__11791),
            .I(N__11785));
    Span4Mux_v I__2070 (
            .O(N__11788),
            .I(N__11782));
    Span12Mux_h I__2069 (
            .O(N__11785),
            .I(N__11779));
    Sp12to4 I__2068 (
            .O(N__11782),
            .I(N__11776));
    Span12Mux_v I__2067 (
            .O(N__11779),
            .I(N__11773));
    Span12Mux_h I__2066 (
            .O(N__11776),
            .I(N__11770));
    Odrv12 I__2065 (
            .O(N__11773),
            .I(port_address_c_1));
    Odrv12 I__2064 (
            .O(N__11770),
            .I(port_address_c_1));
    InMux I__2063 (
            .O(N__11765),
            .I(N__11758));
    InMux I__2062 (
            .O(N__11764),
            .I(N__11758));
    InMux I__2061 (
            .O(N__11763),
            .I(N__11755));
    LocalMux I__2060 (
            .O(N__11758),
            .I(\this_start_data_delay.this_edge_detector.N_275 ));
    LocalMux I__2059 (
            .O(N__11755),
            .I(\this_start_data_delay.this_edge_detector.N_275 ));
    CascadeMux I__2058 (
            .O(N__11750),
            .I(\this_start_data_delay.this_edge_detector.N_259_cascade_ ));
    InMux I__2057 (
            .O(N__11747),
            .I(N__11744));
    LocalMux I__2056 (
            .O(N__11744),
            .I(N__11741));
    Span4Mux_s2_v I__2055 (
            .O(N__11741),
            .I(N__11738));
    Sp12to4 I__2054 (
            .O(N__11738),
            .I(N__11735));
    Span12Mux_s6_v I__2053 (
            .O(N__11735),
            .I(N__11732));
    Span12Mux_v I__2052 (
            .O(N__11732),
            .I(N__11729));
    Odrv12 I__2051 (
            .O(N__11729),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1 ));
    InMux I__2050 (
            .O(N__11726),
            .I(N__11723));
    LocalMux I__2049 (
            .O(N__11723),
            .I(N__11720));
    Span12Mux_s11_v I__2048 (
            .O(N__11720),
            .I(N__11717));
    Odrv12 I__2047 (
            .O(N__11717),
            .I(\this_vga_signals.mult1_un68_sum_i_1_3 ));
    CascadeMux I__2046 (
            .O(N__11714),
            .I(N__11711));
    InMux I__2045 (
            .O(N__11711),
            .I(N__11708));
    LocalMux I__2044 (
            .O(N__11708),
            .I(N__11705));
    Span4Mux_v I__2043 (
            .O(N__11705),
            .I(N__11702));
    Span4Mux_v I__2042 (
            .O(N__11702),
            .I(N__11695));
    CascadeMux I__2041 (
            .O(N__11701),
            .I(N__11691));
    InMux I__2040 (
            .O(N__11700),
            .I(N__11688));
    InMux I__2039 (
            .O(N__11699),
            .I(N__11685));
    CascadeMux I__2038 (
            .O(N__11698),
            .I(N__11682));
    Span4Mux_v I__2037 (
            .O(N__11695),
            .I(N__11679));
    CascadeMux I__2036 (
            .O(N__11694),
            .I(N__11674));
    InMux I__2035 (
            .O(N__11691),
            .I(N__11671));
    LocalMux I__2034 (
            .O(N__11688),
            .I(N__11668));
    LocalMux I__2033 (
            .O(N__11685),
            .I(N__11665));
    InMux I__2032 (
            .O(N__11682),
            .I(N__11662));
    Span4Mux_v I__2031 (
            .O(N__11679),
            .I(N__11659));
    InMux I__2030 (
            .O(N__11678),
            .I(N__11656));
    InMux I__2029 (
            .O(N__11677),
            .I(N__11651));
    InMux I__2028 (
            .O(N__11674),
            .I(N__11651));
    LocalMux I__2027 (
            .O(N__11671),
            .I(N__11648));
    Span4Mux_h I__2026 (
            .O(N__11668),
            .I(N__11641));
    Span4Mux_h I__2025 (
            .O(N__11665),
            .I(N__11641));
    LocalMux I__2024 (
            .O(N__11662),
            .I(N__11641));
    Odrv4 I__2023 (
            .O(N__11659),
            .I(\this_vga_signals.M_haddress_qZ0Z_4 ));
    LocalMux I__2022 (
            .O(N__11656),
            .I(\this_vga_signals.M_haddress_qZ0Z_4 ));
    LocalMux I__2021 (
            .O(N__11651),
            .I(\this_vga_signals.M_haddress_qZ0Z_4 ));
    Odrv4 I__2020 (
            .O(N__11648),
            .I(\this_vga_signals.M_haddress_qZ0Z_4 ));
    Odrv4 I__2019 (
            .O(N__11641),
            .I(\this_vga_signals.M_haddress_qZ0Z_4 ));
    InMux I__2018 (
            .O(N__11630),
            .I(N__11627));
    LocalMux I__2017 (
            .O(N__11627),
            .I(N__11624));
    Span12Mux_s8_v I__2016 (
            .O(N__11624),
            .I(N__11621));
    Odrv12 I__2015 (
            .O(N__11621),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_2 ));
    CascadeMux I__2014 (
            .O(N__11618),
            .I(N__11615));
    CascadeBuf I__2013 (
            .O(N__11615),
            .I(N__11612));
    CascadeMux I__2012 (
            .O(N__11612),
            .I(N__11609));
    CascadeBuf I__2011 (
            .O(N__11609),
            .I(N__11606));
    CascadeMux I__2010 (
            .O(N__11606),
            .I(N__11603));
    CascadeBuf I__2009 (
            .O(N__11603),
            .I(N__11600));
    CascadeMux I__2008 (
            .O(N__11600),
            .I(N__11597));
    CascadeBuf I__2007 (
            .O(N__11597),
            .I(N__11594));
    CascadeMux I__2006 (
            .O(N__11594),
            .I(N__11591));
    CascadeBuf I__2005 (
            .O(N__11591),
            .I(N__11588));
    CascadeMux I__2004 (
            .O(N__11588),
            .I(N__11585));
    CascadeBuf I__2003 (
            .O(N__11585),
            .I(N__11582));
    CascadeMux I__2002 (
            .O(N__11582),
            .I(N__11579));
    CascadeBuf I__2001 (
            .O(N__11579),
            .I(N__11576));
    CascadeMux I__2000 (
            .O(N__11576),
            .I(N__11573));
    CascadeBuf I__1999 (
            .O(N__11573),
            .I(N__11570));
    CascadeMux I__1998 (
            .O(N__11570),
            .I(N__11567));
    CascadeBuf I__1997 (
            .O(N__11567),
            .I(N__11564));
    CascadeMux I__1996 (
            .O(N__11564),
            .I(N__11561));
    CascadeBuf I__1995 (
            .O(N__11561),
            .I(N__11558));
    CascadeMux I__1994 (
            .O(N__11558),
            .I(N__11555));
    CascadeBuf I__1993 (
            .O(N__11555),
            .I(N__11552));
    CascadeMux I__1992 (
            .O(N__11552),
            .I(N__11549));
    CascadeBuf I__1991 (
            .O(N__11549),
            .I(N__11546));
    CascadeMux I__1990 (
            .O(N__11546),
            .I(N__11543));
    CascadeBuf I__1989 (
            .O(N__11543),
            .I(N__11540));
    CascadeMux I__1988 (
            .O(N__11540),
            .I(N__11537));
    CascadeBuf I__1987 (
            .O(N__11537),
            .I(N__11534));
    CascadeMux I__1986 (
            .O(N__11534),
            .I(N__11531));
    CascadeBuf I__1985 (
            .O(N__11531),
            .I(N__11528));
    CascadeMux I__1984 (
            .O(N__11528),
            .I(N__11525));
    InMux I__1983 (
            .O(N__11525),
            .I(N__11522));
    LocalMux I__1982 (
            .O(N__11522),
            .I(N__11519));
    Odrv12 I__1981 (
            .O(N__11519),
            .I(this_vga_signals_un6_address_if_generate_plus_mult1_un68_sum_i_3));
    CascadeMux I__1980 (
            .O(N__11516),
            .I(N__11513));
    InMux I__1979 (
            .O(N__11513),
            .I(N__11510));
    LocalMux I__1978 (
            .O(N__11510),
            .I(N__11507));
    Span12Mux_h I__1977 (
            .O(N__11507),
            .I(N__11504));
    Odrv12 I__1976 (
            .O(N__11504),
            .I(\this_vga_signals.g0_14_N_8L16_sx ));
    InMux I__1975 (
            .O(N__11501),
            .I(N__11498));
    LocalMux I__1974 (
            .O(N__11498),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_0_0 ));
    CascadeMux I__1973 (
            .O(N__11495),
            .I(N__11489));
    InMux I__1972 (
            .O(N__11494),
            .I(N__11486));
    InMux I__1971 (
            .O(N__11493),
            .I(N__11482));
    InMux I__1970 (
            .O(N__11492),
            .I(N__11479));
    InMux I__1969 (
            .O(N__11489),
            .I(N__11476));
    LocalMux I__1968 (
            .O(N__11486),
            .I(N__11473));
    InMux I__1967 (
            .O(N__11485),
            .I(N__11470));
    LocalMux I__1966 (
            .O(N__11482),
            .I(N__11459));
    LocalMux I__1965 (
            .O(N__11479),
            .I(N__11459));
    LocalMux I__1964 (
            .O(N__11476),
            .I(N__11459));
    Span4Mux_h I__1963 (
            .O(N__11473),
            .I(N__11459));
    LocalMux I__1962 (
            .O(N__11470),
            .I(N__11459));
    Span4Mux_v I__1961 (
            .O(N__11459),
            .I(N__11455));
    CascadeMux I__1960 (
            .O(N__11458),
            .I(N__11452));
    Span4Mux_v I__1959 (
            .O(N__11455),
            .I(N__11449));
    InMux I__1958 (
            .O(N__11452),
            .I(N__11446));
    Sp12to4 I__1957 (
            .O(N__11449),
            .I(N__11441));
    LocalMux I__1956 (
            .O(N__11446),
            .I(N__11441));
    Odrv12 I__1955 (
            .O(N__11441),
            .I(M_this_vram_read_data_3));
    InMux I__1954 (
            .O(N__11438),
            .I(N__11434));
    InMux I__1953 (
            .O(N__11437),
            .I(N__11431));
    LocalMux I__1952 (
            .O(N__11434),
            .I(N__11427));
    LocalMux I__1951 (
            .O(N__11431),
            .I(N__11424));
    InMux I__1950 (
            .O(N__11430),
            .I(N__11421));
    Odrv4 I__1949 (
            .O(N__11427),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    Odrv4 I__1948 (
            .O(N__11424),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    LocalMux I__1947 (
            .O(N__11421),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    InMux I__1946 (
            .O(N__11414),
            .I(N__11410));
    InMux I__1945 (
            .O(N__11413),
            .I(N__11405));
    LocalMux I__1944 (
            .O(N__11410),
            .I(N__11402));
    InMux I__1943 (
            .O(N__11409),
            .I(N__11397));
    InMux I__1942 (
            .O(N__11408),
            .I(N__11397));
    LocalMux I__1941 (
            .O(N__11405),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    Odrv4 I__1940 (
            .O(N__11402),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    LocalMux I__1939 (
            .O(N__11397),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    InMux I__1938 (
            .O(N__11390),
            .I(N__11386));
    InMux I__1937 (
            .O(N__11389),
            .I(N__11383));
    LocalMux I__1936 (
            .O(N__11386),
            .I(\this_start_data_delay.this_edge_detector.N_253_0 ));
    LocalMux I__1935 (
            .O(N__11383),
            .I(\this_start_data_delay.this_edge_detector.N_253_0 ));
    CascadeMux I__1934 (
            .O(N__11378),
            .I(N__11375));
    InMux I__1933 (
            .O(N__11375),
            .I(N__11370));
    InMux I__1932 (
            .O(N__11374),
            .I(N__11367));
    CascadeMux I__1931 (
            .O(N__11373),
            .I(N__11363));
    LocalMux I__1930 (
            .O(N__11370),
            .I(N__11358));
    LocalMux I__1929 (
            .O(N__11367),
            .I(N__11355));
    InMux I__1928 (
            .O(N__11366),
            .I(N__11348));
    InMux I__1927 (
            .O(N__11363),
            .I(N__11348));
    InMux I__1926 (
            .O(N__11362),
            .I(N__11348));
    InMux I__1925 (
            .O(N__11361),
            .I(N__11345));
    Span4Mux_v I__1924 (
            .O(N__11358),
            .I(N__11342));
    Span4Mux_v I__1923 (
            .O(N__11355),
            .I(N__11339));
    LocalMux I__1922 (
            .O(N__11348),
            .I(N__11336));
    LocalMux I__1921 (
            .O(N__11345),
            .I(\this_vga_signals.M_haddress_qZ0Z_3 ));
    Odrv4 I__1920 (
            .O(N__11342),
            .I(\this_vga_signals.M_haddress_qZ0Z_3 ));
    Odrv4 I__1919 (
            .O(N__11339),
            .I(\this_vga_signals.M_haddress_qZ0Z_3 ));
    Odrv4 I__1918 (
            .O(N__11336),
            .I(\this_vga_signals.M_haddress_qZ0Z_3 ));
    CascadeMux I__1917 (
            .O(N__11327),
            .I(\this_start_data_delay.this_edge_detector.N_261_cascade_ ));
    InMux I__1916 (
            .O(N__11324),
            .I(N__11321));
    LocalMux I__1915 (
            .O(N__11321),
            .I(\this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0Z0Z_0 ));
    InMux I__1914 (
            .O(N__11318),
            .I(N__11315));
    LocalMux I__1913 (
            .O(N__11315),
            .I(M_this_start_address_delay_out_0));
    InMux I__1912 (
            .O(N__11312),
            .I(N__11308));
    InMux I__1911 (
            .O(N__11311),
            .I(N__11305));
    LocalMux I__1910 (
            .O(N__11308),
            .I(\this_start_data_delay.this_edge_detector.N_267 ));
    LocalMux I__1909 (
            .O(N__11305),
            .I(\this_start_data_delay.this_edge_detector.N_267 ));
    CascadeMux I__1908 (
            .O(N__11300),
            .I(\this_start_data_delay.this_edge_detector.N_275_cascade_ ));
    CascadeMux I__1907 (
            .O(N__11297),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_ ));
    CascadeMux I__1906 (
            .O(N__11294),
            .I(N__11291));
    InMux I__1905 (
            .O(N__11291),
            .I(N__11288));
    LocalMux I__1904 (
            .O(N__11288),
            .I(N__11285));
    Odrv4 I__1903 (
            .O(N__11285),
            .I(\this_vga_signals.g0_0_0_0 ));
    CascadeMux I__1902 (
            .O(N__11282),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_cascade_ ));
    InMux I__1901 (
            .O(N__11279),
            .I(N__11272));
    InMux I__1900 (
            .O(N__11278),
            .I(N__11272));
    InMux I__1899 (
            .O(N__11277),
            .I(N__11269));
    LocalMux I__1898 (
            .O(N__11272),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_0 ));
    LocalMux I__1897 (
            .O(N__11269),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_0 ));
    InMux I__1896 (
            .O(N__11264),
            .I(N__11261));
    LocalMux I__1895 (
            .O(N__11261),
            .I(N__11258));
    Odrv12 I__1894 (
            .O(N__11258),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0 ));
    CascadeMux I__1893 (
            .O(N__11255),
            .I(\this_vga_signals.g0_0_5_1_cascade_ ));
    CascadeMux I__1892 (
            .O(N__11252),
            .I(N__11249));
    InMux I__1891 (
            .O(N__11249),
            .I(N__11246));
    LocalMux I__1890 (
            .O(N__11246),
            .I(\this_vga_signals.g0_3_1 ));
    CascadeMux I__1889 (
            .O(N__11243),
            .I(\this_vga_signals.if_N_2_1_0_cascade_ ));
    InMux I__1888 (
            .O(N__11240),
            .I(N__11236));
    InMux I__1887 (
            .O(N__11239),
            .I(N__11233));
    LocalMux I__1886 (
            .O(N__11236),
            .I(N__11230));
    LocalMux I__1885 (
            .O(N__11233),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0_0_1_1 ));
    Odrv12 I__1884 (
            .O(N__11230),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0_0_1_1 ));
    CascadeMux I__1883 (
            .O(N__11225),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d_cascade_ ));
    CascadeMux I__1882 (
            .O(N__11222),
            .I(\this_vga_signals.if_N_2_1_1_cascade_ ));
    CascadeMux I__1881 (
            .O(N__11219),
            .I(\this_vga_signals.mult1_un54_sum_c3_2_cascade_ ));
    InMux I__1880 (
            .O(N__11216),
            .I(N__11213));
    LocalMux I__1879 (
            .O(N__11213),
            .I(\this_vga_signals.N_3_1_0 ));
    InMux I__1878 (
            .O(N__11210),
            .I(N__11207));
    LocalMux I__1877 (
            .O(N__11207),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_x ));
    CascadeMux I__1876 (
            .O(N__11204),
            .I(\this_vga_signals.g0_3_0_cascade_ ));
    InMux I__1875 (
            .O(N__11201),
            .I(N__11198));
    LocalMux I__1874 (
            .O(N__11198),
            .I(\this_vga_signals.if_N_2_5 ));
    InMux I__1873 (
            .O(N__11195),
            .I(N__11188));
    InMux I__1872 (
            .O(N__11194),
            .I(N__11188));
    InMux I__1871 (
            .O(N__11193),
            .I(N__11185));
    LocalMux I__1870 (
            .O(N__11188),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    LocalMux I__1869 (
            .O(N__11185),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    InMux I__1868 (
            .O(N__11180),
            .I(N__11177));
    LocalMux I__1867 (
            .O(N__11177),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_18 ));
    CascadeMux I__1866 (
            .O(N__11174),
            .I(\this_start_data_delay.this_edge_detector.N_267_cascade_ ));
    InMux I__1865 (
            .O(N__11171),
            .I(N__11168));
    LocalMux I__1864 (
            .O(N__11168),
            .I(N__11165));
    Span12Mux_s3_v I__1863 (
            .O(N__11165),
            .I(N__11162));
    Span12Mux_v I__1862 (
            .O(N__11162),
            .I(N__11159));
    Odrv12 I__1861 (
            .O(N__11159),
            .I(\this_vga_signals.if_m12_bm ));
    InMux I__1860 (
            .O(N__11156),
            .I(N__11153));
    LocalMux I__1859 (
            .O(N__11153),
            .I(N__11150));
    Span4Mux_v I__1858 (
            .O(N__11150),
            .I(N__11147));
    Span4Mux_v I__1857 (
            .O(N__11147),
            .I(N__11144));
    Span4Mux_v I__1856 (
            .O(N__11144),
            .I(N__11141));
    Span4Mux_v I__1855 (
            .O(N__11141),
            .I(N__11138));
    Odrv4 I__1854 (
            .O(N__11138),
            .I(\this_vga_signals.if_m12_am ));
    InMux I__1853 (
            .O(N__11135),
            .I(N__11132));
    LocalMux I__1852 (
            .O(N__11132),
            .I(N__11129));
    Span12Mux_s5_v I__1851 (
            .O(N__11129),
            .I(N__11126));
    Span12Mux_v I__1850 (
            .O(N__11126),
            .I(N__11123));
    Odrv12 I__1849 (
            .O(N__11123),
            .I(\this_vga_signals.if_m13_ns_1 ));
    CascadeMux I__1848 (
            .O(N__11120),
            .I(N__11117));
    CascadeBuf I__1847 (
            .O(N__11117),
            .I(N__11114));
    CascadeMux I__1846 (
            .O(N__11114),
            .I(N__11111));
    CascadeBuf I__1845 (
            .O(N__11111),
            .I(N__11108));
    CascadeMux I__1844 (
            .O(N__11108),
            .I(N__11105));
    CascadeBuf I__1843 (
            .O(N__11105),
            .I(N__11102));
    CascadeMux I__1842 (
            .O(N__11102),
            .I(N__11099));
    CascadeBuf I__1841 (
            .O(N__11099),
            .I(N__11096));
    CascadeMux I__1840 (
            .O(N__11096),
            .I(N__11093));
    CascadeBuf I__1839 (
            .O(N__11093),
            .I(N__11090));
    CascadeMux I__1838 (
            .O(N__11090),
            .I(N__11087));
    CascadeBuf I__1837 (
            .O(N__11087),
            .I(N__11084));
    CascadeMux I__1836 (
            .O(N__11084),
            .I(N__11081));
    CascadeBuf I__1835 (
            .O(N__11081),
            .I(N__11078));
    CascadeMux I__1834 (
            .O(N__11078),
            .I(N__11075));
    CascadeBuf I__1833 (
            .O(N__11075),
            .I(N__11072));
    CascadeMux I__1832 (
            .O(N__11072),
            .I(N__11069));
    CascadeBuf I__1831 (
            .O(N__11069),
            .I(N__11066));
    CascadeMux I__1830 (
            .O(N__11066),
            .I(N__11063));
    CascadeBuf I__1829 (
            .O(N__11063),
            .I(N__11060));
    CascadeMux I__1828 (
            .O(N__11060),
            .I(N__11057));
    CascadeBuf I__1827 (
            .O(N__11057),
            .I(N__11054));
    CascadeMux I__1826 (
            .O(N__11054),
            .I(N__11051));
    CascadeBuf I__1825 (
            .O(N__11051),
            .I(N__11048));
    CascadeMux I__1824 (
            .O(N__11048),
            .I(N__11045));
    CascadeBuf I__1823 (
            .O(N__11045),
            .I(N__11042));
    CascadeMux I__1822 (
            .O(N__11042),
            .I(N__11039));
    CascadeBuf I__1821 (
            .O(N__11039),
            .I(N__11036));
    CascadeMux I__1820 (
            .O(N__11036),
            .I(N__11033));
    CascadeBuf I__1819 (
            .O(N__11033),
            .I(N__11030));
    CascadeMux I__1818 (
            .O(N__11030),
            .I(N__11027));
    InMux I__1817 (
            .O(N__11027),
            .I(N__11024));
    LocalMux I__1816 (
            .O(N__11024),
            .I(N__11021));
    Odrv12 I__1815 (
            .O(N__11021),
            .I(if_m13_ns));
    CascadeMux I__1814 (
            .O(N__11018),
            .I(\this_vga_signals.N_9_0_0_cascade_ ));
    InMux I__1813 (
            .O(N__11015),
            .I(N__11012));
    LocalMux I__1812 (
            .O(N__11012),
            .I(N__11009));
    Span4Mux_v I__1811 (
            .O(N__11009),
            .I(N__11006));
    Odrv4 I__1810 (
            .O(N__11006),
            .I(\this_vga_signals.g0_4_2 ));
    InMux I__1809 (
            .O(N__11003),
            .I(N__11000));
    LocalMux I__1808 (
            .O(N__11000),
            .I(\this_vga_signals.mult1_un40_sum_1_ac0_2 ));
    InMux I__1807 (
            .O(N__10997),
            .I(N__10994));
    LocalMux I__1806 (
            .O(N__10994),
            .I(N__10991));
    Span4Mux_h I__1805 (
            .O(N__10991),
            .I(N__10988));
    Odrv4 I__1804 (
            .O(N__10988),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_15 ));
    InMux I__1803 (
            .O(N__10985),
            .I(N__10982));
    LocalMux I__1802 (
            .O(N__10982),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_18 ));
    InMux I__1801 (
            .O(N__10979),
            .I(N__10976));
    LocalMux I__1800 (
            .O(N__10976),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_16 ));
    InMux I__1799 (
            .O(N__10973),
            .I(N__10970));
    LocalMux I__1798 (
            .O(N__10970),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_17 ));
    InMux I__1797 (
            .O(N__10967),
            .I(N__10964));
    LocalMux I__1796 (
            .O(N__10964),
            .I(M_state_qZ0Z_5));
    CascadeMux I__1795 (
            .O(N__10961),
            .I(N__10958));
    InMux I__1794 (
            .O(N__10958),
            .I(N__10955));
    LocalMux I__1793 (
            .O(N__10955),
            .I(\this_start_data_delay.this_edge_detector.N_252_0 ));
    InMux I__1792 (
            .O(N__10952),
            .I(N__10949));
    LocalMux I__1791 (
            .O(N__10949),
            .I(N__10946));
    Odrv4 I__1790 (
            .O(N__10946),
            .I(\this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0 ));
    CascadeMux I__1789 (
            .O(N__10943),
            .I(\this_start_data_delay.this_edge_detector.N_252_0_cascade_ ));
    InMux I__1788 (
            .O(N__10940),
            .I(N__10936));
    InMux I__1787 (
            .O(N__10939),
            .I(N__10933));
    LocalMux I__1786 (
            .O(N__10936),
            .I(\this_vga_signals.mult1_un40_sum_1_axb1 ));
    LocalMux I__1785 (
            .O(N__10933),
            .I(\this_vga_signals.mult1_un40_sum_1_axb1 ));
    InMux I__1784 (
            .O(N__10928),
            .I(N__10924));
    InMux I__1783 (
            .O(N__10927),
            .I(N__10921));
    LocalMux I__1782 (
            .O(N__10924),
            .I(\this_vga_signals.mult1_un40_sum_1_c2_0 ));
    LocalMux I__1781 (
            .O(N__10921),
            .I(\this_vga_signals.mult1_un40_sum_1_c2_0 ));
    CascadeMux I__1780 (
            .O(N__10916),
            .I(N__10913));
    InMux I__1779 (
            .O(N__10913),
            .I(N__10907));
    InMux I__1778 (
            .O(N__10912),
            .I(N__10907));
    LocalMux I__1777 (
            .O(N__10907),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc2_0 ));
    CascadeMux I__1776 (
            .O(N__10904),
            .I(\this_vga_signals.N_2_1_1_cascade_ ));
    CascadeMux I__1775 (
            .O(N__10901),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_a4_cascade_ ));
    CascadeMux I__1774 (
            .O(N__10898),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_cascade_ ));
    InMux I__1773 (
            .O(N__10895),
            .I(N__10892));
    LocalMux I__1772 (
            .O(N__10892),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_0 ));
    InMux I__1771 (
            .O(N__10889),
            .I(N__10886));
    LocalMux I__1770 (
            .O(N__10886),
            .I(\this_vga_signals.mult1_un40_sum1_0_3 ));
    InMux I__1769 (
            .O(N__10883),
            .I(N__10875));
    InMux I__1768 (
            .O(N__10882),
            .I(N__10868));
    InMux I__1767 (
            .O(N__10881),
            .I(N__10868));
    InMux I__1766 (
            .O(N__10880),
            .I(N__10863));
    CascadeMux I__1765 (
            .O(N__10879),
            .I(N__10855));
    InMux I__1764 (
            .O(N__10878),
            .I(N__10851));
    LocalMux I__1763 (
            .O(N__10875),
            .I(N__10848));
    InMux I__1762 (
            .O(N__10874),
            .I(N__10843));
    InMux I__1761 (
            .O(N__10873),
            .I(N__10843));
    LocalMux I__1760 (
            .O(N__10868),
            .I(N__10840));
    InMux I__1759 (
            .O(N__10867),
            .I(N__10835));
    InMux I__1758 (
            .O(N__10866),
            .I(N__10835));
    LocalMux I__1757 (
            .O(N__10863),
            .I(N__10832));
    InMux I__1756 (
            .O(N__10862),
            .I(N__10829));
    InMux I__1755 (
            .O(N__10861),
            .I(N__10824));
    InMux I__1754 (
            .O(N__10860),
            .I(N__10824));
    InMux I__1753 (
            .O(N__10859),
            .I(N__10815));
    InMux I__1752 (
            .O(N__10858),
            .I(N__10815));
    InMux I__1751 (
            .O(N__10855),
            .I(N__10815));
    InMux I__1750 (
            .O(N__10854),
            .I(N__10815));
    LocalMux I__1749 (
            .O(N__10851),
            .I(\this_vga_signals.M_haddress_qZ0Z_7 ));
    Odrv12 I__1748 (
            .O(N__10848),
            .I(\this_vga_signals.M_haddress_qZ0Z_7 ));
    LocalMux I__1747 (
            .O(N__10843),
            .I(\this_vga_signals.M_haddress_qZ0Z_7 ));
    Odrv4 I__1746 (
            .O(N__10840),
            .I(\this_vga_signals.M_haddress_qZ0Z_7 ));
    LocalMux I__1745 (
            .O(N__10835),
            .I(\this_vga_signals.M_haddress_qZ0Z_7 ));
    Odrv4 I__1744 (
            .O(N__10832),
            .I(\this_vga_signals.M_haddress_qZ0Z_7 ));
    LocalMux I__1743 (
            .O(N__10829),
            .I(\this_vga_signals.M_haddress_qZ0Z_7 ));
    LocalMux I__1742 (
            .O(N__10824),
            .I(\this_vga_signals.M_haddress_qZ0Z_7 ));
    LocalMux I__1741 (
            .O(N__10815),
            .I(\this_vga_signals.M_haddress_qZ0Z_7 ));
    InMux I__1740 (
            .O(N__10796),
            .I(N__10793));
    LocalMux I__1739 (
            .O(N__10793),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_a5 ));
    InMux I__1738 (
            .O(N__10790),
            .I(N__10787));
    LocalMux I__1737 (
            .O(N__10787),
            .I(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_1 ));
    CascadeMux I__1736 (
            .O(N__10784),
            .I(\this_vga_signals.g1_0_1_cascade_ ));
    InMux I__1735 (
            .O(N__10781),
            .I(N__10778));
    LocalMux I__1734 (
            .O(N__10778),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_1 ));
    InMux I__1733 (
            .O(N__10775),
            .I(N__10772));
    LocalMux I__1732 (
            .O(N__10772),
            .I(\this_vga_signals.g0_0_0_2 ));
    CascadeMux I__1731 (
            .O(N__10769),
            .I(N__10766));
    InMux I__1730 (
            .O(N__10766),
            .I(N__10763));
    LocalMux I__1729 (
            .O(N__10763),
            .I(\this_vga_signals.g0_29_1 ));
    InMux I__1728 (
            .O(N__10760),
            .I(N__10757));
    LocalMux I__1727 (
            .O(N__10757),
            .I(\this_vga_signals.N_3_0_0_0 ));
    InMux I__1726 (
            .O(N__10754),
            .I(N__10751));
    LocalMux I__1725 (
            .O(N__10751),
            .I(N__10748));
    Odrv4 I__1724 (
            .O(N__10748),
            .I(\this_vga_signals.if_N_7 ));
    InMux I__1723 (
            .O(N__10745),
            .I(N__10735));
    InMux I__1722 (
            .O(N__10744),
            .I(N__10735));
    InMux I__1721 (
            .O(N__10743),
            .I(N__10735));
    InMux I__1720 (
            .O(N__10742),
            .I(N__10729));
    LocalMux I__1719 (
            .O(N__10735),
            .I(N__10726));
    InMux I__1718 (
            .O(N__10734),
            .I(N__10723));
    InMux I__1717 (
            .O(N__10733),
            .I(N__10720));
    InMux I__1716 (
            .O(N__10732),
            .I(N__10717));
    LocalMux I__1715 (
            .O(N__10729),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    Odrv4 I__1714 (
            .O(N__10726),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__1713 (
            .O(N__10723),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__1712 (
            .O(N__10720),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__1711 (
            .O(N__10717),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    InMux I__1710 (
            .O(N__10706),
            .I(N__10703));
    LocalMux I__1709 (
            .O(N__10703),
            .I(N__10698));
    InMux I__1708 (
            .O(N__10702),
            .I(N__10695));
    InMux I__1707 (
            .O(N__10701),
            .I(N__10692));
    Odrv4 I__1706 (
            .O(N__10698),
            .I(\this_vga_signals.mult1_un40_sum_m_2 ));
    LocalMux I__1705 (
            .O(N__10695),
            .I(\this_vga_signals.mult1_un40_sum_m_2 ));
    LocalMux I__1704 (
            .O(N__10692),
            .I(\this_vga_signals.mult1_un40_sum_m_2 ));
    CascadeMux I__1703 (
            .O(N__10685),
            .I(N__10682));
    CascadeBuf I__1702 (
            .O(N__10682),
            .I(N__10679));
    CascadeMux I__1701 (
            .O(N__10679),
            .I(N__10676));
    CascadeBuf I__1700 (
            .O(N__10676),
            .I(N__10673));
    CascadeMux I__1699 (
            .O(N__10673),
            .I(N__10670));
    CascadeBuf I__1698 (
            .O(N__10670),
            .I(N__10667));
    CascadeMux I__1697 (
            .O(N__10667),
            .I(N__10664));
    CascadeBuf I__1696 (
            .O(N__10664),
            .I(N__10661));
    CascadeMux I__1695 (
            .O(N__10661),
            .I(N__10658));
    CascadeBuf I__1694 (
            .O(N__10658),
            .I(N__10655));
    CascadeMux I__1693 (
            .O(N__10655),
            .I(N__10652));
    CascadeBuf I__1692 (
            .O(N__10652),
            .I(N__10649));
    CascadeMux I__1691 (
            .O(N__10649),
            .I(N__10646));
    CascadeBuf I__1690 (
            .O(N__10646),
            .I(N__10643));
    CascadeMux I__1689 (
            .O(N__10643),
            .I(N__10640));
    CascadeBuf I__1688 (
            .O(N__10640),
            .I(N__10637));
    CascadeMux I__1687 (
            .O(N__10637),
            .I(N__10634));
    CascadeBuf I__1686 (
            .O(N__10634),
            .I(N__10631));
    CascadeMux I__1685 (
            .O(N__10631),
            .I(N__10628));
    CascadeBuf I__1684 (
            .O(N__10628),
            .I(N__10625));
    CascadeMux I__1683 (
            .O(N__10625),
            .I(N__10622));
    CascadeBuf I__1682 (
            .O(N__10622),
            .I(N__10619));
    CascadeMux I__1681 (
            .O(N__10619),
            .I(N__10616));
    CascadeBuf I__1680 (
            .O(N__10616),
            .I(N__10613));
    CascadeMux I__1679 (
            .O(N__10613),
            .I(N__10610));
    CascadeBuf I__1678 (
            .O(N__10610),
            .I(N__10607));
    CascadeMux I__1677 (
            .O(N__10607),
            .I(N__10604));
    CascadeBuf I__1676 (
            .O(N__10604),
            .I(N__10601));
    CascadeMux I__1675 (
            .O(N__10601),
            .I(N__10598));
    CascadeBuf I__1674 (
            .O(N__10598),
            .I(N__10595));
    CascadeMux I__1673 (
            .O(N__10595),
            .I(N__10592));
    InMux I__1672 (
            .O(N__10592),
            .I(N__10589));
    LocalMux I__1671 (
            .O(N__10589),
            .I(N__10586));
    Span4Mux_v I__1670 (
            .O(N__10586),
            .I(N__10583));
    Span4Mux_v I__1669 (
            .O(N__10583),
            .I(N__10580));
    Sp12to4 I__1668 (
            .O(N__10580),
            .I(N__10572));
    InMux I__1667 (
            .O(N__10579),
            .I(N__10569));
    InMux I__1666 (
            .O(N__10578),
            .I(N__10564));
    InMux I__1665 (
            .O(N__10577),
            .I(N__10564));
    InMux I__1664 (
            .O(N__10576),
            .I(N__10559));
    InMux I__1663 (
            .O(N__10575),
            .I(N__10559));
    Span12Mux_h I__1662 (
            .O(N__10572),
            .I(N__10556));
    LocalMux I__1661 (
            .O(N__10569),
            .I(this_vga_signals_un6_address_if_N_5_mux_0));
    LocalMux I__1660 (
            .O(N__10564),
            .I(this_vga_signals_un6_address_if_N_5_mux_0));
    LocalMux I__1659 (
            .O(N__10559),
            .I(this_vga_signals_un6_address_if_N_5_mux_0));
    Odrv12 I__1658 (
            .O(N__10556),
            .I(this_vga_signals_un6_address_if_N_5_mux_0));
    InMux I__1657 (
            .O(N__10547),
            .I(N__10539));
    InMux I__1656 (
            .O(N__10546),
            .I(N__10539));
    InMux I__1655 (
            .O(N__10545),
            .I(N__10534));
    InMux I__1654 (
            .O(N__10544),
            .I(N__10534));
    LocalMux I__1653 (
            .O(N__10539),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0 ));
    LocalMux I__1652 (
            .O(N__10534),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0 ));
    CascadeMux I__1651 (
            .O(N__10529),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_cascade_ ));
    InMux I__1650 (
            .O(N__10526),
            .I(N__10519));
    InMux I__1649 (
            .O(N__10525),
            .I(N__10516));
    InMux I__1648 (
            .O(N__10524),
            .I(N__10509));
    InMux I__1647 (
            .O(N__10523),
            .I(N__10509));
    InMux I__1646 (
            .O(N__10522),
            .I(N__10509));
    LocalMux I__1645 (
            .O(N__10519),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1644 (
            .O(N__10516),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1643 (
            .O(N__10509),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    CascadeMux I__1642 (
            .O(N__10502),
            .I(N__10499));
    CascadeBuf I__1641 (
            .O(N__10499),
            .I(N__10496));
    CascadeMux I__1640 (
            .O(N__10496),
            .I(N__10493));
    CascadeBuf I__1639 (
            .O(N__10493),
            .I(N__10490));
    CascadeMux I__1638 (
            .O(N__10490),
            .I(N__10487));
    CascadeBuf I__1637 (
            .O(N__10487),
            .I(N__10484));
    CascadeMux I__1636 (
            .O(N__10484),
            .I(N__10481));
    CascadeBuf I__1635 (
            .O(N__10481),
            .I(N__10478));
    CascadeMux I__1634 (
            .O(N__10478),
            .I(N__10475));
    CascadeBuf I__1633 (
            .O(N__10475),
            .I(N__10472));
    CascadeMux I__1632 (
            .O(N__10472),
            .I(N__10469));
    CascadeBuf I__1631 (
            .O(N__10469),
            .I(N__10466));
    CascadeMux I__1630 (
            .O(N__10466),
            .I(N__10463));
    CascadeBuf I__1629 (
            .O(N__10463),
            .I(N__10460));
    CascadeMux I__1628 (
            .O(N__10460),
            .I(N__10457));
    CascadeBuf I__1627 (
            .O(N__10457),
            .I(N__10454));
    CascadeMux I__1626 (
            .O(N__10454),
            .I(N__10451));
    CascadeBuf I__1625 (
            .O(N__10451),
            .I(N__10448));
    CascadeMux I__1624 (
            .O(N__10448),
            .I(N__10445));
    CascadeBuf I__1623 (
            .O(N__10445),
            .I(N__10442));
    CascadeMux I__1622 (
            .O(N__10442),
            .I(N__10439));
    CascadeBuf I__1621 (
            .O(N__10439),
            .I(N__10436));
    CascadeMux I__1620 (
            .O(N__10436),
            .I(N__10433));
    CascadeBuf I__1619 (
            .O(N__10433),
            .I(N__10430));
    CascadeMux I__1618 (
            .O(N__10430),
            .I(N__10427));
    CascadeBuf I__1617 (
            .O(N__10427),
            .I(N__10424));
    CascadeMux I__1616 (
            .O(N__10424),
            .I(N__10421));
    CascadeBuf I__1615 (
            .O(N__10421),
            .I(N__10418));
    CascadeMux I__1614 (
            .O(N__10418),
            .I(N__10415));
    CascadeBuf I__1613 (
            .O(N__10415),
            .I(N__10412));
    CascadeMux I__1612 (
            .O(N__10412),
            .I(N__10409));
    InMux I__1611 (
            .O(N__10409),
            .I(N__10406));
    LocalMux I__1610 (
            .O(N__10406),
            .I(N__10403));
    Span4Mux_h I__1609 (
            .O(N__10403),
            .I(N__10400));
    Span4Mux_h I__1608 (
            .O(N__10400),
            .I(N__10397));
    Sp12to4 I__1607 (
            .O(N__10397),
            .I(N__10394));
    Span12Mux_v I__1606 (
            .O(N__10394),
            .I(N__10391));
    Odrv12 I__1605 (
            .O(N__10391),
            .I(this_vga_signals_un6_address_if_generate_plus_mult1_un47_sum_i_3));
    CascadeMux I__1604 (
            .O(N__10388),
            .I(N__10384));
    InMux I__1603 (
            .O(N__10387),
            .I(N__10378));
    InMux I__1602 (
            .O(N__10384),
            .I(N__10378));
    InMux I__1601 (
            .O(N__10383),
            .I(N__10375));
    LocalMux I__1600 (
            .O(N__10378),
            .I(\this_vga_signals.mult1_un40_sum_m_1 ));
    LocalMux I__1599 (
            .O(N__10375),
            .I(\this_vga_signals.mult1_un40_sum_m_1 ));
    InMux I__1598 (
            .O(N__10370),
            .I(N__10360));
    InMux I__1597 (
            .O(N__10369),
            .I(N__10360));
    InMux I__1596 (
            .O(N__10368),
            .I(N__10360));
    InMux I__1595 (
            .O(N__10367),
            .I(N__10357));
    LocalMux I__1594 (
            .O(N__10360),
            .I(\this_vga_signals.CO1_1_0 ));
    LocalMux I__1593 (
            .O(N__10357),
            .I(\this_vga_signals.CO1_1_0 ));
    CascadeMux I__1592 (
            .O(N__10352),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ));
    InMux I__1591 (
            .O(N__10349),
            .I(N__10346));
    LocalMux I__1590 (
            .O(N__10346),
            .I(\this_vga_signals.if_m1 ));
    InMux I__1589 (
            .O(N__10343),
            .I(N__10339));
    InMux I__1588 (
            .O(N__10342),
            .I(N__10336));
    LocalMux I__1587 (
            .O(N__10339),
            .I(\this_vga_signals.mult1_un54_sum_axb1_2 ));
    LocalMux I__1586 (
            .O(N__10336),
            .I(\this_vga_signals.mult1_un54_sum_axb1_2 ));
    InMux I__1585 (
            .O(N__10331),
            .I(N__10328));
    LocalMux I__1584 (
            .O(N__10328),
            .I(\this_vga_signals.g1_N_2L1 ));
    CascadeMux I__1583 (
            .O(N__10325),
            .I(N__10322));
    InMux I__1582 (
            .O(N__10322),
            .I(N__10319));
    LocalMux I__1581 (
            .O(N__10319),
            .I(\this_vga_signals.G_5_0_x2_1 ));
    CascadeMux I__1580 (
            .O(N__10316),
            .I(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ));
    CascadeMux I__1579 (
            .O(N__10313),
            .I(\this_vga_signals.g2_4_cascade_ ));
    CascadeMux I__1578 (
            .O(N__10310),
            .I(N__10307));
    InMux I__1577 (
            .O(N__10307),
            .I(N__10304));
    LocalMux I__1576 (
            .O(N__10304),
            .I(\this_vga_signals.if_m1_3 ));
    CascadeMux I__1575 (
            .O(N__10301),
            .I(\this_vga_signals.if_m1_3_cascade_ ));
    CascadeMux I__1574 (
            .O(N__10298),
            .I(\this_vga_signals.if_m8_am_cascade_ ));
    InMux I__1573 (
            .O(N__10295),
            .I(N__10292));
    LocalMux I__1572 (
            .O(N__10292),
            .I(\this_vga_signals.if_m8_bm ));
    InMux I__1571 (
            .O(N__10289),
            .I(N__10286));
    LocalMux I__1570 (
            .O(N__10286),
            .I(\this_vga_signals.g1_0_0 ));
    CascadeMux I__1569 (
            .O(N__10283),
            .I(\this_vga_signals.g0_0_2_cascade_ ));
    InMux I__1568 (
            .O(N__10280),
            .I(N__10277));
    LocalMux I__1567 (
            .O(N__10277),
            .I(\this_vga_signals.g0_0_3_0 ));
    InMux I__1566 (
            .O(N__10274),
            .I(N__10271));
    LocalMux I__1565 (
            .O(N__10271),
            .I(N__10268));
    Odrv4 I__1564 (
            .O(N__10268),
            .I(\this_vga_signals.g3_2 ));
    InMux I__1563 (
            .O(N__10265),
            .I(N__10262));
    LocalMux I__1562 (
            .O(N__10262),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_0_0_1 ));
    InMux I__1561 (
            .O(N__10259),
            .I(\this_vga_signals.un1_M_haddress_q_cry_9 ));
    InMux I__1560 (
            .O(N__10256),
            .I(\this_vga_signals.un1_M_haddress_q_cry_10 ));
    SRMux I__1559 (
            .O(N__10253),
            .I(N__10249));
    SRMux I__1558 (
            .O(N__10252),
            .I(N__10246));
    LocalMux I__1557 (
            .O(N__10249),
            .I(N__10243));
    LocalMux I__1556 (
            .O(N__10246),
            .I(N__10240));
    Span4Mux_h I__1555 (
            .O(N__10243),
            .I(N__10237));
    Span4Mux_h I__1554 (
            .O(N__10240),
            .I(N__10234));
    Span4Mux_h I__1553 (
            .O(N__10237),
            .I(N__10231));
    Odrv4 I__1552 (
            .O(N__10234),
            .I(\this_vga_signals.M_hstate_q_RNIFIH84Z0Z_5 ));
    Odrv4 I__1551 (
            .O(N__10231),
            .I(\this_vga_signals.M_hstate_q_RNIFIH84Z0Z_5 ));
    InMux I__1550 (
            .O(N__10226),
            .I(N__10223));
    LocalMux I__1549 (
            .O(N__10223),
            .I(N__10220));
    Span4Mux_h I__1548 (
            .O(N__10220),
            .I(N__10217));
    Odrv4 I__1547 (
            .O(N__10217),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_16 ));
    InMux I__1546 (
            .O(N__10214),
            .I(N__10211));
    LocalMux I__1545 (
            .O(N__10211),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_17 ));
    InMux I__1544 (
            .O(N__10208),
            .I(N__10205));
    LocalMux I__1543 (
            .O(N__10205),
            .I(N__10199));
    InMux I__1542 (
            .O(N__10204),
            .I(N__10196));
    InMux I__1541 (
            .O(N__10203),
            .I(N__10193));
    InMux I__1540 (
            .O(N__10202),
            .I(N__10190));
    Odrv12 I__1539 (
            .O(N__10199),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    LocalMux I__1538 (
            .O(N__10196),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    LocalMux I__1537 (
            .O(N__10193),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    LocalMux I__1536 (
            .O(N__10190),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    InMux I__1535 (
            .O(N__10181),
            .I(N__10178));
    LocalMux I__1534 (
            .O(N__10178),
            .I(N__10171));
    InMux I__1533 (
            .O(N__10177),
            .I(N__10166));
    InMux I__1532 (
            .O(N__10176),
            .I(N__10166));
    InMux I__1531 (
            .O(N__10175),
            .I(N__10163));
    InMux I__1530 (
            .O(N__10174),
            .I(N__10160));
    Odrv12 I__1529 (
            .O(N__10171),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0_i ));
    LocalMux I__1528 (
            .O(N__10166),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0_i ));
    LocalMux I__1527 (
            .O(N__10163),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0_i ));
    LocalMux I__1526 (
            .O(N__10160),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0_i ));
    CascadeMux I__1525 (
            .O(N__10151),
            .I(N__10148));
    CascadeBuf I__1524 (
            .O(N__10148),
            .I(N__10145));
    CascadeMux I__1523 (
            .O(N__10145),
            .I(N__10142));
    CascadeBuf I__1522 (
            .O(N__10142),
            .I(N__10139));
    CascadeMux I__1521 (
            .O(N__10139),
            .I(N__10136));
    CascadeBuf I__1520 (
            .O(N__10136),
            .I(N__10133));
    CascadeMux I__1519 (
            .O(N__10133),
            .I(N__10130));
    CascadeBuf I__1518 (
            .O(N__10130),
            .I(N__10127));
    CascadeMux I__1517 (
            .O(N__10127),
            .I(N__10124));
    CascadeBuf I__1516 (
            .O(N__10124),
            .I(N__10121));
    CascadeMux I__1515 (
            .O(N__10121),
            .I(N__10118));
    CascadeBuf I__1514 (
            .O(N__10118),
            .I(N__10115));
    CascadeMux I__1513 (
            .O(N__10115),
            .I(N__10112));
    CascadeBuf I__1512 (
            .O(N__10112),
            .I(N__10109));
    CascadeMux I__1511 (
            .O(N__10109),
            .I(N__10106));
    CascadeBuf I__1510 (
            .O(N__10106),
            .I(N__10103));
    CascadeMux I__1509 (
            .O(N__10103),
            .I(N__10100));
    CascadeBuf I__1508 (
            .O(N__10100),
            .I(N__10097));
    CascadeMux I__1507 (
            .O(N__10097),
            .I(N__10094));
    CascadeBuf I__1506 (
            .O(N__10094),
            .I(N__10091));
    CascadeMux I__1505 (
            .O(N__10091),
            .I(N__10088));
    CascadeBuf I__1504 (
            .O(N__10088),
            .I(N__10085));
    CascadeMux I__1503 (
            .O(N__10085),
            .I(N__10082));
    CascadeBuf I__1502 (
            .O(N__10082),
            .I(N__10079));
    CascadeMux I__1501 (
            .O(N__10079),
            .I(N__10076));
    CascadeBuf I__1500 (
            .O(N__10076),
            .I(N__10073));
    CascadeMux I__1499 (
            .O(N__10073),
            .I(N__10070));
    CascadeBuf I__1498 (
            .O(N__10070),
            .I(N__10067));
    CascadeMux I__1497 (
            .O(N__10067),
            .I(N__10064));
    CascadeBuf I__1496 (
            .O(N__10064),
            .I(N__10061));
    CascadeMux I__1495 (
            .O(N__10061),
            .I(N__10058));
    InMux I__1494 (
            .O(N__10058),
            .I(N__10055));
    LocalMux I__1493 (
            .O(N__10055),
            .I(N__10052));
    Sp12to4 I__1492 (
            .O(N__10052),
            .I(N__10049));
    Span12Mux_h I__1491 (
            .O(N__10049),
            .I(N__10046));
    Span12Mux_v I__1490 (
            .O(N__10046),
            .I(N__10043));
    Odrv12 I__1489 (
            .O(N__10043),
            .I(this_vga_signals_un6_address_if_generate_plus_mult1_un54_sum_i_3));
    CascadeMux I__1488 (
            .O(N__10040),
            .I(\this_vga_signals.g1_3_1_cascade_ ));
    CascadeMux I__1487 (
            .O(N__10037),
            .I(\this_vga_signals.if_N_7_cascade_ ));
    InMux I__1486 (
            .O(N__10034),
            .I(\this_vga_signals.un1_M_haddress_q_cry_0 ));
    InMux I__1485 (
            .O(N__10031),
            .I(N__10027));
    InMux I__1484 (
            .O(N__10030),
            .I(N__10024));
    LocalMux I__1483 (
            .O(N__10027),
            .I(N__10021));
    LocalMux I__1482 (
            .O(N__10024),
            .I(\this_vga_signals.M_haddress_qZ0Z_2 ));
    Odrv4 I__1481 (
            .O(N__10021),
            .I(\this_vga_signals.M_haddress_qZ0Z_2 ));
    InMux I__1480 (
            .O(N__10016),
            .I(\this_vga_signals.un1_M_haddress_q_cry_1 ));
    InMux I__1479 (
            .O(N__10013),
            .I(\this_vga_signals.un1_M_haddress_q_cry_2 ));
    InMux I__1478 (
            .O(N__10010),
            .I(\this_vga_signals.un1_M_haddress_q_cry_3 ));
    InMux I__1477 (
            .O(N__10007),
            .I(N__10002));
    CascadeMux I__1476 (
            .O(N__10006),
            .I(N__9996));
    CascadeMux I__1475 (
            .O(N__10005),
            .I(N__9992));
    LocalMux I__1474 (
            .O(N__10002),
            .I(N__9988));
    InMux I__1473 (
            .O(N__10001),
            .I(N__9985));
    CascadeMux I__1472 (
            .O(N__10000),
            .I(N__9981));
    InMux I__1471 (
            .O(N__9999),
            .I(N__9978));
    InMux I__1470 (
            .O(N__9996),
            .I(N__9975));
    InMux I__1469 (
            .O(N__9995),
            .I(N__9968));
    InMux I__1468 (
            .O(N__9992),
            .I(N__9968));
    InMux I__1467 (
            .O(N__9991),
            .I(N__9968));
    Span4Mux_h I__1466 (
            .O(N__9988),
            .I(N__9965));
    LocalMux I__1465 (
            .O(N__9985),
            .I(N__9962));
    InMux I__1464 (
            .O(N__9984),
            .I(N__9957));
    InMux I__1463 (
            .O(N__9981),
            .I(N__9957));
    LocalMux I__1462 (
            .O(N__9978),
            .I(\this_vga_signals.M_haddress_qZ0Z_5 ));
    LocalMux I__1461 (
            .O(N__9975),
            .I(\this_vga_signals.M_haddress_qZ0Z_5 ));
    LocalMux I__1460 (
            .O(N__9968),
            .I(\this_vga_signals.M_haddress_qZ0Z_5 ));
    Odrv4 I__1459 (
            .O(N__9965),
            .I(\this_vga_signals.M_haddress_qZ0Z_5 ));
    Odrv4 I__1458 (
            .O(N__9962),
            .I(\this_vga_signals.M_haddress_qZ0Z_5 ));
    LocalMux I__1457 (
            .O(N__9957),
            .I(\this_vga_signals.M_haddress_qZ0Z_5 ));
    InMux I__1456 (
            .O(N__9944),
            .I(\this_vga_signals.un1_M_haddress_q_cry_4 ));
    CascadeMux I__1455 (
            .O(N__9941),
            .I(N__9937));
    CascadeMux I__1454 (
            .O(N__9940),
            .I(N__9934));
    InMux I__1453 (
            .O(N__9937),
            .I(N__9925));
    InMux I__1452 (
            .O(N__9934),
            .I(N__9925));
    InMux I__1451 (
            .O(N__9933),
            .I(N__9925));
    InMux I__1450 (
            .O(N__9932),
            .I(N__9917));
    LocalMux I__1449 (
            .O(N__9925),
            .I(N__9914));
    InMux I__1448 (
            .O(N__9924),
            .I(N__9911));
    InMux I__1447 (
            .O(N__9923),
            .I(N__9908));
    InMux I__1446 (
            .O(N__9922),
            .I(N__9901));
    InMux I__1445 (
            .O(N__9921),
            .I(N__9901));
    InMux I__1444 (
            .O(N__9920),
            .I(N__9901));
    LocalMux I__1443 (
            .O(N__9917),
            .I(\this_vga_signals.M_haddress_qZ0Z_6 ));
    Odrv4 I__1442 (
            .O(N__9914),
            .I(\this_vga_signals.M_haddress_qZ0Z_6 ));
    LocalMux I__1441 (
            .O(N__9911),
            .I(\this_vga_signals.M_haddress_qZ0Z_6 ));
    LocalMux I__1440 (
            .O(N__9908),
            .I(\this_vga_signals.M_haddress_qZ0Z_6 ));
    LocalMux I__1439 (
            .O(N__9901),
            .I(\this_vga_signals.M_haddress_qZ0Z_6 ));
    InMux I__1438 (
            .O(N__9890),
            .I(\this_vga_signals.un1_M_haddress_q_cry_5 ));
    InMux I__1437 (
            .O(N__9887),
            .I(\this_vga_signals.un1_M_haddress_q_cry_6 ));
    InMux I__1436 (
            .O(N__9884),
            .I(bfn_18_16_0_));
    InMux I__1435 (
            .O(N__9881),
            .I(\this_vga_signals.un1_M_haddress_q_cry_8 ));
    InMux I__1434 (
            .O(N__9878),
            .I(N__9875));
    LocalMux I__1433 (
            .O(N__9875),
            .I(N__9871));
    InMux I__1432 (
            .O(N__9874),
            .I(N__9868));
    Odrv4 I__1431 (
            .O(N__9871),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_3_1 ));
    LocalMux I__1430 (
            .O(N__9868),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_3_1 ));
    CascadeMux I__1429 (
            .O(N__9863),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_1_0_cascade_ ));
    InMux I__1428 (
            .O(N__9860),
            .I(N__9857));
    LocalMux I__1427 (
            .O(N__9857),
            .I(\this_vga_signals.if_N_4_i ));
    CascadeMux I__1426 (
            .O(N__9854),
            .I(this_vga_signals_un6_address_if_N_5_mux_0_cascade_));
    CascadeMux I__1425 (
            .O(N__9851),
            .I(\this_vga_signals.mult1_un47_sum_c3_cascade_ ));
    InMux I__1424 (
            .O(N__9848),
            .I(N__9845));
    LocalMux I__1423 (
            .O(N__9845),
            .I(\this_vga_signals.if_m1_1 ));
    CascadeMux I__1422 (
            .O(N__9842),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_ ));
    InMux I__1421 (
            .O(N__9839),
            .I(N__9836));
    LocalMux I__1420 (
            .O(N__9836),
            .I(\this_vga_signals.if_m1_9_1 ));
    InMux I__1419 (
            .O(N__9833),
            .I(N__9828));
    InMux I__1418 (
            .O(N__9832),
            .I(N__9825));
    CascadeMux I__1417 (
            .O(N__9831),
            .I(N__9820));
    LocalMux I__1416 (
            .O(N__9828),
            .I(N__9817));
    LocalMux I__1415 (
            .O(N__9825),
            .I(N__9813));
    CascadeMux I__1414 (
            .O(N__9824),
            .I(N__9810));
    InMux I__1413 (
            .O(N__9823),
            .I(N__9807));
    InMux I__1412 (
            .O(N__9820),
            .I(N__9804));
    Sp12to4 I__1411 (
            .O(N__9817),
            .I(N__9801));
    CascadeMux I__1410 (
            .O(N__9816),
            .I(N__9798));
    Span4Mux_v I__1409 (
            .O(N__9813),
            .I(N__9795));
    InMux I__1408 (
            .O(N__9810),
            .I(N__9792));
    LocalMux I__1407 (
            .O(N__9807),
            .I(N__9787));
    LocalMux I__1406 (
            .O(N__9804),
            .I(N__9787));
    Span12Mux_v I__1405 (
            .O(N__9801),
            .I(N__9784));
    InMux I__1404 (
            .O(N__9798),
            .I(N__9781));
    Span4Mux_h I__1403 (
            .O(N__9795),
            .I(N__9774));
    LocalMux I__1402 (
            .O(N__9792),
            .I(N__9774));
    Span4Mux_h I__1401 (
            .O(N__9787),
            .I(N__9774));
    Odrv12 I__1400 (
            .O(N__9784),
            .I(\this_vga_signals.M_hstate_qZ0Z_1 ));
    LocalMux I__1399 (
            .O(N__9781),
            .I(\this_vga_signals.M_hstate_qZ0Z_1 ));
    Odrv4 I__1398 (
            .O(N__9774),
            .I(\this_vga_signals.M_hstate_qZ0Z_1 ));
    InMux I__1397 (
            .O(N__9767),
            .I(N__9764));
    LocalMux I__1396 (
            .O(N__9764),
            .I(\this_vga_signals.M_haddress_qZ0Z_0 ));
    InMux I__1395 (
            .O(N__9761),
            .I(N__9758));
    LocalMux I__1394 (
            .O(N__9758),
            .I(\this_vga_signals.M_haddress_qZ0Z_1 ));
    InMux I__1393 (
            .O(N__9755),
            .I(N__9752));
    LocalMux I__1392 (
            .O(N__9752),
            .I(\this_vga_signals.if_m2_0_1 ));
    InMux I__1391 (
            .O(N__9749),
            .I(N__9746));
    LocalMux I__1390 (
            .O(N__9746),
            .I(\this_vga_signals.if_N_3_0_i ));
    CascadeMux I__1389 (
            .O(N__9743),
            .I(\this_vga_signals.if_N_3_0_i_cascade_ ));
    InMux I__1388 (
            .O(N__9740),
            .I(N__9737));
    LocalMux I__1387 (
            .O(N__9737),
            .I(\this_vga_signals.mult1_un75_sum_c3_0 ));
    InMux I__1386 (
            .O(N__9734),
            .I(N__9731));
    LocalMux I__1385 (
            .O(N__9731),
            .I(\this_vga_signals.if_i1_mux_0 ));
    InMux I__1384 (
            .O(N__9728),
            .I(N__9725));
    LocalMux I__1383 (
            .O(N__9725),
            .I(\this_vga_signals.if_m2 ));
    CascadeMux I__1382 (
            .O(N__9722),
            .I(\this_vga_signals.M_haddress_q_RNILVKM8Z0Z_6_cascade_ ));
    CascadeMux I__1381 (
            .O(N__9719),
            .I(\this_vga_signals.mult1_un54_sum_c3_cascade_ ));
    InMux I__1380 (
            .O(N__9716),
            .I(N__9713));
    LocalMux I__1379 (
            .O(N__9713),
            .I(\this_vga_signals.if_N_8_i ));
    InMux I__1378 (
            .O(N__9710),
            .I(N__9707));
    LocalMux I__1377 (
            .O(N__9707),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_1_0 ));
    InMux I__1376 (
            .O(N__9704),
            .I(N__9701));
    LocalMux I__1375 (
            .O(N__9701),
            .I(N__9698));
    Odrv4 I__1374 (
            .O(N__9698),
            .I(\this_vga_signals.g1_2_1 ));
    CascadeMux I__1373 (
            .O(N__9695),
            .I(N__9692));
    InMux I__1372 (
            .O(N__9692),
            .I(N__9689));
    LocalMux I__1371 (
            .O(N__9689),
            .I(N__9686));
    Odrv4 I__1370 (
            .O(N__9686),
            .I(\this_vga_signals.g2_5_0 ));
    InMux I__1369 (
            .O(N__9683),
            .I(N__9680));
    LocalMux I__1368 (
            .O(N__9680),
            .I(\this_vga_signals.M_vaddress_q_RNI85LKP4Z0Z_2 ));
    CascadeMux I__1367 (
            .O(N__9677),
            .I(\this_vga_signals.mult1_un54_sum_axb1_1_0_cascade_ ));
    CascadeMux I__1366 (
            .O(N__9674),
            .I(\this_vga_signals.mult1_un61_sum_c3_1_1_0_cascade_ ));
    CascadeMux I__1365 (
            .O(N__9671),
            .I(\this_vga_signals.g3_0_0_0_1_cascade_ ));
    InMux I__1364 (
            .O(N__9668),
            .I(N__9665));
    LocalMux I__1363 (
            .O(N__9665),
            .I(\this_vga_signals.g1_2 ));
    InMux I__1362 (
            .O(N__9662),
            .I(N__9659));
    LocalMux I__1361 (
            .O(N__9659),
            .I(\this_vga_signals.g2 ));
    InMux I__1360 (
            .O(N__9656),
            .I(N__9653));
    LocalMux I__1359 (
            .O(N__9653),
            .I(\this_vga_signals.g1_0_1_0_0 ));
    InMux I__1358 (
            .O(N__9650),
            .I(N__9647));
    LocalMux I__1357 (
            .O(N__9647),
            .I(\this_vga_signals.N_4_i ));
    InMux I__1356 (
            .O(N__9644),
            .I(N__9641));
    LocalMux I__1355 (
            .O(N__9641),
            .I(\this_vga_signals.g0_14_N_7L14_1 ));
    CascadeMux I__1354 (
            .O(N__9638),
            .I(\this_vga_signals.g2_3_0_cascade_ ));
    CascadeMux I__1353 (
            .O(N__9635),
            .I(\this_vga_signals.if_N_2_4_cascade_ ));
    CascadeMux I__1352 (
            .O(N__9632),
            .I(\this_vga_signals.mult1_un61_sum_c3_2_cascade_ ));
    CascadeMux I__1351 (
            .O(N__9629),
            .I(\this_vga_signals.g0_0_6_cascade_ ));
    InMux I__1350 (
            .O(N__9626),
            .I(N__9623));
    LocalMux I__1349 (
            .O(N__9623),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    InMux I__1348 (
            .O(N__9620),
            .I(N__9617));
    LocalMux I__1347 (
            .O(N__9617),
            .I(\this_vga_signals.g0_1_0 ));
    CascadeMux I__1346 (
            .O(N__9614),
            .I(\this_vga_signals.mult1_un61_sum_c3_cascade_ ));
    InMux I__1345 (
            .O(N__9611),
            .I(N__9608));
    LocalMux I__1344 (
            .O(N__9608),
            .I(\this_vga_signals.mult1_un68_sum_axb2_i ));
    CascadeMux I__1343 (
            .O(N__9605),
            .I(N__9602));
    InMux I__1342 (
            .O(N__9602),
            .I(N__9599));
    LocalMux I__1341 (
            .O(N__9599),
            .I(\this_vga_signals.g0_14_N_4L6 ));
    InMux I__1340 (
            .O(N__9596),
            .I(N__9591));
    InMux I__1339 (
            .O(N__9595),
            .I(N__9588));
    InMux I__1338 (
            .O(N__9594),
            .I(N__9585));
    LocalMux I__1337 (
            .O(N__9591),
            .I(N__9582));
    LocalMux I__1336 (
            .O(N__9588),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1335 (
            .O(N__9585),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__1334 (
            .O(N__9582),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__1333 (
            .O(N__9575),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__1332 (
            .O(N__9572),
            .I(N__9567));
    InMux I__1331 (
            .O(N__9571),
            .I(N__9564));
    InMux I__1330 (
            .O(N__9570),
            .I(N__9561));
    LocalMux I__1329 (
            .O(N__9567),
            .I(N__9558));
    LocalMux I__1328 (
            .O(N__9564),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1327 (
            .O(N__9561),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__1326 (
            .O(N__9558),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    InMux I__1325 (
            .O(N__9551),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__1324 (
            .O(N__9548),
            .I(N__9542));
    InMux I__1323 (
            .O(N__9547),
            .I(N__9537));
    InMux I__1322 (
            .O(N__9546),
            .I(N__9537));
    InMux I__1321 (
            .O(N__9545),
            .I(N__9534));
    LocalMux I__1320 (
            .O(N__9542),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1319 (
            .O(N__9537),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1318 (
            .O(N__9534),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    InMux I__1317 (
            .O(N__9527),
            .I(bfn_17_18_0_));
    InMux I__1316 (
            .O(N__9524),
            .I(N__9517));
    InMux I__1315 (
            .O(N__9523),
            .I(N__9512));
    InMux I__1314 (
            .O(N__9522),
            .I(N__9512));
    InMux I__1313 (
            .O(N__9521),
            .I(N__9507));
    InMux I__1312 (
            .O(N__9520),
            .I(N__9507));
    LocalMux I__1311 (
            .O(N__9517),
            .I(N__9499));
    LocalMux I__1310 (
            .O(N__9512),
            .I(N__9499));
    LocalMux I__1309 (
            .O(N__9507),
            .I(N__9499));
    InMux I__1308 (
            .O(N__9506),
            .I(N__9496));
    Span4Mux_v I__1307 (
            .O(N__9499),
            .I(N__9493));
    LocalMux I__1306 (
            .O(N__9496),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    Odrv4 I__1305 (
            .O(N__9493),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    InMux I__1304 (
            .O(N__9488),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_9 ));
    InMux I__1303 (
            .O(N__9485),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_10 ));
    InMux I__1302 (
            .O(N__9482),
            .I(N__9477));
    InMux I__1301 (
            .O(N__9481),
            .I(N__9472));
    InMux I__1300 (
            .O(N__9480),
            .I(N__9472));
    LocalMux I__1299 (
            .O(N__9477),
            .I(\this_vga_signals.M_hcounter_qZ0Z_11 ));
    LocalMux I__1298 (
            .O(N__9472),
            .I(\this_vga_signals.M_hcounter_qZ0Z_11 ));
    InMux I__1297 (
            .O(N__9467),
            .I(N__9464));
    LocalMux I__1296 (
            .O(N__9464),
            .I(\this_vga_signals.g1_1_1 ));
    CascadeMux I__1295 (
            .O(N__9461),
            .I(\this_vga_signals.g2_1_0_cascade_ ));
    CascadeMux I__1294 (
            .O(N__9458),
            .I(\this_vga_signals.mult1_un40_sum_0_ac0_3_0_a1_0_cascade_ ));
    InMux I__1293 (
            .O(N__9455),
            .I(N__9452));
    LocalMux I__1292 (
            .O(N__9452),
            .I(\this_vga_signals.if_m3_0_0 ));
    InMux I__1291 (
            .O(N__9449),
            .I(N__9446));
    LocalMux I__1290 (
            .O(N__9446),
            .I(\this_vga_signals.mult1_un40_sum_0_ac0_3_1 ));
    CascadeMux I__1289 (
            .O(N__9443),
            .I(\this_vga_signals.mult1_un40_sum_0_ac0_3_0_cascade_ ));
    InMux I__1288 (
            .O(N__9440),
            .I(N__9437));
    LocalMux I__1287 (
            .O(N__9437),
            .I(\this_vga_signals.mult1_un40_sum_0_ac0_3_2 ));
    InMux I__1286 (
            .O(N__9434),
            .I(N__9431));
    LocalMux I__1285 (
            .O(N__9431),
            .I(N__9428));
    Odrv4 I__1284 (
            .O(N__9428),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_14 ));
    InMux I__1283 (
            .O(N__9425),
            .I(N__9422));
    LocalMux I__1282 (
            .O(N__9422),
            .I(N__9419));
    Span4Mux_v I__1281 (
            .O(N__9419),
            .I(N__9416));
    Odrv4 I__1280 (
            .O(N__9416),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_15 ));
    InMux I__1279 (
            .O(N__9413),
            .I(N__9404));
    InMux I__1278 (
            .O(N__9412),
            .I(N__9404));
    InMux I__1277 (
            .O(N__9411),
            .I(N__9401));
    InMux I__1276 (
            .O(N__9410),
            .I(N__9396));
    InMux I__1275 (
            .O(N__9409),
            .I(N__9396));
    LocalMux I__1274 (
            .O(N__9404),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1273 (
            .O(N__9401),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1272 (
            .O(N__9396),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    CascadeMux I__1271 (
            .O(N__9389),
            .I(N__9386));
    InMux I__1270 (
            .O(N__9386),
            .I(N__9382));
    InMux I__1269 (
            .O(N__9385),
            .I(N__9378));
    LocalMux I__1268 (
            .O(N__9382),
            .I(N__9375));
    InMux I__1267 (
            .O(N__9381),
            .I(N__9372));
    LocalMux I__1266 (
            .O(N__9378),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__1265 (
            .O(N__9375),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__1264 (
            .O(N__9372),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    InMux I__1263 (
            .O(N__9365),
            .I(N__9361));
    InMux I__1262 (
            .O(N__9364),
            .I(N__9358));
    LocalMux I__1261 (
            .O(N__9361),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__1260 (
            .O(N__9358),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__1259 (
            .O(N__9353),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__1258 (
            .O(N__9350),
            .I(N__9346));
    InMux I__1257 (
            .O(N__9349),
            .I(N__9343));
    LocalMux I__1256 (
            .O(N__9346),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1255 (
            .O(N__9343),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__1254 (
            .O(N__9338),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    CascadeMux I__1253 (
            .O(N__9335),
            .I(N__9331));
    InMux I__1252 (
            .O(N__9334),
            .I(N__9328));
    InMux I__1251 (
            .O(N__9331),
            .I(N__9325));
    LocalMux I__1250 (
            .O(N__9328),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1249 (
            .O(N__9325),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__1248 (
            .O(N__9320),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__1247 (
            .O(N__9317),
            .I(N__9312));
    InMux I__1246 (
            .O(N__9316),
            .I(N__9309));
    InMux I__1245 (
            .O(N__9315),
            .I(N__9306));
    LocalMux I__1244 (
            .O(N__9312),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1243 (
            .O(N__9309),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1242 (
            .O(N__9306),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    InMux I__1241 (
            .O(N__9299),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__1240 (
            .O(N__9296),
            .I(N__9290));
    InMux I__1239 (
            .O(N__9295),
            .I(N__9283));
    InMux I__1238 (
            .O(N__9294),
            .I(N__9283));
    InMux I__1237 (
            .O(N__9293),
            .I(N__9283));
    LocalMux I__1236 (
            .O(N__9290),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1235 (
            .O(N__9283),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    InMux I__1234 (
            .O(N__9278),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__1233 (
            .O(N__9275),
            .I(N__9272));
    LocalMux I__1232 (
            .O(N__9272),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_13 ));
    CascadeMux I__1231 (
            .O(N__9269),
            .I(\this_vga_signals.mult1_un40_sum_0_ac0_3_2_1_cascade_ ));
    CascadeMux I__1230 (
            .O(N__9266),
            .I(\this_vga_signals.if_N_2_6_cascade_ ));
    InMux I__1229 (
            .O(N__9263),
            .I(N__9260));
    LocalMux I__1228 (
            .O(N__9260),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    InMux I__1227 (
            .O(N__9257),
            .I(N__9254));
    LocalMux I__1226 (
            .O(N__9254),
            .I(\this_vga_signals.g0_14_N_7L14 ));
    CascadeMux I__1225 (
            .O(N__9251),
            .I(\this_vga_signals.if_N_9_0_cascade_ ));
    InMux I__1224 (
            .O(N__9248),
            .I(N__9245));
    LocalMux I__1223 (
            .O(N__9245),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    CascadeMux I__1222 (
            .O(N__9242),
            .I(\this_vga_signals.mult1_un61_sum_axb1_cascade_ ));
    CascadeMux I__1221 (
            .O(N__9239),
            .I(\this_vga_signals.if_m3_1_2_cascade_ ));
    InMux I__1220 (
            .O(N__9236),
            .I(N__9233));
    LocalMux I__1219 (
            .O(N__9233),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_out ));
    InMux I__1218 (
            .O(N__9230),
            .I(N__9227));
    LocalMux I__1217 (
            .O(N__9227),
            .I(\this_vga_signals.if_i2_mux_0 ));
    CascadeMux I__1216 (
            .O(N__9224),
            .I(\this_vga_signals.if_N_6_0_0_cascade_ ));
    CascadeMux I__1215 (
            .O(N__9221),
            .I(N__9218));
    CascadeBuf I__1214 (
            .O(N__9218),
            .I(N__9215));
    CascadeMux I__1213 (
            .O(N__9215),
            .I(N__9212));
    CascadeBuf I__1212 (
            .O(N__9212),
            .I(N__9209));
    CascadeMux I__1211 (
            .O(N__9209),
            .I(N__9206));
    CascadeBuf I__1210 (
            .O(N__9206),
            .I(N__9203));
    CascadeMux I__1209 (
            .O(N__9203),
            .I(N__9200));
    CascadeBuf I__1208 (
            .O(N__9200),
            .I(N__9197));
    CascadeMux I__1207 (
            .O(N__9197),
            .I(N__9194));
    CascadeBuf I__1206 (
            .O(N__9194),
            .I(N__9191));
    CascadeMux I__1205 (
            .O(N__9191),
            .I(N__9188));
    CascadeBuf I__1204 (
            .O(N__9188),
            .I(N__9185));
    CascadeMux I__1203 (
            .O(N__9185),
            .I(N__9182));
    CascadeBuf I__1202 (
            .O(N__9182),
            .I(N__9179));
    CascadeMux I__1201 (
            .O(N__9179),
            .I(N__9176));
    CascadeBuf I__1200 (
            .O(N__9176),
            .I(N__9173));
    CascadeMux I__1199 (
            .O(N__9173),
            .I(N__9170));
    CascadeBuf I__1198 (
            .O(N__9170),
            .I(N__9167));
    CascadeMux I__1197 (
            .O(N__9167),
            .I(N__9164));
    CascadeBuf I__1196 (
            .O(N__9164),
            .I(N__9161));
    CascadeMux I__1195 (
            .O(N__9161),
            .I(N__9158));
    CascadeBuf I__1194 (
            .O(N__9158),
            .I(N__9155));
    CascadeMux I__1193 (
            .O(N__9155),
            .I(N__9152));
    CascadeBuf I__1192 (
            .O(N__9152),
            .I(N__9149));
    CascadeMux I__1191 (
            .O(N__9149),
            .I(N__9146));
    CascadeBuf I__1190 (
            .O(N__9146),
            .I(N__9143));
    CascadeMux I__1189 (
            .O(N__9143),
            .I(N__9140));
    CascadeBuf I__1188 (
            .O(N__9140),
            .I(N__9137));
    CascadeMux I__1187 (
            .O(N__9137),
            .I(N__9134));
    CascadeBuf I__1186 (
            .O(N__9134),
            .I(N__9131));
    CascadeMux I__1185 (
            .O(N__9131),
            .I(N__9128));
    InMux I__1184 (
            .O(N__9128),
            .I(N__9125));
    LocalMux I__1183 (
            .O(N__9125),
            .I(N__9122));
    Span12Mux_h I__1182 (
            .O(N__9122),
            .I(N__9119));
    Span12Mux_v I__1181 (
            .O(N__9119),
            .I(N__9116));
    Odrv12 I__1180 (
            .O(N__9116),
            .I(this_vga_signals_un6_address_if_generate_plus_mult1_un75_sum_i_3));
    CascadeMux I__1179 (
            .O(N__9113),
            .I(\this_vga_signals.g2_2_cascade_ ));
    CascadeMux I__1178 (
            .O(N__9110),
            .I(\this_vga_signals.g1_cascade_ ));
    CascadeMux I__1177 (
            .O(N__9107),
            .I(\this_vga_signals.g2_5_cascade_ ));
    InMux I__1176 (
            .O(N__9104),
            .I(N__9101));
    LocalMux I__1175 (
            .O(N__9101),
            .I(\this_vga_signals.g1_1_4 ));
    CascadeMux I__1174 (
            .O(N__9098),
            .I(\this_vga_signals.g0_14_N_8L16_cascade_ ));
    CascadeMux I__1173 (
            .O(N__9095),
            .I(\this_vga_signals.mult1_un75_sum_c3_0_0_cascade_ ));
    CascadeMux I__1172 (
            .O(N__9092),
            .I(N__9089));
    CascadeBuf I__1171 (
            .O(N__9089),
            .I(N__9086));
    CascadeMux I__1170 (
            .O(N__9086),
            .I(N__9083));
    CascadeBuf I__1169 (
            .O(N__9083),
            .I(N__9080));
    CascadeMux I__1168 (
            .O(N__9080),
            .I(N__9077));
    CascadeBuf I__1167 (
            .O(N__9077),
            .I(N__9074));
    CascadeMux I__1166 (
            .O(N__9074),
            .I(N__9071));
    CascadeBuf I__1165 (
            .O(N__9071),
            .I(N__9068));
    CascadeMux I__1164 (
            .O(N__9068),
            .I(N__9065));
    CascadeBuf I__1163 (
            .O(N__9065),
            .I(N__9062));
    CascadeMux I__1162 (
            .O(N__9062),
            .I(N__9059));
    CascadeBuf I__1161 (
            .O(N__9059),
            .I(N__9056));
    CascadeMux I__1160 (
            .O(N__9056),
            .I(N__9053));
    CascadeBuf I__1159 (
            .O(N__9053),
            .I(N__9050));
    CascadeMux I__1158 (
            .O(N__9050),
            .I(N__9047));
    CascadeBuf I__1157 (
            .O(N__9047),
            .I(N__9044));
    CascadeMux I__1156 (
            .O(N__9044),
            .I(N__9041));
    CascadeBuf I__1155 (
            .O(N__9041),
            .I(N__9038));
    CascadeMux I__1154 (
            .O(N__9038),
            .I(N__9035));
    CascadeBuf I__1153 (
            .O(N__9035),
            .I(N__9032));
    CascadeMux I__1152 (
            .O(N__9032),
            .I(N__9029));
    CascadeBuf I__1151 (
            .O(N__9029),
            .I(N__9026));
    CascadeMux I__1150 (
            .O(N__9026),
            .I(N__9023));
    CascadeBuf I__1149 (
            .O(N__9023),
            .I(N__9020));
    CascadeMux I__1148 (
            .O(N__9020),
            .I(N__9017));
    CascadeBuf I__1147 (
            .O(N__9017),
            .I(N__9014));
    CascadeMux I__1146 (
            .O(N__9014),
            .I(N__9011));
    CascadeBuf I__1145 (
            .O(N__9011),
            .I(N__9008));
    CascadeMux I__1144 (
            .O(N__9008),
            .I(N__9005));
    CascadeBuf I__1143 (
            .O(N__9005),
            .I(N__9002));
    CascadeMux I__1142 (
            .O(N__9002),
            .I(N__8999));
    InMux I__1141 (
            .O(N__8999),
            .I(N__8996));
    LocalMux I__1140 (
            .O(N__8996),
            .I(N__8993));
    Span4Mux_v I__1139 (
            .O(N__8993),
            .I(N__8990));
    Span4Mux_h I__1138 (
            .O(N__8990),
            .I(N__8987));
    Span4Mux_h I__1137 (
            .O(N__8987),
            .I(N__8984));
    Sp12to4 I__1136 (
            .O(N__8984),
            .I(N__8981));
    Span12Mux_s11_v I__1135 (
            .O(N__8981),
            .I(N__8978));
    Odrv12 I__1134 (
            .O(N__8978),
            .I(this_vga_signals_un14_address_if_generate_plus_mult1_un75_sum_i_3));
    CascadeMux I__1133 (
            .O(N__8975),
            .I(\this_vga_signals.N_386_0_cascade_ ));
    InMux I__1132 (
            .O(N__8972),
            .I(N__8968));
    InMux I__1131 (
            .O(N__8971),
            .I(N__8965));
    LocalMux I__1130 (
            .O(N__8968),
            .I(N__8960));
    LocalMux I__1129 (
            .O(N__8965),
            .I(N__8960));
    Odrv4 I__1128 (
            .O(N__8960),
            .I(\this_vga_signals.M_hstate_q_srsts_0_o3_2_1 ));
    InMux I__1127 (
            .O(N__8957),
            .I(N__8952));
    InMux I__1126 (
            .O(N__8956),
            .I(N__8949));
    InMux I__1125 (
            .O(N__8955),
            .I(N__8946));
    LocalMux I__1124 (
            .O(N__8952),
            .I(\this_vga_signals.N_388_0 ));
    LocalMux I__1123 (
            .O(N__8949),
            .I(\this_vga_signals.N_388_0 ));
    LocalMux I__1122 (
            .O(N__8946),
            .I(\this_vga_signals.N_388_0 ));
    CascadeMux I__1121 (
            .O(N__8939),
            .I(N__8936));
    InMux I__1120 (
            .O(N__8936),
            .I(N__8933));
    LocalMux I__1119 (
            .O(N__8933),
            .I(\this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5 ));
    InMux I__1118 (
            .O(N__8930),
            .I(N__8925));
    InMux I__1117 (
            .O(N__8929),
            .I(N__8920));
    InMux I__1116 (
            .O(N__8928),
            .I(N__8920));
    LocalMux I__1115 (
            .O(N__8925),
            .I(\this_vga_signals.N_393_0 ));
    LocalMux I__1114 (
            .O(N__8920),
            .I(\this_vga_signals.N_393_0 ));
    InMux I__1113 (
            .O(N__8915),
            .I(N__8912));
    LocalMux I__1112 (
            .O(N__8912),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    InMux I__1111 (
            .O(N__8909),
            .I(N__8897));
    InMux I__1110 (
            .O(N__8908),
            .I(N__8897));
    InMux I__1109 (
            .O(N__8907),
            .I(N__8897));
    InMux I__1108 (
            .O(N__8906),
            .I(N__8897));
    LocalMux I__1107 (
            .O(N__8897),
            .I(N__8894));
    Odrv12 I__1106 (
            .O(N__8894),
            .I(rst_n_c));
    InMux I__1105 (
            .O(N__8891),
            .I(N__8888));
    LocalMux I__1104 (
            .O(N__8888),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__1103 (
            .O(N__8885),
            .I(N__8882));
    LocalMux I__1102 (
            .O(N__8882),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    CascadeMux I__1101 (
            .O(N__8879),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa_cascade_ ));
    InMux I__1100 (
            .O(N__8876),
            .I(N__8873));
    LocalMux I__1099 (
            .O(N__8873),
            .I(\this_vga_signals.N_405_0 ));
    InMux I__1098 (
            .O(N__8870),
            .I(N__8864));
    InMux I__1097 (
            .O(N__8869),
            .I(N__8864));
    LocalMux I__1096 (
            .O(N__8864),
            .I(\this_vga_signals.M_hstate_qZ0Z_0 ));
    CascadeMux I__1095 (
            .O(N__8861),
            .I(\this_vga_signals.N_405_0_cascade_ ));
    InMux I__1094 (
            .O(N__8858),
            .I(N__8855));
    LocalMux I__1093 (
            .O(N__8855),
            .I(\this_vga_signals.N_409 ));
    InMux I__1092 (
            .O(N__8852),
            .I(N__8847));
    InMux I__1091 (
            .O(N__8851),
            .I(N__8842));
    InMux I__1090 (
            .O(N__8850),
            .I(N__8842));
    LocalMux I__1089 (
            .O(N__8847),
            .I(\this_vga_signals.N_397_0 ));
    LocalMux I__1088 (
            .O(N__8842),
            .I(\this_vga_signals.N_397_0 ));
    InMux I__1087 (
            .O(N__8837),
            .I(N__8832));
    InMux I__1086 (
            .O(N__8836),
            .I(N__8829));
    InMux I__1085 (
            .O(N__8835),
            .I(N__8826));
    LocalMux I__1084 (
            .O(N__8832),
            .I(\this_vga_signals.M_hstate_qZ0Z_5 ));
    LocalMux I__1083 (
            .O(N__8829),
            .I(\this_vga_signals.M_hstate_qZ0Z_5 ));
    LocalMux I__1082 (
            .O(N__8826),
            .I(\this_vga_signals.M_hstate_qZ0Z_5 ));
    CascadeMux I__1081 (
            .O(N__8819),
            .I(\this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5_cascade_ ));
    InMux I__1080 (
            .O(N__8816),
            .I(N__8810));
    InMux I__1079 (
            .O(N__8815),
            .I(N__8810));
    LocalMux I__1078 (
            .O(N__8810),
            .I(\this_vga_signals.N_385_0 ));
    CascadeMux I__1077 (
            .O(N__8807),
            .I(\this_vga_signals.N_385_0_cascade_ ));
    InMux I__1076 (
            .O(N__8804),
            .I(N__8801));
    LocalMux I__1075 (
            .O(N__8801),
            .I(N__8795));
    InMux I__1074 (
            .O(N__8800),
            .I(N__8792));
    InMux I__1073 (
            .O(N__8799),
            .I(N__8787));
    InMux I__1072 (
            .O(N__8798),
            .I(N__8787));
    Odrv4 I__1071 (
            .O(N__8795),
            .I(\this_vga_signals.N_391_0 ));
    LocalMux I__1070 (
            .O(N__8792),
            .I(\this_vga_signals.N_391_0 ));
    LocalMux I__1069 (
            .O(N__8787),
            .I(\this_vga_signals.N_391_0 ));
    InMux I__1068 (
            .O(N__8780),
            .I(N__8775));
    CascadeMux I__1067 (
            .O(N__8779),
            .I(N__8771));
    CascadeMux I__1066 (
            .O(N__8778),
            .I(N__8768));
    LocalMux I__1065 (
            .O(N__8775),
            .I(N__8765));
    InMux I__1064 (
            .O(N__8774),
            .I(N__8762));
    InMux I__1063 (
            .O(N__8771),
            .I(N__8759));
    InMux I__1062 (
            .O(N__8768),
            .I(N__8756));
    Odrv4 I__1061 (
            .O(N__8765),
            .I(\this_vga_signals.N_386_0 ));
    LocalMux I__1060 (
            .O(N__8762),
            .I(\this_vga_signals.N_386_0 ));
    LocalMux I__1059 (
            .O(N__8759),
            .I(\this_vga_signals.N_386_0 ));
    LocalMux I__1058 (
            .O(N__8756),
            .I(\this_vga_signals.N_386_0 ));
    CascadeMux I__1057 (
            .O(N__8747),
            .I(\this_vga_signals.N_390_0_cascade_ ));
    InMux I__1056 (
            .O(N__8744),
            .I(N__8738));
    InMux I__1055 (
            .O(N__8743),
            .I(N__8738));
    LocalMux I__1054 (
            .O(N__8738),
            .I(\this_vga_signals.N_390_0 ));
    InMux I__1053 (
            .O(N__8735),
            .I(N__8731));
    InMux I__1052 (
            .O(N__8734),
            .I(N__8728));
    LocalMux I__1051 (
            .O(N__8731),
            .I(\this_vga_signals.M_hstate_qZ0Z_2 ));
    LocalMux I__1050 (
            .O(N__8728),
            .I(\this_vga_signals.M_hstate_qZ0Z_2 ));
    CascadeMux I__1049 (
            .O(N__8723),
            .I(\this_vga_signals.N_413_cascade_ ));
    InMux I__1048 (
            .O(N__8720),
            .I(N__8716));
    InMux I__1047 (
            .O(N__8719),
            .I(N__8713));
    LocalMux I__1046 (
            .O(N__8716),
            .I(\this_vga_signals.N_398_0 ));
    LocalMux I__1045 (
            .O(N__8713),
            .I(\this_vga_signals.N_398_0 ));
    CascadeMux I__1044 (
            .O(N__8708),
            .I(N__8704));
    CascadeMux I__1043 (
            .O(N__8707),
            .I(N__8701));
    InMux I__1042 (
            .O(N__8704),
            .I(N__8696));
    InMux I__1041 (
            .O(N__8701),
            .I(N__8696));
    LocalMux I__1040 (
            .O(N__8696),
            .I(\this_vga_signals.M_hstate_qZ0Z_3 ));
    InMux I__1039 (
            .O(N__8693),
            .I(N__8690));
    LocalMux I__1038 (
            .O(N__8690),
            .I(N__8687));
    Odrv4 I__1037 (
            .O(N__8687),
            .I(\this_vga_signals.M_hstate_q_srsts_0_a3_0_4 ));
    InMux I__1036 (
            .O(N__8684),
            .I(N__8681));
    LocalMux I__1035 (
            .O(N__8681),
            .I(\this_vga_signals.N_416 ));
    CascadeMux I__1034 (
            .O(N__8678),
            .I(\this_vga_signals.M_hstate_q_srsts_0_a3_0_4_cascade_ ));
    InMux I__1033 (
            .O(N__8675),
            .I(N__8672));
    LocalMux I__1032 (
            .O(N__8672),
            .I(N__8669));
    Span4Mux_v I__1031 (
            .O(N__8669),
            .I(N__8666));
    Span4Mux_h I__1030 (
            .O(N__8666),
            .I(N__8663));
    Span4Mux_v I__1029 (
            .O(N__8663),
            .I(N__8659));
    InMux I__1028 (
            .O(N__8662),
            .I(N__8656));
    Odrv4 I__1027 (
            .O(N__8659),
            .I(\this_vga_signals.M_hstate_qZ0Z_4 ));
    LocalMux I__1026 (
            .O(N__8656),
            .I(\this_vga_signals.M_hstate_qZ0Z_4 ));
    InMux I__1025 (
            .O(N__8651),
            .I(N__8648));
    LocalMux I__1024 (
            .O(N__8648),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_12 ));
    InMux I__1023 (
            .O(N__8645),
            .I(N__8642));
    LocalMux I__1022 (
            .O(N__8642),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_11 ));
    InMux I__1021 (
            .O(N__8639),
            .I(N__8636));
    LocalMux I__1020 (
            .O(N__8636),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_8 ));
    InMux I__1019 (
            .O(N__8633),
            .I(N__8630));
    LocalMux I__1018 (
            .O(N__8630),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_9 ));
    InMux I__1017 (
            .O(N__8627),
            .I(N__8624));
    LocalMux I__1016 (
            .O(N__8624),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_14 ));
    CascadeMux I__1015 (
            .O(N__8621),
            .I(\this_vga_signals.N_417_cascade_ ));
    CascadeMux I__1014 (
            .O(N__8618),
            .I(\this_vga_signals.N_412_cascade_ ));
    CascadeMux I__1013 (
            .O(N__8615),
            .I(N__8609));
    InMux I__1012 (
            .O(N__8614),
            .I(N__8606));
    InMux I__1011 (
            .O(N__8613),
            .I(N__8603));
    InMux I__1010 (
            .O(N__8612),
            .I(N__8600));
    InMux I__1009 (
            .O(N__8609),
            .I(N__8597));
    LocalMux I__1008 (
            .O(N__8606),
            .I(N__8592));
    LocalMux I__1007 (
            .O(N__8603),
            .I(N__8592));
    LocalMux I__1006 (
            .O(N__8600),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__1005 (
            .O(N__8597),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__1004 (
            .O(N__8592),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    InMux I__1003 (
            .O(N__8585),
            .I(N__8578));
    InMux I__1002 (
            .O(N__8584),
            .I(N__8573));
    InMux I__1001 (
            .O(N__8583),
            .I(N__8573));
    InMux I__1000 (
            .O(N__8582),
            .I(N__8570));
    InMux I__999 (
            .O(N__8581),
            .I(N__8567));
    LocalMux I__998 (
            .O(N__8578),
            .I(N__8564));
    LocalMux I__997 (
            .O(N__8573),
            .I(N__8559));
    LocalMux I__996 (
            .O(N__8570),
            .I(N__8559));
    LocalMux I__995 (
            .O(N__8567),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__994 (
            .O(N__8564),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__993 (
            .O(N__8559),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    InMux I__992 (
            .O(N__8552),
            .I(N__8548));
    InMux I__991 (
            .O(N__8551),
            .I(N__8545));
    LocalMux I__990 (
            .O(N__8548),
            .I(\this_vga_signals.N_230_0 ));
    LocalMux I__989 (
            .O(N__8545),
            .I(\this_vga_signals.N_230_0 ));
    CascadeMux I__988 (
            .O(N__8540),
            .I(\this_vga_signals.M_vstate_q_srsts_0_o2_2_5_cascade_ ));
    CascadeMux I__987 (
            .O(N__8537),
            .I(N__8531));
    InMux I__986 (
            .O(N__8536),
            .I(N__8527));
    InMux I__985 (
            .O(N__8535),
            .I(N__8524));
    InMux I__984 (
            .O(N__8534),
            .I(N__8517));
    InMux I__983 (
            .O(N__8531),
            .I(N__8517));
    InMux I__982 (
            .O(N__8530),
            .I(N__8517));
    LocalMux I__981 (
            .O(N__8527),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__980 (
            .O(N__8524),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__979 (
            .O(N__8517),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    InMux I__978 (
            .O(N__8510),
            .I(N__8503));
    InMux I__977 (
            .O(N__8509),
            .I(N__8493));
    InMux I__976 (
            .O(N__8508),
            .I(N__8493));
    InMux I__975 (
            .O(N__8507),
            .I(N__8493));
    InMux I__974 (
            .O(N__8506),
            .I(N__8493));
    LocalMux I__973 (
            .O(N__8503),
            .I(N__8490));
    InMux I__972 (
            .O(N__8502),
            .I(N__8487));
    LocalMux I__971 (
            .O(N__8493),
            .I(\this_vga_signals.N_248_0 ));
    Odrv4 I__970 (
            .O(N__8490),
            .I(\this_vga_signals.N_248_0 ));
    LocalMux I__969 (
            .O(N__8487),
            .I(\this_vga_signals.N_248_0 ));
    CascadeMux I__968 (
            .O(N__8480),
            .I(\this_vga_signals.N_248_0_cascade_ ));
    CascadeMux I__967 (
            .O(N__8477),
            .I(N__8473));
    InMux I__966 (
            .O(N__8476),
            .I(N__8467));
    InMux I__965 (
            .O(N__8473),
            .I(N__8464));
    CascadeMux I__964 (
            .O(N__8472),
            .I(N__8461));
    CascadeMux I__963 (
            .O(N__8471),
            .I(N__8458));
    CascadeMux I__962 (
            .O(N__8470),
            .I(N__8455));
    LocalMux I__961 (
            .O(N__8467),
            .I(N__8450));
    LocalMux I__960 (
            .O(N__8464),
            .I(N__8447));
    InMux I__959 (
            .O(N__8461),
            .I(N__8440));
    InMux I__958 (
            .O(N__8458),
            .I(N__8440));
    InMux I__957 (
            .O(N__8455),
            .I(N__8440));
    InMux I__956 (
            .O(N__8454),
            .I(N__8437));
    InMux I__955 (
            .O(N__8453),
            .I(N__8434));
    Odrv4 I__954 (
            .O(N__8450),
            .I(\this_vga_signals.M_vstate_qZ0Z_5 ));
    Odrv4 I__953 (
            .O(N__8447),
            .I(\this_vga_signals.M_vstate_qZ0Z_5 ));
    LocalMux I__952 (
            .O(N__8440),
            .I(\this_vga_signals.M_vstate_qZ0Z_5 ));
    LocalMux I__951 (
            .O(N__8437),
            .I(\this_vga_signals.M_vstate_qZ0Z_5 ));
    LocalMux I__950 (
            .O(N__8434),
            .I(\this_vga_signals.M_vstate_qZ0Z_5 ));
    InMux I__949 (
            .O(N__8423),
            .I(N__8420));
    LocalMux I__948 (
            .O(N__8420),
            .I(\this_vga_signals.N_252 ));
    InMux I__947 (
            .O(N__8417),
            .I(N__8412));
    InMux I__946 (
            .O(N__8416),
            .I(N__8409));
    InMux I__945 (
            .O(N__8415),
            .I(N__8403));
    LocalMux I__944 (
            .O(N__8412),
            .I(N__8398));
    LocalMux I__943 (
            .O(N__8409),
            .I(N__8398));
    InMux I__942 (
            .O(N__8408),
            .I(N__8395));
    InMux I__941 (
            .O(N__8407),
            .I(N__8392));
    InMux I__940 (
            .O(N__8406),
            .I(N__8389));
    LocalMux I__939 (
            .O(N__8403),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__938 (
            .O(N__8398),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__937 (
            .O(N__8395),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__936 (
            .O(N__8392),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__935 (
            .O(N__8389),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    CascadeMux I__934 (
            .O(N__8378),
            .I(N__8373));
    InMux I__933 (
            .O(N__8377),
            .I(N__8368));
    InMux I__932 (
            .O(N__8376),
            .I(N__8365));
    InMux I__931 (
            .O(N__8373),
            .I(N__8362));
    InMux I__930 (
            .O(N__8372),
            .I(N__8359));
    InMux I__929 (
            .O(N__8371),
            .I(N__8356));
    LocalMux I__928 (
            .O(N__8368),
            .I(N__8353));
    LocalMux I__927 (
            .O(N__8365),
            .I(N__8350));
    LocalMux I__926 (
            .O(N__8362),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__925 (
            .O(N__8359),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__924 (
            .O(N__8356),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__923 (
            .O(N__8353),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__922 (
            .O(N__8350),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    CascadeMux I__921 (
            .O(N__8339),
            .I(N__8335));
    CascadeMux I__920 (
            .O(N__8338),
            .I(N__8332));
    InMux I__919 (
            .O(N__8335),
            .I(N__8326));
    InMux I__918 (
            .O(N__8332),
            .I(N__8323));
    InMux I__917 (
            .O(N__8331),
            .I(N__8320));
    InMux I__916 (
            .O(N__8330),
            .I(N__8317));
    InMux I__915 (
            .O(N__8329),
            .I(N__8314));
    LocalMux I__914 (
            .O(N__8326),
            .I(N__8309));
    LocalMux I__913 (
            .O(N__8323),
            .I(N__8309));
    LocalMux I__912 (
            .O(N__8320),
            .I(N__8304));
    LocalMux I__911 (
            .O(N__8317),
            .I(N__8304));
    LocalMux I__910 (
            .O(N__8314),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__909 (
            .O(N__8309),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__908 (
            .O(N__8304),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    InMux I__907 (
            .O(N__8297),
            .I(N__8291));
    InMux I__906 (
            .O(N__8296),
            .I(N__8287));
    InMux I__905 (
            .O(N__8295),
            .I(N__8284));
    InMux I__904 (
            .O(N__8294),
            .I(N__8281));
    LocalMux I__903 (
            .O(N__8291),
            .I(N__8278));
    InMux I__902 (
            .O(N__8290),
            .I(N__8275));
    LocalMux I__901 (
            .O(N__8287),
            .I(N__8272));
    LocalMux I__900 (
            .O(N__8284),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__899 (
            .O(N__8281),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__898 (
            .O(N__8278),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__897 (
            .O(N__8275),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__896 (
            .O(N__8272),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    CascadeMux I__895 (
            .O(N__8261),
            .I(\this_vga_signals.M_vstate_q_srsts_0_o2_2_3_cascade_ ));
    InMux I__894 (
            .O(N__8258),
            .I(N__8255));
    LocalMux I__893 (
            .O(N__8255),
            .I(N__8252));
    Odrv4 I__892 (
            .O(N__8252),
            .I(\this_vga_signals.N_255 ));
    InMux I__891 (
            .O(N__8249),
            .I(N__8246));
    LocalMux I__890 (
            .O(N__8246),
            .I(\this_vga_signals.M_vstate_q_srsts_0_o2_2_3 ));
    CascadeMux I__889 (
            .O(N__8243),
            .I(N__8239));
    InMux I__888 (
            .O(N__8242),
            .I(N__8234));
    InMux I__887 (
            .O(N__8239),
            .I(N__8234));
    LocalMux I__886 (
            .O(N__8234),
            .I(\this_vga_signals.M_vstate_qZ0Z_3 ));
    InMux I__885 (
            .O(N__8231),
            .I(N__8222));
    InMux I__884 (
            .O(N__8230),
            .I(N__8222));
    InMux I__883 (
            .O(N__8229),
            .I(N__8217));
    InMux I__882 (
            .O(N__8228),
            .I(N__8217));
    InMux I__881 (
            .O(N__8227),
            .I(N__8214));
    LocalMux I__880 (
            .O(N__8222),
            .I(\this_vga_signals.N_226_0 ));
    LocalMux I__879 (
            .O(N__8217),
            .I(\this_vga_signals.N_226_0 ));
    LocalMux I__878 (
            .O(N__8214),
            .I(\this_vga_signals.N_226_0 ));
    InMux I__877 (
            .O(N__8207),
            .I(N__8204));
    LocalMux I__876 (
            .O(N__8204),
            .I(\this_vga_signals.N_256 ));
    InMux I__875 (
            .O(N__8201),
            .I(N__8198));
    LocalMux I__874 (
            .O(N__8198),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_7 ));
    InMux I__873 (
            .O(N__8195),
            .I(N__8192));
    LocalMux I__872 (
            .O(N__8192),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_10 ));
    IoInMux I__871 (
            .O(N__8189),
            .I(N__8186));
    LocalMux I__870 (
            .O(N__8186),
            .I(N__8183));
    Span12Mux_s11_h I__869 (
            .O(N__8183),
            .I(N__8180));
    Odrv12 I__868 (
            .O(N__8180),
            .I(\this_vga_signals.M_vstate_q_RNI3M6M4Z0Z_0 ));
    CascadeMux I__867 (
            .O(N__8177),
            .I(\this_vga_signals.N_251_cascade_ ));
    InMux I__866 (
            .O(N__8174),
            .I(N__8170));
    InMux I__865 (
            .O(N__8173),
            .I(N__8167));
    LocalMux I__864 (
            .O(N__8170),
            .I(N__8164));
    LocalMux I__863 (
            .O(N__8167),
            .I(\this_vga_signals.N_237_0 ));
    Odrv4 I__862 (
            .O(N__8164),
            .I(\this_vga_signals.N_237_0 ));
    InMux I__861 (
            .O(N__8159),
            .I(N__8155));
    InMux I__860 (
            .O(N__8158),
            .I(N__8151));
    LocalMux I__859 (
            .O(N__8155),
            .I(N__8148));
    InMux I__858 (
            .O(N__8154),
            .I(N__8145));
    LocalMux I__857 (
            .O(N__8151),
            .I(\this_vga_signals.M_vstate_qZ0Z_0 ));
    Odrv4 I__856 (
            .O(N__8148),
            .I(\this_vga_signals.M_vstate_qZ0Z_0 ));
    LocalMux I__855 (
            .O(N__8145),
            .I(\this_vga_signals.M_vstate_qZ0Z_0 ));
    CascadeMux I__854 (
            .O(N__8138),
            .I(\this_vga_signals.M_vstate_q_srsts_0_a4_0_4_cascade_ ));
    InMux I__853 (
            .O(N__8135),
            .I(N__8132));
    LocalMux I__852 (
            .O(N__8132),
            .I(\this_vga_signals.M_vstate_q_srsts_0_a4_0_4 ));
    CascadeMux I__851 (
            .O(N__8129),
            .I(\this_vga_signals.N_230_0_cascade_ ));
    IoInMux I__850 (
            .O(N__8126),
            .I(N__8123));
    LocalMux I__849 (
            .O(N__8123),
            .I(N__8120));
    IoSpan4Mux I__848 (
            .O(N__8120),
            .I(N__8117));
    Span4Mux_s2_v I__847 (
            .O(N__8117),
            .I(N__8114));
    Sp12to4 I__846 (
            .O(N__8114),
            .I(N__8110));
    InMux I__845 (
            .O(N__8113),
            .I(N__8107));
    Span12Mux_h I__844 (
            .O(N__8110),
            .I(N__8104));
    LocalMux I__843 (
            .O(N__8107),
            .I(N__8101));
    Odrv12 I__842 (
            .O(N__8104),
            .I(vsync_c));
    Odrv4 I__841 (
            .O(N__8101),
            .I(vsync_c));
    InMux I__840 (
            .O(N__8096),
            .I(N__8091));
    InMux I__839 (
            .O(N__8095),
            .I(N__8088));
    InMux I__838 (
            .O(N__8094),
            .I(N__8085));
    LocalMux I__837 (
            .O(N__8091),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__836 (
            .O(N__8088),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__835 (
            .O(N__8085),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    InMux I__834 (
            .O(N__8078),
            .I(N__8073));
    InMux I__833 (
            .O(N__8077),
            .I(N__8070));
    InMux I__832 (
            .O(N__8076),
            .I(N__8067));
    LocalMux I__831 (
            .O(N__8073),
            .I(N__8064));
    LocalMux I__830 (
            .O(N__8070),
            .I(N__8061));
    LocalMux I__829 (
            .O(N__8067),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__828 (
            .O(N__8064),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__827 (
            .O(N__8061),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    CascadeMux I__826 (
            .O(N__8054),
            .I(N__8050));
    CascadeMux I__825 (
            .O(N__8053),
            .I(N__8046));
    InMux I__824 (
            .O(N__8050),
            .I(N__8042));
    InMux I__823 (
            .O(N__8049),
            .I(N__8037));
    InMux I__822 (
            .O(N__8046),
            .I(N__8037));
    InMux I__821 (
            .O(N__8045),
            .I(N__8034));
    LocalMux I__820 (
            .O(N__8042),
            .I(N__8031));
    LocalMux I__819 (
            .O(N__8037),
            .I(N__8028));
    LocalMux I__818 (
            .O(N__8034),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__817 (
            .O(N__8031),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__816 (
            .O(N__8028),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    InMux I__815 (
            .O(N__8021),
            .I(N__8018));
    LocalMux I__814 (
            .O(N__8018),
            .I(N__8015));
    Span4Mux_v I__813 (
            .O(N__8015),
            .I(N__8012));
    Odrv4 I__812 (
            .O(N__8012),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_1 ));
    InMux I__811 (
            .O(N__8009),
            .I(N__8006));
    LocalMux I__810 (
            .O(N__8006),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_6 ));
    InMux I__809 (
            .O(N__8003),
            .I(N__8000));
    LocalMux I__808 (
            .O(N__8000),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_2 ));
    InMux I__807 (
            .O(N__7997),
            .I(N__7994));
    LocalMux I__806 (
            .O(N__7994),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_3 ));
    InMux I__805 (
            .O(N__7991),
            .I(N__7988));
    LocalMux I__804 (
            .O(N__7988),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_4 ));
    InMux I__803 (
            .O(N__7985),
            .I(N__7982));
    LocalMux I__802 (
            .O(N__7982),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_5 ));
    InMux I__801 (
            .O(N__7979),
            .I(N__7976));
    LocalMux I__800 (
            .O(N__7976),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_13 ));
    InMux I__799 (
            .O(N__7973),
            .I(N__7970));
    LocalMux I__798 (
            .O(N__7970),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_11 ));
    InMux I__797 (
            .O(N__7967),
            .I(N__7964));
    LocalMux I__796 (
            .O(N__7964),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_12 ));
    InMux I__795 (
            .O(N__7961),
            .I(N__7958));
    LocalMux I__794 (
            .O(N__7958),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_9 ));
    InMux I__793 (
            .O(N__7955),
            .I(N__7952));
    LocalMux I__792 (
            .O(N__7952),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_10 ));
    CascadeMux I__791 (
            .O(N__7949),
            .I(\this_vga_signals.N_237_0_cascade_ ));
    InMux I__790 (
            .O(N__7946),
            .I(N__7943));
    LocalMux I__789 (
            .O(N__7943),
            .I(\this_vga_signals.M_vstate_d_0_sqmuxa ));
    CascadeMux I__788 (
            .O(N__7940),
            .I(N__7937));
    InMux I__787 (
            .O(N__7937),
            .I(N__7931));
    InMux I__786 (
            .O(N__7936),
            .I(N__7931));
    LocalMux I__785 (
            .O(N__7931),
            .I(\this_vga_signals.N_221_0 ));
    InMux I__784 (
            .O(N__7928),
            .I(N__7925));
    LocalMux I__783 (
            .O(N__7925),
            .I(\this_vga_signals.N_225_0 ));
    CascadeMux I__782 (
            .O(N__7922),
            .I(\this_vga_signals.N_225_0_cascade_ ));
    InMux I__781 (
            .O(N__7919),
            .I(N__7916));
    LocalMux I__780 (
            .O(N__7916),
            .I(\this_vga_signals.N_239_0 ));
    CascadeMux I__779 (
            .O(N__7913),
            .I(\this_vga_signals.N_239_0_cascade_ ));
    IoInMux I__778 (
            .O(N__7910),
            .I(N__7907));
    LocalMux I__777 (
            .O(N__7907),
            .I(N__7904));
    Span4Mux_s0_h I__776 (
            .O(N__7904),
            .I(N__7900));
    InMux I__775 (
            .O(N__7903),
            .I(N__7897));
    Sp12to4 I__774 (
            .O(N__7900),
            .I(N__7894));
    LocalMux I__773 (
            .O(N__7897),
            .I(N__7891));
    Span12Mux_v I__772 (
            .O(N__7894),
            .I(N__7887));
    Sp12to4 I__771 (
            .O(N__7891),
            .I(N__7884));
    InMux I__770 (
            .O(N__7890),
            .I(N__7881));
    Span12Mux_h I__769 (
            .O(N__7887),
            .I(N__7876));
    Span12Mux_v I__768 (
            .O(N__7884),
            .I(N__7873));
    LocalMux I__767 (
            .O(N__7881),
            .I(N__7870));
    InMux I__766 (
            .O(N__7880),
            .I(N__7867));
    InMux I__765 (
            .O(N__7879),
            .I(N__7864));
    Odrv12 I__764 (
            .O(N__7876),
            .I(port_nmib_c));
    Odrv12 I__763 (
            .O(N__7873),
            .I(port_nmib_c));
    Odrv4 I__762 (
            .O(N__7870),
            .I(port_nmib_c));
    LocalMux I__761 (
            .O(N__7867),
            .I(port_nmib_c));
    LocalMux I__760 (
            .O(N__7864),
            .I(port_nmib_c));
    CascadeMux I__759 (
            .O(N__7853),
            .I(\this_vga_signals.N_258_cascade_ ));
    InMux I__758 (
            .O(N__7850),
            .I(N__7847));
    LocalMux I__757 (
            .O(N__7847),
            .I(\this_vga_signals.N_238_0 ));
    InMux I__756 (
            .O(N__7844),
            .I(N__7838));
    InMux I__755 (
            .O(N__7843),
            .I(N__7838));
    LocalMux I__754 (
            .O(N__7838),
            .I(\this_vga_signals.M_vstate_qZ0Z_2 ));
    InMux I__753 (
            .O(N__7835),
            .I(bfn_13_18_0_));
    InMux I__752 (
            .O(N__7832),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_8 ));
    InMux I__751 (
            .O(N__7829),
            .I(N__7826));
    LocalMux I__750 (
            .O(N__7826),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_CO ));
    InMux I__749 (
            .O(N__7823),
            .I(N__7820));
    LocalMux I__748 (
            .O(N__7820),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_CO ));
    InMux I__747 (
            .O(N__7817),
            .I(N__7814));
    LocalMux I__746 (
            .O(N__7814),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_CO ));
    CascadeMux I__745 (
            .O(N__7811),
            .I(\this_vga_signals.N_238_0_cascade_ ));
    CascadeMux I__744 (
            .O(N__7808),
            .I(\this_vga_signals.N_221_0_cascade_ ));
    InMux I__743 (
            .O(N__7805),
            .I(N__7799));
    InMux I__742 (
            .O(N__7804),
            .I(N__7799));
    LocalMux I__741 (
            .O(N__7799),
            .I(\this_vga_signals.N_232_0 ));
    InMux I__740 (
            .O(N__7796),
            .I(N__7793));
    LocalMux I__739 (
            .O(N__7793),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_3 ));
    InMux I__738 (
            .O(N__7790),
            .I(N__7787));
    LocalMux I__737 (
            .O(N__7787),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_4 ));
    InMux I__736 (
            .O(N__7784),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_0 ));
    InMux I__735 (
            .O(N__7781),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_1 ));
    InMux I__734 (
            .O(N__7778),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_2 ));
    InMux I__733 (
            .O(N__7775),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_3 ));
    InMux I__732 (
            .O(N__7772),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_4 ));
    InMux I__731 (
            .O(N__7769),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_5 ));
    InMux I__730 (
            .O(N__7766),
            .I(\this_vga_signals.un1_M_vcounter_q_10_cry_6 ));
    InMux I__729 (
            .O(N__7763),
            .I(N__7756));
    InMux I__728 (
            .O(N__7762),
            .I(N__7756));
    InMux I__727 (
            .O(N__7761),
            .I(N__7753));
    LocalMux I__726 (
            .O(N__7756),
            .I(N__7748));
    LocalMux I__725 (
            .O(N__7753),
            .I(N__7748));
    Span4Mux_v I__724 (
            .O(N__7748),
            .I(N__7745));
    Span4Mux_v I__723 (
            .O(N__7745),
            .I(N__7742));
    Sp12to4 I__722 (
            .O(N__7742),
            .I(N__7739));
    Span12Mux_h I__721 (
            .O(N__7739),
            .I(N__7736));
    Odrv12 I__720 (
            .O(N__7736),
            .I(port_clk_c));
    InMux I__719 (
            .O(N__7733),
            .I(N__7729));
    InMux I__718 (
            .O(N__7732),
            .I(N__7726));
    LocalMux I__717 (
            .O(N__7729),
            .I(this_start_data_delay_this_edge_detector_M_last_q));
    LocalMux I__716 (
            .O(N__7726),
            .I(this_start_data_delay_this_edge_detector_M_last_q));
    InMux I__715 (
            .O(N__7721),
            .I(N__7718));
    LocalMux I__714 (
            .O(N__7718),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_0 ));
    InMux I__713 (
            .O(N__7715),
            .I(N__7712));
    LocalMux I__712 (
            .O(N__7712),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_1 ));
    InMux I__711 (
            .O(N__7709),
            .I(N__7706));
    LocalMux I__710 (
            .O(N__7706),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_2 ));
    InMux I__709 (
            .O(N__7703),
            .I(N__7700));
    LocalMux I__708 (
            .O(N__7700),
            .I(m16));
    InMux I__707 (
            .O(N__7697),
            .I(N__7694));
    LocalMux I__706 (
            .O(N__7694),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_8 ));
    InMux I__705 (
            .O(N__7691),
            .I(N__7688));
    LocalMux I__704 (
            .O(N__7688),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_6 ));
    InMux I__703 (
            .O(N__7685),
            .I(N__7682));
    LocalMux I__702 (
            .O(N__7682),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_7 ));
    InMux I__701 (
            .O(N__7679),
            .I(N__7676));
    LocalMux I__700 (
            .O(N__7676),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_5 ));
    InMux I__699 (
            .O(N__7673),
            .I(N__7670));
    LocalMux I__698 (
            .O(N__7670),
            .I(N__7667));
    Span4Mux_v I__697 (
            .O(N__7667),
            .I(N__7664));
    Odrv4 I__696 (
            .O(N__7664),
            .I(rgb_2_5_0__i2_mux_0));
    InMux I__695 (
            .O(N__7661),
            .I(N__7658));
    LocalMux I__694 (
            .O(N__7658),
            .I(N__7655));
    Odrv12 I__693 (
            .O(N__7655),
            .I(rgb_2_5_0__i2_mux));
    InMux I__692 (
            .O(N__7652),
            .I(N__7649));
    LocalMux I__691 (
            .O(N__7649),
            .I(N__7646));
    Span4Mux_v I__690 (
            .O(N__7646),
            .I(N__7643));
    Odrv4 I__689 (
            .O(N__7643),
            .I(m19));
    InMux I__688 (
            .O(N__7640),
            .I(N__7634));
    InMux I__687 (
            .O(N__7639),
            .I(N__7631));
    InMux I__686 (
            .O(N__7638),
            .I(N__7628));
    InMux I__685 (
            .O(N__7637),
            .I(N__7625));
    LocalMux I__684 (
            .O(N__7634),
            .I(N__7622));
    LocalMux I__683 (
            .O(N__7631),
            .I(N__7618));
    LocalMux I__682 (
            .O(N__7628),
            .I(N__7615));
    LocalMux I__681 (
            .O(N__7625),
            .I(N__7612));
    Span4Mux_v I__680 (
            .O(N__7622),
            .I(N__7608));
    InMux I__679 (
            .O(N__7621),
            .I(N__7605));
    Span4Mux_v I__678 (
            .O(N__7618),
            .I(N__7600));
    Span4Mux_v I__677 (
            .O(N__7615),
            .I(N__7600));
    Span4Mux_v I__676 (
            .O(N__7612),
            .I(N__7597));
    InMux I__675 (
            .O(N__7611),
            .I(N__7594));
    Span4Mux_v I__674 (
            .O(N__7608),
            .I(N__7589));
    LocalMux I__673 (
            .O(N__7605),
            .I(N__7589));
    Odrv4 I__672 (
            .O(N__7600),
            .I(rgb72));
    Odrv4 I__671 (
            .O(N__7597),
            .I(rgb72));
    LocalMux I__670 (
            .O(N__7594),
            .I(rgb72));
    Odrv4 I__669 (
            .O(N__7589),
            .I(rgb72));
    IoInMux I__668 (
            .O(N__7580),
            .I(N__7577));
    LocalMux I__667 (
            .O(N__7577),
            .I(N__7574));
    IoSpan4Mux I__666 (
            .O(N__7574),
            .I(N__7571));
    Sp12to4 I__665 (
            .O(N__7571),
            .I(N__7568));
    Span12Mux_s6_h I__664 (
            .O(N__7568),
            .I(N__7565));
    Odrv12 I__663 (
            .O(N__7565),
            .I(rgb_c_3));
    InMux I__662 (
            .O(N__7562),
            .I(N__7559));
    LocalMux I__661 (
            .O(N__7559),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_0 ));
    IoInMux I__660 (
            .O(N__7556),
            .I(N__7553));
    LocalMux I__659 (
            .O(N__7553),
            .I(N__7550));
    Span4Mux_s1_v I__658 (
            .O(N__7550),
            .I(N__7547));
    Span4Mux_v I__657 (
            .O(N__7547),
            .I(N__7544));
    Span4Mux_v I__656 (
            .O(N__7544),
            .I(N__7541));
    Odrv4 I__655 (
            .O(N__7541),
            .I(this_vga_signals_M_hstate_q_i_1));
    IoInMux I__654 (
            .O(N__7538),
            .I(N__7535));
    LocalMux I__653 (
            .O(N__7535),
            .I(N__7532));
    Span12Mux_s2_v I__652 (
            .O(N__7532),
            .I(N__7529));
    Odrv12 I__651 (
            .O(N__7529),
            .I(port_nmib_c_i));
    IoInMux I__650 (
            .O(N__7526),
            .I(N__7523));
    LocalMux I__649 (
            .O(N__7523),
            .I(N__7520));
    Odrv12 I__648 (
            .O(N__7520),
            .I(rgb_c_2));
    IoInMux I__647 (
            .O(N__7517),
            .I(N__7514));
    LocalMux I__646 (
            .O(N__7514),
            .I(N__7511));
    Span4Mux_s2_h I__645 (
            .O(N__7511),
            .I(N__7508));
    Span4Mux_h I__644 (
            .O(N__7508),
            .I(N__7505));
    Span4Mux_v I__643 (
            .O(N__7505),
            .I(N__7502));
    Odrv4 I__642 (
            .O(N__7502),
            .I(rgb_c_5));
    IoInMux I__641 (
            .O(N__7499),
            .I(N__7496));
    LocalMux I__640 (
            .O(N__7496),
            .I(N__7493));
    IoSpan4Mux I__639 (
            .O(N__7493),
            .I(N__7490));
    Span4Mux_s1_v I__638 (
            .O(N__7490),
            .I(N__7487));
    Span4Mux_v I__637 (
            .O(N__7487),
            .I(N__7484));
    Odrv4 I__636 (
            .O(N__7484),
            .I(this_vga_signals_M_hstate_q_i_4));
    IoInMux I__635 (
            .O(N__7481),
            .I(N__7478));
    LocalMux I__634 (
            .O(N__7478),
            .I(N__7475));
    Span12Mux_s8_h I__633 (
            .O(N__7475),
            .I(N__7472));
    Odrv12 I__632 (
            .O(N__7472),
            .I(rgb_c_4));
    IoInMux I__631 (
            .O(N__7469),
            .I(N__7466));
    LocalMux I__630 (
            .O(N__7466),
            .I(N__7463));
    IoSpan4Mux I__629 (
            .O(N__7463),
            .I(N__7460));
    IoSpan4Mux I__628 (
            .O(N__7460),
            .I(N__7457));
    Span4Mux_s3_h I__627 (
            .O(N__7457),
            .I(N__7454));
    Span4Mux_h I__626 (
            .O(N__7454),
            .I(N__7451));
    Odrv4 I__625 (
            .O(N__7451),
            .I(rgb_c_0));
    InMux I__624 (
            .O(N__7448),
            .I(N__7445));
    LocalMux I__623 (
            .O(N__7445),
            .I(N__7442));
    Odrv4 I__622 (
            .O(N__7442),
            .I(m5));
    IoInMux I__621 (
            .O(N__7439),
            .I(N__7436));
    LocalMux I__620 (
            .O(N__7436),
            .I(N__7433));
    Span12Mux_s9_h I__619 (
            .O(N__7433),
            .I(N__7430));
    Odrv12 I__618 (
            .O(N__7430),
            .I(rgb_c_1));
    IoInMux I__617 (
            .O(N__7427),
            .I(N__7424));
    LocalMux I__616 (
            .O(N__7424),
            .I(port_rw_c_i));
    SRMux I__615 (
            .O(N__7421),
            .I(N__7418));
    LocalMux I__614 (
            .O(N__7418),
            .I(N__7413));
    SRMux I__613 (
            .O(N__7417),
            .I(N__7410));
    SRMux I__612 (
            .O(N__7416),
            .I(N__7407));
    Span4Mux_v I__611 (
            .O(N__7413),
            .I(N__7397));
    LocalMux I__610 (
            .O(N__7410),
            .I(N__7397));
    LocalMux I__609 (
            .O(N__7407),
            .I(N__7397));
    SRMux I__608 (
            .O(N__7406),
            .I(N__7394));
    SRMux I__607 (
            .O(N__7405),
            .I(N__7391));
    SRMux I__606 (
            .O(N__7404),
            .I(N__7386));
    Span4Mux_v I__605 (
            .O(N__7397),
            .I(N__7377));
    LocalMux I__604 (
            .O(N__7394),
            .I(N__7377));
    LocalMux I__603 (
            .O(N__7391),
            .I(N__7377));
    SRMux I__602 (
            .O(N__7390),
            .I(N__7374));
    SRMux I__601 (
            .O(N__7389),
            .I(N__7370));
    LocalMux I__600 (
            .O(N__7386),
            .I(N__7367));
    SRMux I__599 (
            .O(N__7385),
            .I(N__7364));
    SRMux I__598 (
            .O(N__7384),
            .I(N__7361));
    Span4Mux_v I__597 (
            .O(N__7377),
            .I(N__7354));
    LocalMux I__596 (
            .O(N__7374),
            .I(N__7354));
    SRMux I__595 (
            .O(N__7373),
            .I(N__7351));
    LocalMux I__594 (
            .O(N__7370),
            .I(N__7346));
    Span4Mux_s1_v I__593 (
            .O(N__7367),
            .I(N__7339));
    LocalMux I__592 (
            .O(N__7364),
            .I(N__7339));
    LocalMux I__591 (
            .O(N__7361),
            .I(N__7339));
    SRMux I__590 (
            .O(N__7360),
            .I(N__7336));
    SRMux I__589 (
            .O(N__7359),
            .I(N__7333));
    Span4Mux_h I__588 (
            .O(N__7354),
            .I(N__7324));
    LocalMux I__587 (
            .O(N__7351),
            .I(N__7324));
    SRMux I__586 (
            .O(N__7350),
            .I(N__7321));
    SRMux I__585 (
            .O(N__7349),
            .I(N__7317));
    Span4Mux_v I__584 (
            .O(N__7346),
            .I(N__7305));
    Span4Mux_v I__583 (
            .O(N__7339),
            .I(N__7305));
    LocalMux I__582 (
            .O(N__7336),
            .I(N__7305));
    LocalMux I__581 (
            .O(N__7333),
            .I(N__7305));
    SRMux I__580 (
            .O(N__7332),
            .I(N__7302));
    SRMux I__579 (
            .O(N__7331),
            .I(N__7299));
    IoInMux I__578 (
            .O(N__7330),
            .I(N__7295));
    SRMux I__577 (
            .O(N__7329),
            .I(N__7292));
    Span4Mux_v I__576 (
            .O(N__7324),
            .I(N__7287));
    LocalMux I__575 (
            .O(N__7321),
            .I(N__7287));
    SRMux I__574 (
            .O(N__7320),
            .I(N__7284));
    LocalMux I__573 (
            .O(N__7317),
            .I(N__7278));
    SRMux I__572 (
            .O(N__7316),
            .I(N__7275));
    SRMux I__571 (
            .O(N__7315),
            .I(N__7270));
    SRMux I__570 (
            .O(N__7314),
            .I(N__7266));
    Span4Mux_v I__569 (
            .O(N__7305),
            .I(N__7259));
    LocalMux I__568 (
            .O(N__7302),
            .I(N__7259));
    LocalMux I__567 (
            .O(N__7299),
            .I(N__7259));
    SRMux I__566 (
            .O(N__7298),
            .I(N__7256));
    LocalMux I__565 (
            .O(N__7295),
            .I(N__7252));
    LocalMux I__564 (
            .O(N__7292),
            .I(N__7245));
    Span4Mux_h I__563 (
            .O(N__7287),
            .I(N__7245));
    LocalMux I__562 (
            .O(N__7284),
            .I(N__7245));
    SRMux I__561 (
            .O(N__7283),
            .I(N__7242));
    SRMux I__560 (
            .O(N__7282),
            .I(N__7239));
    SRMux I__559 (
            .O(N__7281),
            .I(N__7236));
    Span4Mux_v I__558 (
            .O(N__7278),
            .I(N__7231));
    LocalMux I__557 (
            .O(N__7275),
            .I(N__7231));
    SRMux I__556 (
            .O(N__7274),
            .I(N__7228));
    SRMux I__555 (
            .O(N__7273),
            .I(N__7225));
    LocalMux I__554 (
            .O(N__7270),
            .I(N__7222));
    SRMux I__553 (
            .O(N__7269),
            .I(N__7219));
    LocalMux I__552 (
            .O(N__7266),
            .I(N__7215));
    Span4Mux_v I__551 (
            .O(N__7259),
            .I(N__7210));
    LocalMux I__550 (
            .O(N__7256),
            .I(N__7210));
    SRMux I__549 (
            .O(N__7255),
            .I(N__7206));
    IoSpan4Mux I__548 (
            .O(N__7252),
            .I(N__7203));
    Span4Mux_v I__547 (
            .O(N__7245),
            .I(N__7198));
    LocalMux I__546 (
            .O(N__7242),
            .I(N__7198));
    LocalMux I__545 (
            .O(N__7239),
            .I(N__7195));
    LocalMux I__544 (
            .O(N__7236),
            .I(N__7192));
    Span4Mux_v I__543 (
            .O(N__7231),
            .I(N__7185));
    LocalMux I__542 (
            .O(N__7228),
            .I(N__7185));
    LocalMux I__541 (
            .O(N__7225),
            .I(N__7185));
    Span4Mux_v I__540 (
            .O(N__7222),
            .I(N__7180));
    LocalMux I__539 (
            .O(N__7219),
            .I(N__7180));
    SRMux I__538 (
            .O(N__7218),
            .I(N__7177));
    Span12Mux_h I__537 (
            .O(N__7215),
            .I(N__7174));
    Span4Mux_v I__536 (
            .O(N__7210),
            .I(N__7171));
    SRMux I__535 (
            .O(N__7209),
            .I(N__7168));
    LocalMux I__534 (
            .O(N__7206),
            .I(N__7165));
    Span4Mux_s2_h I__533 (
            .O(N__7203),
            .I(N__7162));
    Span4Mux_h I__532 (
            .O(N__7198),
            .I(N__7159));
    Span4Mux_s3_v I__531 (
            .O(N__7195),
            .I(N__7156));
    Span4Mux_s3_v I__530 (
            .O(N__7192),
            .I(N__7147));
    Span4Mux_v I__529 (
            .O(N__7185),
            .I(N__7147));
    Span4Mux_s3_v I__528 (
            .O(N__7180),
            .I(N__7147));
    LocalMux I__527 (
            .O(N__7177),
            .I(N__7147));
    Span12Mux_h I__526 (
            .O(N__7174),
            .I(N__7144));
    Sp12to4 I__525 (
            .O(N__7171),
            .I(N__7139));
    LocalMux I__524 (
            .O(N__7168),
            .I(N__7139));
    Span12Mux_h I__523 (
            .O(N__7165),
            .I(N__7136));
    Span4Mux_h I__522 (
            .O(N__7162),
            .I(N__7133));
    Span4Mux_v I__521 (
            .O(N__7159),
            .I(N__7126));
    Span4Mux_h I__520 (
            .O(N__7156),
            .I(N__7126));
    Span4Mux_h I__519 (
            .O(N__7147),
            .I(N__7126));
    Span12Mux_v I__518 (
            .O(N__7144),
            .I(N__7123));
    Span12Mux_h I__517 (
            .O(N__7139),
            .I(N__7120));
    Span12Mux_h I__516 (
            .O(N__7136),
            .I(N__7115));
    Sp12to4 I__515 (
            .O(N__7133),
            .I(N__7115));
    Sp12to4 I__514 (
            .O(N__7126),
            .I(N__7112));
    Span12Mux_v I__513 (
            .O(N__7123),
            .I(N__7109));
    Span12Mux_h I__512 (
            .O(N__7120),
            .I(N__7104));
    Span12Mux_v I__511 (
            .O(N__7115),
            .I(N__7104));
    Span12Mux_h I__510 (
            .O(N__7112),
            .I(N__7101));
    Odrv12 I__509 (
            .O(N__7109),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__508 (
            .O(N__7104),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__507 (
            .O(N__7101),
            .I(CONSTANT_ONE_NET));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_10_cry_7 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_23_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_9_0_));
    defparam IN_MUX_bfv_23_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_10_0_ (
            .carryinitin(\this_vga_signals.un1_M_vaddress_q_cry_7 ),
            .carryinitout(bfn_23_10_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(\this_vga_signals.un1_M_haddress_q_cry_7 ),
            .carryinitout(bfn_18_16_0_));
    ICE_GB \this_vga_signals.M_vstate_q_RNI3M6M4_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__8189),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_583_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNI6VB7_3  (
            .USERSIGNALTOGLOBALBUFFER(N__19510),
            .GLOBALBUFFEROUTPUT(N_631_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam port_data_rw_obuf_RNO_LC_1_22_4.C_ON=1'b0;
    defparam port_data_rw_obuf_RNO_LC_1_22_4.SEQ_MODE=4'b0000;
    defparam port_data_rw_obuf_RNO_LC_1_22_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 port_data_rw_obuf_RNO_LC_1_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18859),
            .lcout(port_rw_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_3_29_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_3_29_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_3_29_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_3_29_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNI1DID_1_LC_5_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNI1DID_1_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNI1DID_1_LC_5_23_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_hstate_q_RNI1DID_1_LC_5_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9833),
            .lcout(this_vga_signals_M_hstate_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNIFPC1_1_LC_5_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNIFPC1_1_LC_5_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNIFPC1_1_LC_5_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_vstate_q_RNIFPC1_1_LC_5_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7903),
            .lcout(port_nmib_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_obuf_RNO_2_LC_7_17_4.C_ON=1'b0;
    defparam rgb_obuf_RNO_2_LC_7_17_4.SEQ_MODE=4'b0000;
    defparam rgb_obuf_RNO_2_LC_7_17_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_obuf_RNO_2_LC_7_17_4 (
            .in0(N__7661),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7639),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_obuf_RNO_5_LC_7_20_6.C_ON=1'b0;
    defparam rgb_obuf_RNO_5_LC_7_20_6.SEQ_MODE=4'b0000;
    defparam rgb_obuf_RNO_5_LC_7_20_6.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_obuf_RNO_5_LC_7_20_6 (
            .in0(N__7673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7638),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNI4GID_4_LC_7_27_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNI4GID_4_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNI4GID_4_LC_7_27_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_hstate_q_RNI4GID_4_LC_7_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8675),
            .lcout(this_vga_signals_M_hstate_q_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_obuf_RNO_4_LC_9_21_1.C_ON=1'b0;
    defparam rgb_obuf_RNO_4_LC_9_21_1.SEQ_MODE=4'b0000;
    defparam rgb_obuf_RNO_4_LC_9_21_1.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_obuf_RNO_4_LC_9_21_1 (
            .in0(N__7652),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7637),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_obuf_RNO_0_LC_10_12_1.C_ON=1'b0;
    defparam rgb_obuf_RNO_0_LC_10_12_1.SEQ_MODE=4'b0000;
    defparam rgb_obuf_RNO_0_LC_10_12_1.LUT_INIT=16'b0001101000000000;
    LogicCell40 rgb_obuf_RNO_0_LC_10_12_1 (
            .in0(N__15566),
            .in1(N__11939),
            .in2(N__11458),
            .in3(N__7640),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m5_LC_10_16_0.C_ON=1'b0;
    defparam rgb_2_5_0__m5_LC_10_16_0.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m5_LC_10_16_0.LUT_INIT=16'b1010101000100010;
    LogicCell40 rgb_2_5_0__m5_LC_10_16_0 (
            .in0(N__11940),
            .in1(N__15584),
            .in2(_gnd_net_),
            .in3(N__15856),
            .lcout(m5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_obuf_RNO_1_LC_10_18_4.C_ON=1'b0;
    defparam rgb_obuf_RNO_1_LC_10_18_4.SEQ_MODE=4'b0000;
    defparam rgb_obuf_RNO_1_LC_10_18_4.LUT_INIT=16'b1010110000000000;
    LogicCell40 rgb_obuf_RNO_1_LC_10_18_4 (
            .in0(N__15865),
            .in1(N__7448),
            .in2(N__11495),
            .in3(N__7611),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m22_LC_10_19_5.C_ON=1'b0;
    defparam rgb_2_5_0__m22_LC_10_19_5.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m22_LC_10_19_5.LUT_INIT=16'b0001100001001111;
    LogicCell40 rgb_2_5_0__m22_LC_10_19_5 (
            .in0(N__11941),
            .in1(N__15590),
            .in2(N__15869),
            .in3(N__11493),
            .lcout(rgb_2_5_0__i2_mux_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m10_LC_11_17_7.C_ON=1'b0;
    defparam rgb_2_5_0__m10_LC_11_17_7.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m10_LC_11_17_7.LUT_INIT=16'b0001001101001111;
    LogicCell40 rgb_2_5_0__m10_LC_11_17_7 (
            .in0(N__15588),
            .in1(N__11958),
            .in2(N__15855),
            .in3(N__11485),
            .lcout(rgb_2_5_0__i2_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNIG6VE_1_LC_11_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNIG6VE_1_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNIG6VE_1_LC_11_19_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNIG6VE_1_LC_11_19_7  (
            .in0(N__9832),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7890),
            .lcout(rgb72),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m19_LC_11_20_4.C_ON=1'b0;
    defparam rgb_2_5_0__m19_LC_11_20_4.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m19_LC_11_20_4.LUT_INIT=16'b0011100001011011;
    LogicCell40 rgb_2_5_0__m19_LC_11_20_4 (
            .in0(N__15589),
            .in1(N__11962),
            .in2(N__15863),
            .in3(N__11492),
            .lcout(m19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_obuf_RNO_3_LC_11_21_0.C_ON=1'b0;
    defparam rgb_obuf_RNO_3_LC_11_21_0.SEQ_MODE=4'b0000;
    defparam rgb_obuf_RNO_3_LC_11_21_0.LUT_INIT=16'b0010001000100010;
    LogicCell40 rgb_obuf_RNO_3_LC_11_21_0 (
            .in0(N__7621),
            .in1(N__7703),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_1_LC_12_14_1 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_1_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_1_LC_12_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_1_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7562),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19139),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_last_q_LC_12_14_2 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_last_q_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_edge_detector.M_last_q_LC_12_14_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_last_q_LC_12_14_2  (
            .in0(N__7763),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13168),
            .lcout(this_start_data_delay_this_edge_detector_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19139),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_0_LC_12_14_7 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_0_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_0_LC_12_14_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_0_LC_12_14_7  (
            .in0(N__13167),
            .in1(N__7762),
            .in2(_gnd_net_),
            .in3(N__7732),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19139),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_3_LC_12_15_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_3_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_3_LC_12_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_3_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7709),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19146),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_0_LC_12_15_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_0_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_0_LC_12_15_5 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_0_LC_12_15_5  (
            .in0(N__13166),
            .in1(N__7761),
            .in2(_gnd_net_),
            .in3(N__7733),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19146),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_1_LC_12_15_6 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_1_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_1_LC_12_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_1_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7721),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19146),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_2_LC_12_15_7 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_2_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_2_LC_12_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_2_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7715),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19146),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m16_LC_12_20_1.C_ON=1'b0;
    defparam rgb_2_5_0__m16_LC_12_20_1.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m16_LC_12_20_1.LUT_INIT=16'b0100100100011111;
    LogicCell40 rgb_2_5_0__m16_LC_12_20_1 (
            .in0(N__15565),
            .in1(N__15864),
            .in2(N__11966),
            .in3(N__11494),
            .lcout(m16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_6_LC_13_14_2 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_6_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_6_LC_13_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_6_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7679),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19132),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_8_LC_13_14_3 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_8_LC_13_14_3 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_8_LC_13_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_8_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7685),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19132),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_9_LC_13_14_4 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_9_LC_13_14_4 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_9_LC_13_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_9_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7697),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19132),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_7_LC_13_14_6 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_7_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_7_LC_13_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_7_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7691),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19132),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_5_LC_13_14_7 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_5_LC_13_14_7 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_5_LC_13_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_5_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7790),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19132),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_4_LC_13_15_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_4_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_4_LC_13_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_4_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7796),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19140),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_0_c_LC_13_17_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_0_c_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_0_c_LC_13_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_10_cry_0_c_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__14099),
            .in2(N__8615),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_10_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_LUT4_0_LC_13_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_LUT4_0_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_LUT4_0_LC_13_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_LUT4_0_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__8408),
            .in2(_gnd_net_),
            .in3(N__7784),
            .lcout(\this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_10_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_10_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_LUT4_0_LC_13_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_LUT4_0_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_LUT4_0_LC_13_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_LUT4_0_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__8372),
            .in2(_gnd_net_),
            .in3(N__7781),
            .lcout(\this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_10_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_10_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_LUT4_0_LC_13_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_LUT4_0_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_LUT4_0_LC_13_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_LUT4_0_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__8294),
            .in2(_gnd_net_),
            .in3(N__7778),
            .lcout(\this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_10_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_10_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_LC_13_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_4_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_LC_13_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__8329),
            .in2(_gnd_net_),
            .in3(N__7775),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_10_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_10_cry_4 ),
            .clk(N__19153),
            .ce(),
            .sr(N__17803));
    defparam \this_vga_signals.M_vcounter_q_5_LC_13_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_5_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_LC_13_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__8076),
            .in2(_gnd_net_),
            .in3(N__7772),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_10_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_10_cry_5 ),
            .clk(N__19153),
            .ce(),
            .sr(N__17803));
    defparam \this_vga_signals.M_vcounter_q_6_LC_13_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_6_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_LC_13_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__8045),
            .in2(_gnd_net_),
            .in3(N__7769),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_10_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_10_cry_6 ),
            .clk(N__19153),
            .ce(),
            .sr(N__17803));
    defparam \this_vga_signals.M_vcounter_q_7_LC_13_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_7_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_LC_13_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__8581),
            .in2(_gnd_net_),
            .in3(N__7766),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_10_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_10_cry_7 ),
            .clk(N__19153),
            .ce(),
            .sr(N__17803));
    defparam \this_vga_signals.M_vcounter_q_8_LC_13_18_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_8_LC_13_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_LC_13_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__8536),
            .in2(_gnd_net_),
            .in3(N__7835),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_10_cry_8 ),
            .clk(N__19160),
            .ce(),
            .sr(N__17800));
    defparam \this_vga_signals.M_vcounter_q_9_LC_13_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_9_LC_13_18_1 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_LC_13_18_1  (
            .in0(N__8509),
            .in1(N__8096),
            .in2(N__8470),
            .in3(N__7832),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19160),
            .ce(),
            .sr(N__17800));
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_18_3 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_13_18_3  (
            .in0(N__8508),
            .in1(N__8295),
            .in2(N__8472),
            .in3(N__7829),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19160),
            .ce(),
            .sr(N__17800));
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_18_4 .LUT_INIT=16'b0000011101110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_13_18_4  (
            .in0(N__8476),
            .in1(N__8507),
            .in2(N__8378),
            .in3(N__7823),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19160),
            .ce(),
            .sr(N__17800));
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_18_5 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_13_18_5  (
            .in0(N__8506),
            .in1(N__8415),
            .in2(N__8471),
            .in3(N__7817),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19160),
            .ce(),
            .sr(N__17800));
    defparam \this_vga_signals.M_vcounter_q_RNIHOM62_6_LC_13_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIHOM62_6_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIHOM62_6_LC_13_19_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIHOM62_6_LC_13_19_0  (
            .in0(N__8330),
            .in1(N__8406),
            .in2(N__8053),
            .in3(N__7928),
            .lcout(\this_vga_signals.N_232_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_7_LC_13_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_7_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_7_LC_13_19_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIFUDD4_7_LC_13_19_2  (
            .in0(N__7805),
            .in1(N__8534),
            .in2(N__7940),
            .in3(N__8584),
            .lcout(\this_vga_signals.N_238_0 ),
            .ltout(\this_vga_signals.N_238_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_1_LC_13_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_1_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_1_LC_13_19_3 .LUT_INIT=16'b0011001100000010;
    LogicCell40 \this_vga_signals.M_vstate_q_1_LC_13_19_3  (
            .in0(N__7879),
            .in1(N__19476),
            .in2(N__7811),
            .in3(N__7946),
            .lcout(port_nmib_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19164),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNILPDA1_9_LC_13_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNILPDA1_9_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNILPDA1_9_LC_13_19_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNILPDA1_9_LC_13_19_4  (
            .in0(N__8094),
            .in1(N__8077),
            .in2(_gnd_net_),
            .in3(N__8613),
            .lcout(\this_vga_signals.N_221_0 ),
            .ltout(\this_vga_signals.N_221_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_1_7_LC_13_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_1_7_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_1_7_LC_13_19_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIFUDD4_1_7_LC_13_19_5  (
            .in0(N__8530),
            .in1(N__8582),
            .in2(N__7808),
            .in3(N__7804),
            .lcout(\this_vga_signals.N_237_0 ),
            .ltout(\this_vga_signals.N_237_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_0_1_LC_13_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_0_1_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_0_1_LC_13_19_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_0_1_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7949),
            .in3(N__8159),
            .lcout(\this_vga_signals.M_vstate_d_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIHQRK2_6_LC_13_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIHQRK2_6_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIHQRK2_6_LC_13_19_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIHQRK2_6_LC_13_19_7  (
            .in0(N__8583),
            .in1(N__7936),
            .in2(N__8537),
            .in3(N__8049),
            .lcout(\this_vga_signals.N_226_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_3_LC_13_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_3_LC_13_20_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_3_LC_13_20_0 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \this_vga_signals.M_vstate_q_3_LC_13_20_0  (
            .in0(N__8207),
            .in1(N__7844),
            .in2(N__19509),
            .in3(N__7919),
            .lcout(\this_vga_signals.M_vstate_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19168),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_13_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_13_20_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__8296),
            .in2(_gnd_net_),
            .in3(N__8376),
            .lcout(\this_vga_signals.N_225_0 ),
            .ltout(\this_vga_signals.N_225_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_1_LC_13_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_1_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_1_LC_13_20_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIFUDD4_1_LC_13_20_5  (
            .in0(N__8227),
            .in1(N__8331),
            .in2(N__7922),
            .in3(N__8417),
            .lcout(\this_vga_signals.N_239_0 ),
            .ltout(\this_vga_signals.N_239_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_0_2_LC_13_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_0_2_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_0_2_LC_13_20_6 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_0_2_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__7843),
            .in2(N__7913),
            .in3(N__19479),
            .lcout(),
            .ltout(\this_vga_signals.N_258_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_2_LC_13_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_2_LC_13_20_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_2_LC_13_20_7 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \this_vga_signals.M_vstate_q_2_LC_13_20_7  (
            .in0(N__19480),
            .in1(N__7880),
            .in2(N__7853),
            .in3(N__7850),
            .lcout(\this_vga_signals.M_vstate_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19168),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_7_LC_14_13_0 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_7_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_7_LC_14_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_7_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8009),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19121),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_2_LC_14_13_3 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_2_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_2_LC_14_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_2_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8021),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19121),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_6_LC_14_13_4 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_6_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_6_LC_14_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_6_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7985),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19121),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_3_LC_14_13_5 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_3_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_3_LC_14_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_3_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8003),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19121),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_4_LC_14_13_6 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_4_LC_14_13_6 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_4_LC_14_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_4_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7997),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19121),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_5_LC_14_13_7 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_5_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_5_LC_14_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_5_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7991),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19121),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_14_LC_14_14_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_14_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_14_LC_14_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_14_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7979),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19127),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_11_LC_14_14_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_11_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_11_LC_14_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_11_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7955),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19127),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_13_LC_14_14_3 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_13_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_13_LC_14_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_13_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7967),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19127),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_12_LC_14_14_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_12_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_12_LC_14_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_12_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7973),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19127),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_10_LC_14_14_7 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_10_LC_14_14_7 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_10_LC_14_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_10_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7961),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19127),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNI3M6M4_0_LC_14_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNI3M6M4_0_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNI3M6M4_0_LC_14_17_1 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \this_vga_signals.M_vstate_q_RNI3M6M4_0_LC_14_17_1  (
            .in0(N__8154),
            .in1(N__19468),
            .in2(_gnd_net_),
            .in3(N__8174),
            .lcout(\this_vga_signals.M_vstate_q_RNI3M6M4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_14_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_0_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_14_17_7 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_14_17_7  (
            .in0(N__8510),
            .in1(N__8612),
            .in2(N__8477),
            .in3(N__14100),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19147),
            .ce(),
            .sr(N__17801));
    defparam \this_vga_signals.M_vstate_q_RNO_0_0_LC_14_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_0_0_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_0_0_LC_14_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_0_0_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__8454),
            .in2(_gnd_net_),
            .in3(N__8502),
            .lcout(),
            .ltout(\this_vga_signals.N_251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_0_LC_14_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_0_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_0_LC_14_18_4 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \this_vga_signals.M_vstate_q_0_LC_14_18_4  (
            .in0(N__19481),
            .in1(N__8158),
            .in2(N__8177),
            .in3(N__8173),
            .lcout(\this_vga_signals.M_vstate_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19154),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNIORO8_4_LC_14_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNIORO8_4_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNIORO8_4_LC_14_19_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNIORO8_4_LC_14_19_0  (
            .in0(N__19474),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8113),
            .lcout(\this_vga_signals.M_vstate_q_srsts_0_a4_0_4 ),
            .ltout(\this_vga_signals.M_vstate_q_srsts_0_a4_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_5_LC_14_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_5_LC_14_19_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_5_LC_14_19_1 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \this_vga_signals.M_vstate_q_5_LC_14_19_1  (
            .in0(N__8552),
            .in1(N__8423),
            .in2(N__8138),
            .in3(N__8231),
            .lcout(\this_vga_signals.M_vstate_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19161),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIU3IO1_2_LC_14_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIU3IO1_2_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIU3IO1_2_LC_14_19_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIU3IO1_2_LC_14_19_2  (
            .in0(N__8407),
            .in1(N__8290),
            .in2(N__8338),
            .in3(N__8371),
            .lcout(\this_vga_signals.N_230_0 ),
            .ltout(\this_vga_signals.N_230_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_4_LC_14_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_4_LC_14_19_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_4_LC_14_19_3 .LUT_INIT=16'b1100111011101110;
    LogicCell40 \this_vga_signals.M_vstate_q_4_LC_14_19_3  (
            .in0(N__8135),
            .in1(N__8258),
            .in2(N__8129),
            .in3(N__8230),
            .lcout(vsync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19161),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI8EIO1_9_LC_14_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI8EIO1_9_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI8EIO1_9_LC_14_19_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI8EIO1_9_LC_14_19_4  (
            .in0(N__8095),
            .in1(N__8078),
            .in2(N__8054),
            .in3(N__8614),
            .lcout(),
            .ltout(\this_vga_signals.M_vstate_q_srsts_0_o2_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_0_7_LC_14_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_0_7_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIFUDD4_0_7_LC_14_19_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIFUDD4_0_7_LC_14_19_5  (
            .in0(N__8585),
            .in1(N__8551),
            .in2(N__8540),
            .in3(N__8535),
            .lcout(\this_vga_signals.N_248_0 ),
            .ltout(\this_vga_signals.N_248_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_0_5_LC_14_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_0_5_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_0_5_LC_14_19_6 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_0_5_LC_14_19_6  (
            .in0(N__19475),
            .in1(_gnd_net_),
            .in2(N__8480),
            .in3(N__8453),
            .lcout(\this_vga_signals.N_252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIU3IO1_0_2_LC_14_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIU3IO1_0_2_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIU3IO1_0_2_LC_14_20_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIU3IO1_0_2_LC_14_20_2  (
            .in0(N__8416),
            .in1(N__8377),
            .in2(N__8339),
            .in3(N__8297),
            .lcout(\this_vga_signals.M_vstate_q_srsts_0_o2_2_3 ),
            .ltout(\this_vga_signals.M_vstate_q_srsts_0_o2_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_0_4_LC_14_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_0_4_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_0_4_LC_14_20_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_0_4_LC_14_20_3  (
            .in0(N__8242),
            .in1(N__19477),
            .in2(N__8261),
            .in3(N__8229),
            .lcout(\this_vga_signals.N_255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_0_3_LC_14_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_0_3_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_0_3_LC_14_20_7 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_0_3_LC_14_20_7  (
            .in0(N__8249),
            .in1(N__19478),
            .in2(N__8243),
            .in3(N__8228),
            .lcout(\this_vga_signals.N_256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_8_LC_15_13_0 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_8_LC_15_13_0 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_8_LC_15_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_8_LC_15_13_0  (
            .in0(N__8201),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19117),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_11_LC_15_13_2 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_11_LC_15_13_2 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_11_LC_15_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_11_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8195),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19117),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_10_LC_15_13_3 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_10_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_10_LC_15_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_10_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8633),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19117),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_12_LC_15_13_4 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_12_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_12_LC_15_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_12_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8645),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19117),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_9_LC_15_13_6 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_9_LC_15_13_6 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_9_LC_15_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_9_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8639),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19117),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_15_LC_15_14_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_15_LC_15_14_1 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_15_LC_15_14_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_15_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__8627),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19122),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_0_5_LC_15_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_0_5_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_0_5_LC_15_16_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_0_5_LC_15_16_4  (
            .in0(N__19445),
            .in1(N__8837),
            .in2(_gnd_net_),
            .in3(N__8852),
            .lcout(),
            .ltout(\this_vga_signals.N_417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_5_LC_15_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_5_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_5_LC_15_16_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \this_vga_signals.M_hstate_q_5_LC_15_16_5  (
            .in0(N__8693),
            .in1(N__8774),
            .in2(N__8621),
            .in3(N__8800),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19133),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI42JJ3_1_10_LC_15_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI42JJ3_1_10_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI42JJ3_1_10_LC_15_17_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI42JJ3_1_10_LC_15_17_0  (
            .in0(N__8816),
            .in1(N__9521),
            .in2(N__8778),
            .in3(N__8956),
            .lcout(\this_vga_signals.N_398_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_16_LC_15_17_2 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_16_LC_15_17_2 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_16_LC_15_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_16_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9425),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19141),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_0_2_LC_15_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_0_2_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_0_2_LC_15_17_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_0_2_LC_15_17_3  (
            .in0(N__8972),
            .in1(N__8930),
            .in2(N__9824),
            .in3(N__19469),
            .lcout(),
            .ltout(\this_vga_signals.N_412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_2_LC_15_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_2_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_2_LC_15_17_4 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \this_vga_signals.M_hstate_q_2_LC_15_17_4  (
            .in0(N__19470),
            .in1(N__8734),
            .in2(N__8618),
            .in3(N__8719),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19141),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_0_7_LC_15_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_0_7_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_0_7_LC_15_17_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIDR6I_0_7_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__9572),
            .in2(_gnd_net_),
            .in3(N__9596),
            .lcout(\this_vga_signals.N_390_0 ),
            .ltout(\this_vga_signals.N_390_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI42JJ3_10_LC_15_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI42JJ3_10_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI42JJ3_10_LC_15_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI42JJ3_10_LC_15_17_7  (
            .in0(N__9520),
            .in1(N__8955),
            .in2(N__8747),
            .in3(N__8815),
            .lcout(\this_vga_signals.N_397_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_0_4_LC_15_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_0_4_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_0_4_LC_15_18_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_0_4_LC_15_18_1  (
            .in0(N__8743),
            .in1(N__19533),
            .in2(N__8707),
            .in3(N__8798),
            .lcout(\this_vga_signals.N_416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_0_3_LC_15_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_0_3_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_0_3_LC_15_18_3 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_0_3_LC_15_18_3  (
            .in0(N__8744),
            .in1(N__19534),
            .in2(N__8708),
            .in3(N__8799),
            .lcout(),
            .ltout(\this_vga_signals.N_413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_3_LC_15_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_3_LC_15_18_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_3_LC_15_18_4 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \this_vga_signals.M_hstate_q_3_LC_15_18_4  (
            .in0(N__19535),
            .in1(N__8735),
            .in2(N__8723),
            .in3(N__8720),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19148),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNIAFUK_4_LC_15_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNIAFUK_4_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNIAFUK_4_LC_15_19_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hstate_q_RNIAFUK_4_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__8662),
            .in2(_gnd_net_),
            .in3(N__19473),
            .lcout(\this_vga_signals.M_hstate_q_srsts_0_a3_0_4 ),
            .ltout(\this_vga_signals.M_hstate_q_srsts_0_a3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_4_LC_15_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_4_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_4_LC_15_19_2 .LUT_INIT=16'b1101110011111100;
    LogicCell40 \this_vga_signals.M_hstate_q_4_LC_15_19_2  (
            .in0(N__8804),
            .in1(N__8684),
            .in2(N__8678),
            .in3(N__8780),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19155),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_13_LC_16_13_7 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_13_LC_16_13_7 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_13_LC_16_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_13_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8651),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19116),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_0_1_LC_16_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_0_1_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_0_1_LC_16_16_1 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_0_1_LC_16_16_1  (
            .in0(N__8929),
            .in1(N__8971),
            .in2(N__9816),
            .in3(N__19376),
            .lcout(\this_vga_signals.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNI9J514_5_LC_16_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNI9J514_5_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNI9J514_5_LC_16_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hstate_q_RNI9J514_5_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__8835),
            .in2(_gnd_net_),
            .in3(N__8850),
            .lcout(\this_vga_signals.M_hstate_d_0_sqmuxa ),
            .ltout(\this_vga_signals.M_hstate_d_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_0_LC_16_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_0_LC_16_16_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_0_LC_16_16_3 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \this_vga_signals.M_hstate_q_0_LC_16_16_3  (
            .in0(N__8870),
            .in1(N__8876),
            .in2(N__8879),
            .in3(N__19378),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19126),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI42JJ3_0_10_LC_16_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI42JJ3_0_10_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI42JJ3_0_10_LC_16_16_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI42JJ3_0_10_LC_16_16_5  (
            .in0(N__8928),
            .in1(N__9524),
            .in2(N__8779),
            .in3(N__8957),
            .lcout(\this_vga_signals.N_405_0 ),
            .ltout(\this_vga_signals.N_405_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_1_LC_16_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_1_LC_16_16_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_1_LC_16_16_6 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \this_vga_signals.M_hstate_q_1_LC_16_16_6  (
            .in0(N__19377),
            .in1(N__8869),
            .in2(N__8861),
            .in3(N__8858),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19126),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNIFIH84_5_LC_16_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNIFIH84_5_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNIFIH84_5_LC_16_16_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \this_vga_signals.M_hstate_q_RNIFIH84_5_LC_16_16_7  (
            .in0(N__8851),
            .in1(N__19375),
            .in2(_gnd_net_),
            .in3(N__8836),
            .lcout(\this_vga_signals.M_hstate_q_RNIFIH84Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_16_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_16_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_16_17_1  (
            .in0(N__9349),
            .in1(N__9364),
            .in2(N__9335),
            .in3(N__9381),
            .lcout(\this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5 ),
            .ltout(\this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_16_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_16_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_16_17_2  (
            .in0(N__9480),
            .in1(N__9409),
            .in2(N__8819),
            .in3(N__9315),
            .lcout(\this_vga_signals.N_385_0 ),
            .ltout(\this_vga_signals.N_385_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIN6C13_6_LC_16_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIN6C13_6_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIN6C13_6_LC_16_17_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIN6C13_6_LC_16_17_3  (
            .in0(N__9295),
            .in1(N__9523),
            .in2(N__8807),
            .in3(N__9547),
            .lcout(\this_vga_signals.N_391_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_7_LC_16_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_7_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_7_LC_16_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIDR6I_7_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__9570),
            .in2(_gnd_net_),
            .in3(N__9594),
            .lcout(\this_vga_signals.N_386_0 ),
            .ltout(\this_vga_signals.N_386_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_16_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_16_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_16_17_5  (
            .in0(N__9294),
            .in1(N__9522),
            .in2(N__8975),
            .in3(N__9546),
            .lcout(\this_vga_signals.M_hstate_q_srsts_0_o3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_6_LC_16_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_6_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_6_LC_16_17_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIDR6I_6_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__9545),
            .in2(_gnd_net_),
            .in3(N__9293),
            .lcout(\this_vga_signals.N_388_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_0_11_LC_16_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_0_11_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_0_11_LC_16_17_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIQFS22_0_11_LC_16_17_7  (
            .in0(N__9410),
            .in1(N__9481),
            .in2(N__8939),
            .in3(N__9316),
            .lcout(\this_vga_signals.N_393_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_0_LC_16_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_16_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_16_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9412),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19138),
            .ce(),
            .sr(N__17795));
    defparam \this_vga_signals.M_hcounter_q_1_LC_16_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_16_18_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_16_18_2  (
            .in0(N__9413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9385),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19138),
            .ce(),
            .sr(N__17795));
    defparam \this_reset_cond.M_stage_q_2_LC_17_9_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_17_9_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_17_9_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__8908),
            .in2(_gnd_net_),
            .in3(N__8885),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19110),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_17_9_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_17_9_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__8909),
            .in2(_gnd_net_),
            .in3(N__8915),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19110),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_17_9_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_17_9_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_17_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8906),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19110),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_17_9_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_17_9_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_17_9_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_17_9_7  (
            .in0(N__8907),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8891),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19110),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g2_2_LC_17_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g2_2_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g2_2_LC_17_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un14_address_g2_2_LC_17_10_1  (
            .in0(N__15353),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12357),
            .lcout(),
            .ltout(\this_vga_signals.g2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_4_LC_17_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_4_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_4_LC_17_10_2 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \this_vga_signals.un14_address_g1_4_LC_17_10_2  (
            .in0(N__15124),
            .in1(N__14502),
            .in2(N__9113),
            .in3(N__12677),
            .lcout(),
            .ltout(\this_vga_signals.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_1_4_LC_17_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_1_4_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_1_4_LC_17_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un14_address_g1_1_4_LC_17_10_3  (
            .in0(N__9467),
            .in1(N__10274),
            .in2(N__9110),
            .in3(N__17658),
            .lcout(\this_vga_signals.g1_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g2_4_LC_17_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g2_4_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g2_4_LC_17_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un14_address_g2_4_LC_17_10_6  (
            .in0(N__12356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15352),
            .lcout(),
            .ltout(\this_vga_signals.g2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_6_LC_17_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_6_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_6_LC_17_10_7 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \this_vga_signals.un14_address_g1_6_LC_17_10_7  (
            .in0(N__14501),
            .in1(N__15123),
            .in2(N__9107),
            .in3(N__11240),
            .lcout(\this_vga_signals.g1_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_14_N_8L16_LC_17_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_14_N_8L16_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_14_N_8L16_LC_17_11_0 .LUT_INIT=16'b0000011000001001;
    LogicCell40 \this_vga_signals.un14_address_g0_14_N_8L16_LC_17_11_0  (
            .in0(N__9257),
            .in1(N__17662),
            .in2(N__11516),
            .in3(N__9263),
            .lcout(),
            .ltout(\this_vga_signals.g0_14_N_8L16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_14_LC_17_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_14_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_14_LC_17_11_1 .LUT_INIT=16'b0000011011110110;
    LogicCell40 \this_vga_signals.un14_address_g0_14_LC_17_11_1  (
            .in0(N__12659),
            .in1(N__9104),
            .in2(N__9098),
            .in3(N__9683),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_LC_17_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_LC_17_11_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un14_address_g0_LC_17_11_2  (
            .in0(N__9620),
            .in1(N__9611),
            .in2(N__9095),
            .in3(N__9662),
            .lcout(this_vga_signals_un14_address_if_generate_plus_mult1_un75_sum_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_1_LC_17_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_1_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_1_LC_17_11_3 .LUT_INIT=16'b0000111011110001;
    LogicCell40 \this_vga_signals.un14_address_g0_1_LC_17_11_3  (
            .in0(N__12362),
            .in1(N__12630),
            .in2(N__15389),
            .in3(N__14906),
            .lcout(),
            .ltout(\this_vga_signals.if_N_2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_0_LC_17_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_0_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_0_LC_17_11_4 .LUT_INIT=16'b0011001011101100;
    LogicCell40 \this_vga_signals.un14_address_g0_0_LC_17_11_4  (
            .in0(N__13963),
            .in1(N__11264),
            .in2(N__9266),
            .in3(N__14507),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_14_N_7L14_LC_17_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_14_N_7L14_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_14_N_7L14_LC_17_11_5 .LUT_INIT=16'b0001111011100001;
    LogicCell40 \this_vga_signals.un14_address_g0_14_N_7L14_LC_17_11_5  (
            .in0(N__12363),
            .in1(N__12631),
            .in2(N__9605),
            .in3(N__9644),
            .lcout(\this_vga_signals.g0_14_N_7L14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m5_e_LC_17_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m5_e_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m5_e_LC_17_13_0 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \this_vga_signals.un6_address_if_m5_e_LC_17_13_0  (
            .in0(N__11699),
            .in1(_gnd_net_),
            .in2(N__11373),
            .in3(N__9248),
            .lcout(),
            .ltout(\this_vga_signals.if_N_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m5_LC_17_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m5_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m5_LC_17_13_1 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \this_vga_signals.un6_address_if_m5_LC_17_13_1  (
            .in0(N__19852),
            .in1(N__11366),
            .in2(N__9251),
            .in3(N__19904),
            .lcout(\this_vga_signals.if_i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_3_s_LC_17_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_3_s_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_3_s_LC_17_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_3_s_LC_17_13_2  (
            .in0(N__11437),
            .in1(N__11408),
            .in2(_gnd_net_),
            .in3(N__19851),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_3_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axb1_LC_17_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axb1_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axb1_LC_17_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axb1_LC_17_13_3  (
            .in0(N__10007),
            .in1(N__10202),
            .in2(_gnd_net_),
            .in3(N__10175),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m3_1_2_LC_17_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m3_1_2_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m3_1_2_LC_17_13_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un6_address_if_m3_1_2_LC_17_13_4  (
            .in0(N__11362),
            .in1(N__11430),
            .in2(N__9242),
            .in3(N__19850),
            .lcout(),
            .ltout(\this_vga_signals.if_m3_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m5_i_LC_17_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m5_i_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m5_i_LC_17_13_5 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \this_vga_signals.un6_address_if_m5_i_LC_17_13_5  (
            .in0(N__11409),
            .in1(N__10031),
            .in2(N__9239),
            .in3(N__9749),
            .lcout(),
            .ltout(\this_vga_signals.if_N_6_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un75_sum_i_3_LC_17_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un75_sum_i_3_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un75_sum_i_3_LC_17_13_6 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un75_sum_i_3_LC_17_13_6  (
            .in0(N__9236),
            .in1(N__9230),
            .in2(N__9224),
            .in3(N__9740),
            .lcout(this_vga_signals_un6_address_if_generate_plus_mult1_un75_sum_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m2_LC_17_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m2_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m2_LC_17_14_1 .LUT_INIT=16'b0010100000010100;
    LogicCell40 \this_vga_signals.un6_address_if_m2_LC_17_14_1  (
            .in0(N__10874),
            .in1(N__9924),
            .in2(N__10000),
            .in3(N__10577),
            .lcout(\this_vga_signals.if_m2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m3_3_LC_17_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m3_3_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m3_3_LC_17_14_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \this_vga_signals.un6_address_if_m3_3_LC_17_14_2  (
            .in0(N__10578),
            .in1(N__9923),
            .in2(_gnd_net_),
            .in3(N__10873),
            .lcout(\this_vga_signals.if_i1_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_17_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_17_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_17_14_4  (
            .in0(N__10177),
            .in1(N__11677),
            .in2(N__10006),
            .in3(N__10204),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_c2_LC_17_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_c2_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_c2_LC_17_14_5 .LUT_INIT=16'b0010101110001110;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_c2_LC_17_14_5  (
            .in0(N__9984),
            .in1(N__10203),
            .in2(N__11694),
            .in3(N__10176),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_14_LC_17_14_7 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_14_LC_17_14_7 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_14_LC_17_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_14_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9275),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19123),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m3_0_0_LC_17_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m3_0_0_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m3_0_0_LC_17_15_0 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \this_vga_signals.un6_address_if_m3_0_0_LC_17_15_0  (
            .in0(N__13470),
            .in1(N__13659),
            .in2(_gnd_net_),
            .in3(N__13578),
            .lcout(\this_vga_signals.if_m3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_1_LC_17_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_1_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_1_LC_17_15_1 .LUT_INIT=16'b1101111011001110;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_1_LC_17_15_1  (
            .in0(N__13657),
            .in1(N__13576),
            .in2(N__13503),
            .in3(N__13380),
            .lcout(\this_vga_signals.mult1_un40_sum_0_ac0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_1_LC_17_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_1_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_1_LC_17_15_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_1_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__13575),
            .in2(_gnd_net_),
            .in3(N__13379),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_0_ac0_3_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_LC_17_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_LC_17_15_4 .LUT_INIT=16'b1111110011110111;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_LC_17_15_4  (
            .in0(N__10861),
            .in1(N__13483),
            .in2(N__9269),
            .in3(N__13658),
            .lcout(\this_vga_signals.mult1_un40_sum_0_ac0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_a1_0_LC_17_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_a1_0_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_a1_0_LC_17_15_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_a1_0_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__13471),
            .in2(_gnd_net_),
            .in3(N__10860),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_0_ac0_3_0_a1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_17_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_17_15_6 .LUT_INIT=16'b0011111101111111;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_17_15_6  (
            .in0(N__13381),
            .in1(N__13656),
            .in2(N__9458),
            .in3(N__13577),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_0_ac0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m3_0_LC_17_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m3_0_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m3_0_LC_17_15_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_vga_signals.un6_address_if_m3_0_LC_17_15_7  (
            .in0(N__9455),
            .in1(N__9449),
            .in2(N__9443),
            .in3(N__9440),
            .lcout(\this_vga_signals.if_N_4_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_15_LC_17_16_5 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_15_LC_17_16_5 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_15_LC_17_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_15_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9434),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19134),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_17_17_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_17_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__9411),
            .in2(N__9389),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_17_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_17_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_17_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__9365),
            .in2(_gnd_net_),
            .in3(N__9353),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__19142),
            .ce(),
            .sr(N__17798));
    defparam \this_vga_signals.M_hcounter_q_3_LC_17_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_17_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_17_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__9350),
            .in2(_gnd_net_),
            .in3(N__9338),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__19142),
            .ce(),
            .sr(N__17798));
    defparam \this_vga_signals.M_hcounter_q_4_LC_17_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_17_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_17_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__9334),
            .in2(_gnd_net_),
            .in3(N__9320),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__19142),
            .ce(),
            .sr(N__17798));
    defparam \this_vga_signals.M_hcounter_q_5_LC_17_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_17_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_17_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__9317),
            .in2(_gnd_net_),
            .in3(N__9299),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__19142),
            .ce(),
            .sr(N__17798));
    defparam \this_vga_signals.M_hcounter_q_6_LC_17_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_17_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_17_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__9296),
            .in2(_gnd_net_),
            .in3(N__9278),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__19142),
            .ce(),
            .sr(N__17798));
    defparam \this_vga_signals.M_hcounter_q_7_LC_17_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_17_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_17_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_17_17_6  (
            .in0(N__14082),
            .in1(N__9595),
            .in2(_gnd_net_),
            .in3(N__9575),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__19142),
            .ce(),
            .sr(N__17798));
    defparam \this_vga_signals.M_hcounter_q_8_LC_17_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_17_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__9571),
            .in2(_gnd_net_),
            .in3(N__9551),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__19142),
            .ce(),
            .sr(N__17798));
    defparam \this_vga_signals.M_hcounter_q_9_LC_17_18_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_9_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_9_LC_17_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_9_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__9548),
            .in2(_gnd_net_),
            .in3(N__9527),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_9 ),
            .clk(N__19149),
            .ce(),
            .sr(N__17796));
    defparam \this_vga_signals.M_hcounter_q_10_LC_17_18_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_10_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_10_LC_17_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_10_LC_17_18_1  (
            .in0(N__14093),
            .in1(N__9506),
            .in2(_gnd_net_),
            .in3(N__9488),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_10 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_9 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_10 ),
            .clk(N__19149),
            .ce(),
            .sr(N__17796));
    defparam \this_vga_signals.M_hcounter_q_11_LC_17_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_11_LC_17_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_11_LC_17_18_2 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \this_vga_signals.M_hcounter_q_11_LC_17_18_2  (
            .in0(N__9482),
            .in1(N__14092),
            .in2(_gnd_net_),
            .in3(N__9485),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19149),
            .ce(),
            .sr(N__17796));
    defparam \this_vga_signals.un14_address_g1_1_1_0_LC_18_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_1_1_0_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_1_1_0_LC_18_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un14_address_g1_1_1_0_LC_18_9_0  (
            .in0(N__13895),
            .in1(N__14027),
            .in2(_gnd_net_),
            .in3(N__15348),
            .lcout(\this_vga_signals.g1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g2_1_0_LC_18_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g2_1_0_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g2_1_0_LC_18_9_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un14_address_g2_1_0_LC_18_9_5  (
            .in0(_gnd_net_),
            .in1(N__15105),
            .in2(_gnd_net_),
            .in3(N__16369),
            .lcout(),
            .ltout(\this_vga_signals.g2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g2_3_0_LC_18_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g2_3_0_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g2_3_0_LC_18_9_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un14_address_g2_3_0_LC_18_9_6  (
            .in0(N__13894),
            .in1(N__14505),
            .in2(N__9461),
            .in3(N__15214),
            .lcout(),
            .ltout(\this_vga_signals.g2_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g2_5_LC_18_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g2_5_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g2_5_LC_18_9_7 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \this_vga_signals.un14_address_g2_5_LC_18_9_7  (
            .in0(N__15347),
            .in1(N__12628),
            .in2(N__9638),
            .in3(N__12358),
            .lcout(\this_vga_signals.g2_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_18_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_18_10_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_18_10_0  (
            .in0(N__17724),
            .in1(N__17683),
            .in2(_gnd_net_),
            .in3(N__17638),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_11_LC_18_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_11_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_11_LC_18_10_1 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \this_vga_signals.un14_address_g0_11_LC_18_10_1  (
            .in0(N__12620),
            .in1(N__12455),
            .in2(N__12427),
            .in3(N__12367),
            .lcout(),
            .ltout(\this_vga_signals.if_N_2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_10_LC_18_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_10_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_10_LC_18_10_2 .LUT_INIT=16'b0101010111101000;
    LogicCell40 \this_vga_signals.un14_address_g0_10_LC_18_10_2  (
            .in0(N__14500),
            .in1(N__13958),
            .in2(N__9635),
            .in3(N__10343),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_0_6_LC_18_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_0_6_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_0_6_LC_18_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un14_address_g0_0_6_LC_18_10_3  (
            .in0(N__17639),
            .in1(N__10280),
            .in2(N__9632),
            .in3(N__10289),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_1_0_LC_18_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_1_0_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_1_0_LC_18_10_4 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \this_vga_signals.un14_address_g0_1_0_LC_18_10_4  (
            .in0(N__14036),
            .in1(N__13959),
            .in2(N__9629),
            .in3(N__9626),
            .lcout(\this_vga_signals.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m5_1_LC_18_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m5_1_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m5_1_LC_18_10_5 .LUT_INIT=16'b0111011001100100;
    LogicCell40 \this_vga_signals.un14_address_if_m5_1_LC_18_10_5  (
            .in0(N__14503),
            .in1(N__10734),
            .in2(N__13974),
            .in3(N__10349),
            .lcout(\this_vga_signals.mult1_un61_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un68_sum_axb2_LC_18_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un68_sum_axb2_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un68_sum_axb2_LC_18_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un68_sum_axb2_LC_18_10_6  (
            .in0(N__17725),
            .in1(N__13960),
            .in2(N__9614),
            .in3(N__14504),
            .lcout(\this_vga_signals.mult1_un68_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_14_N_4L6_LC_18_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_14_N_4L6_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_14_N_4L6_LC_18_10_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un14_address_g0_14_N_4L6_LC_18_10_7  (
            .in0(N__15111),
            .in1(N__16370),
            .in2(N__13973),
            .in3(N__15215),
            .lcout(\this_vga_signals.g0_14_N_4L6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_2_LC_18_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_2_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_2_LC_18_11_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \this_vga_signals.un14_address_g1_2_LC_18_11_0  (
            .in0(N__10265),
            .in1(N__9704),
            .in2(N__9695),
            .in3(N__10775),
            .lcout(\this_vga_signals.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_RNI85LKP4_2_LC_18_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_RNI85LKP4_2_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_RNI85LKP4_2_LC_18_11_1 .LUT_INIT=16'b1000011111100001;
    LogicCell40 \this_vga_signals.M_vaddress_q_RNI85LKP4_2_LC_18_11_1  (
            .in0(N__17644),
            .in1(N__13965),
            .in2(N__10325),
            .in3(N__14498),
            .lcout(\this_vga_signals.M_vaddress_q_RNI85LKP4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_30_LC_18_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_30_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_30_LC_18_11_2 .LUT_INIT=16'b0011110001101001;
    LogicCell40 \this_vga_signals.un14_address_g0_30_LC_18_11_2  (
            .in0(N__12629),
            .in1(N__15351),
            .in2(N__15125),
            .in3(N__12348),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_33_LC_18_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_33_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_33_LC_18_11_3 .LUT_INIT=16'b0101100001011110;
    LogicCell40 \this_vga_signals.un14_address_g0_33_LC_18_11_3  (
            .in0(N__14506),
            .in1(N__13964),
            .in2(N__9677),
            .in3(N__10760),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_32_LC_18_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_32_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_32_LC_18_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un14_address_g0_32_LC_18_11_4  (
            .in0(N__9656),
            .in1(N__11015),
            .in2(N__9674),
            .in3(N__17643),
            .lcout(),
            .ltout(\this_vga_signals.g3_0_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_17_LC_18_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_17_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_17_LC_18_11_5 .LUT_INIT=16'b1111111100011001;
    LogicCell40 \this_vga_signals.un14_address_g0_17_LC_18_11_5  (
            .in0(N__13975),
            .in1(N__9650),
            .in2(N__9671),
            .in3(N__9668),
            .lcout(\this_vga_signals.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_29_LC_18_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_29_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_29_LC_18_11_7 .LUT_INIT=16'b1000010010101101;
    LogicCell40 \this_vga_signals.un14_address_g0_29_LC_18_11_7  (
            .in0(N__15350),
            .in1(N__14497),
            .in2(N__10769),
            .in3(N__15117),
            .lcout(\this_vga_signals.g1_0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_0_x2_LC_18_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_0_x2_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_0_x2_LC_18_12_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un14_address_g0_0_x2_LC_18_12_1  (
            .in0(N__17654),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14499),
            .lcout(\this_vga_signals.N_4_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_14_N_7L14_1_LC_18_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_14_N_7L14_1_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_14_N_7L14_1_LC_18_12_3 .LUT_INIT=16'b0010101100110001;
    LogicCell40 \this_vga_signals.un14_address_g0_14_N_7L14_1_LC_18_12_3  (
            .in0(N__15112),
            .in1(N__10331),
            .in2(N__14516),
            .in3(N__15349),
            .lcout(\this_vga_signals.g0_14_N_7L14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m2_0_1_LC_18_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m2_0_1_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m2_0_1_LC_18_12_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un6_address_if_m2_0_1_LC_18_12_4  (
            .in0(N__10702),
            .in1(N__9874),
            .in2(_gnd_net_),
            .in3(N__10883),
            .lcout(\this_vga_signals.if_m2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m2_0_LC_18_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m2_0_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m2_0_LC_18_13_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un6_address_if_m2_0_LC_18_13_0  (
            .in0(N__9755),
            .in1(N__19849),
            .in2(N__11701),
            .in3(N__9710),
            .lcout(\this_vga_signals.if_N_3_0_i ),
            .ltout(\this_vga_signals.if_N_3_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m4_LC_18_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m4_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m4_LC_18_13_1 .LUT_INIT=16'b0010010110000101;
    LogicCell40 \this_vga_signals.un6_address_if_m4_LC_18_13_1  (
            .in0(N__11374),
            .in1(N__9839),
            .in2(N__9743),
            .in3(N__11413),
            .lcout(\this_vga_signals.mult1_un75_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m7_0_x4_LC_18_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m7_0_x4_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m7_0_x4_LC_18_13_2 .LUT_INIT=16'b0011011010010011;
    LogicCell40 \this_vga_signals.un6_address_if_m7_0_x4_LC_18_13_2  (
            .in0(N__10882),
            .in1(N__10387),
            .in2(N__9940),
            .in3(N__10575),
            .lcout(\this_vga_signals.if_N_8_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_18_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_18_13_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_18_13_3  (
            .in0(N__10701),
            .in1(N__9734),
            .in2(N__10388),
            .in3(N__10522),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_3_1_LC_18_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_3_1_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_3_1_LC_18_13_4 .LUT_INIT=16'b0001011111010100;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_3_1_LC_18_13_4  (
            .in0(N__10524),
            .in1(N__10001),
            .in2(N__9941),
            .in3(N__10547),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_haddress_q_RNILVKM8_6_LC_18_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_haddress_q_RNILVKM8_6_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_haddress_q_RNILVKM8_6_LC_18_13_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.M_haddress_q_RNILVKM8_6_LC_18_13_5  (
            .in0(N__10576),
            .in1(N__9933),
            .in2(_gnd_net_),
            .in3(N__10881),
            .lcout(),
            .ltout(\this_vga_signals.M_haddress_q_RNILVKM8Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_ac0_3_LC_18_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_ac0_3_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_ac0_3_LC_18_13_6 .LUT_INIT=16'b1000101101000111;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_ac0_3_LC_18_13_6  (
            .in0(N__10523),
            .in1(N__9728),
            .in2(N__9722),
            .in3(N__10546),
            .lcout(\this_vga_signals.mult1_un54_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_18_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_18_13_7 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9719),
            .in3(N__10174),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_1_0_LC_18_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_1_0_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_1_0_LC_18_14_0 .LUT_INIT=16'b0101010110110010;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_1_0_LC_18_14_0  (
            .in0(N__9991),
            .in1(N__9716),
            .in2(N__11698),
            .in3(N__9848),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_1_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_18_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_18_14_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_18_14_1  (
            .in0(N__10706),
            .in1(N__9878),
            .in2(N__9863),
            .in3(N__10867),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m3_2_ns_LC_18_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m3_2_ns_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m3_2_ns_LC_18_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vga_signals.un6_address_if_m3_2_ns_LC_18_14_2  (
            .in0(N__10367),
            .in1(N__9860),
            .in2(_gnd_net_),
            .in3(N__10889),
            .lcout(this_vga_signals_un6_address_if_N_5_mux_0),
            .ltout(this_vga_signals_un6_address_if_N_5_mux_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_ac0_3_LC_18_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_ac0_3_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_ac0_3_LC_18_14_3 .LUT_INIT=16'b1100100011101100;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_ac0_3_LC_18_14_3  (
            .in0(N__9920),
            .in1(N__10383),
            .in2(N__9854),
            .in3(N__10866),
            .lcout(\this_vga_signals.mult1_un47_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m1_LC_18_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m1_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m1_LC_18_14_4 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un6_address_if_m1_LC_18_14_4  (
            .in0(N__10544),
            .in1(_gnd_net_),
            .in2(N__9851),
            .in3(N__9921),
            .lcout(\this_vga_signals.if_m1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axb1_LC_18_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axb1_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axb1_LC_18_14_5 .LUT_INIT=16'b0100001110010100;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axb1_LC_18_14_5  (
            .in0(N__13673),
            .in1(N__13595),
            .in2(N__13515),
            .in3(N__13404),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_18_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_18_14_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_18_14_6  (
            .in0(N__10545),
            .in1(N__9922),
            .in2(N__10005),
            .in3(N__10525),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_0 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_m1_9_1_LC_18_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_m1_9_1_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_m1_9_1_LC_18_14_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un6_address_if_m1_9_1_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9842),
            .in3(N__9995),
            .lcout(\this_vga_signals.if_m1_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_haddress_q_0_LC_18_15_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_0_LC_18_15_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_0_LC_18_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_0_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__9767),
            .in2(N__9831),
            .in3(N__9823),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_0 ),
            .clk(N__19135),
            .ce(),
            .sr(N__10252));
    defparam \this_vga_signals.M_haddress_q_1_LC_18_15_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_1_LC_18_15_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_1_LC_18_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_1_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__9761),
            .in2(_gnd_net_),
            .in3(N__10034),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_haddress_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_1 ),
            .clk(N__19135),
            .ce(),
            .sr(N__10252));
    defparam \this_vga_signals.M_haddress_q_2_LC_18_15_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_2_LC_18_15_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_2_LC_18_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_2_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__10030),
            .in2(_gnd_net_),
            .in3(N__10016),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_haddress_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_2 ),
            .clk(N__19135),
            .ce(),
            .sr(N__10252));
    defparam \this_vga_signals.M_haddress_q_3_LC_18_15_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_3_LC_18_15_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_3_LC_18_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_3_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__11361),
            .in2(_gnd_net_),
            .in3(N__10013),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_haddress_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_3 ),
            .clk(N__19135),
            .ce(),
            .sr(N__10252));
    defparam \this_vga_signals.M_haddress_q_4_LC_18_15_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_4_LC_18_15_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_4_LC_18_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_4_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__11678),
            .in2(_gnd_net_),
            .in3(N__10010),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_haddress_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_4 ),
            .clk(N__19135),
            .ce(),
            .sr(N__10252));
    defparam \this_vga_signals.M_haddress_q_5_LC_18_15_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_5_LC_18_15_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_5_LC_18_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_5_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__9999),
            .in2(_gnd_net_),
            .in3(N__9944),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_haddress_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_5 ),
            .clk(N__19135),
            .ce(),
            .sr(N__10252));
    defparam \this_vga_signals.M_haddress_q_6_LC_18_15_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_6_LC_18_15_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_6_LC_18_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_6_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__9932),
            .in2(_gnd_net_),
            .in3(N__9890),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_haddress_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_6 ),
            .clk(N__19135),
            .ce(),
            .sr(N__10252));
    defparam \this_vga_signals.M_haddress_q_7_LC_18_15_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_7_LC_18_15_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_7_LC_18_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_7_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__10878),
            .in2(_gnd_net_),
            .in3(N__9887),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_haddress_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_7 ),
            .clk(N__19135),
            .ce(),
            .sr(N__10252));
    defparam \this_vga_signals.M_haddress_q_8_LC_18_16_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_8_LC_18_16_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_8_LC_18_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_8_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__13591),
            .in2(_gnd_net_),
            .in3(N__9884),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_8 ),
            .clk(N__19143),
            .ce(),
            .sr(N__10253));
    defparam \this_vga_signals.M_haddress_q_9_LC_18_16_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_9_LC_18_16_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_9_LC_18_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_9_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__13669),
            .in2(_gnd_net_),
            .in3(N__9881),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_9 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_haddress_q_cry_8 ),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_9 ),
            .clk(N__19143),
            .ce(),
            .sr(N__10253));
    defparam \this_vga_signals.M_haddress_q_10_LC_18_16_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_haddress_q_10_LC_18_16_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_10_LC_18_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_haddress_q_10_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__13493),
            .in2(_gnd_net_),
            .in3(N__10259),
            .lcout(\this_vga_signals.M_haddress_qZ0Z_10 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_haddress_q_cry_9 ),
            .carryout(\this_vga_signals.un1_M_haddress_q_cry_10 ),
            .clk(N__19143),
            .ce(),
            .sr(N__10253));
    defparam \this_vga_signals.M_haddress_q_11_LC_18_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_haddress_q_11_LC_18_16_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_haddress_q_11_LC_18_16_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_haddress_q_11_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__13398),
            .in2(_gnd_net_),
            .in3(N__10256),
            .lcout(\this_vga_signals.CO0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19143),
            .ce(),
            .sr(N__10253));
    defparam \this_start_address_delay.this_delay.M_pipe_q_17_LC_18_18_4 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_17_LC_18_18_4 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_17_LC_18_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_17_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10226),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19156),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_18_LC_18_18_6 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_18_LC_18_18_6 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_18_LC_18_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_18_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10214),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19156),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_i_3_LC_18_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_i_3_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_i_3_LC_18_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_i_3_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__10208),
            .in2(_gnd_net_),
            .in3(N__10181),
            .lcout(this_vga_signals_un6_address_if_generate_plus_mult1_un54_sum_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m12_bm_LC_19_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m12_bm_LC_19_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m12_bm_LC_19_9_0 .LUT_INIT=16'b0001000001011110;
    LogicCell40 \this_vga_signals.un14_address_if_m12_bm_LC_19_9_0  (
            .in0(N__10745),
            .in1(N__14030),
            .in2(N__10310),
            .in3(N__14476),
            .lcout(\this_vga_signals.if_m12_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m6_0_N_2L1_LC_19_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m6_0_N_2L1_LC_19_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m6_0_N_2L1_LC_19_9_1 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \this_vga_signals.un14_address_if_m6_0_N_2L1_LC_19_9_1  (
            .in0(N__12398),
            .in1(N__12594),
            .in2(_gnd_net_),
            .in3(N__12353),
            .lcout(),
            .ltout(\this_vga_signals.g1_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m6_0_LC_19_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m6_0_LC_19_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m6_0_LC_19_9_2 .LUT_INIT=16'b0100001000100100;
    LogicCell40 \this_vga_signals.un14_address_if_m6_0_LC_19_9_2  (
            .in0(N__14494),
            .in1(N__14028),
            .in2(N__10040),
            .in3(N__12456),
            .lcout(\this_vga_signals.if_N_7 ),
            .ltout(\this_vga_signals.if_N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m8_bm_LC_19_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m8_bm_LC_19_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m8_bm_LC_19_9_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vga_signals.un14_address_if_m8_bm_LC_19_9_3  (
            .in0(_gnd_net_),
            .in1(N__14495),
            .in2(N__10037),
            .in3(N__10743),
            .lcout(\this_vga_signals.if_m8_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m1_3_LC_19_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m1_3_LC_19_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m1_3_LC_19_9_4 .LUT_INIT=16'b1100100100110110;
    LogicCell40 \this_vga_signals.un14_address_if_m1_3_LC_19_9_4  (
            .in0(N__12354),
            .in1(N__12399),
            .in2(N__12623),
            .in3(N__12457),
            .lcout(\this_vga_signals.if_m1_3 ),
            .ltout(\this_vga_signals.if_m1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m8_am_LC_19_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m8_am_LC_19_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m8_am_LC_19_9_5 .LUT_INIT=16'b0011111110110001;
    LogicCell40 \this_vga_signals.un14_address_if_m8_am_LC_19_9_5  (
            .in0(N__14029),
            .in1(N__14496),
            .in2(N__10301),
            .in3(N__10744),
            .lcout(),
            .ltout(\this_vga_signals.if_m8_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m13_ns_1_LC_19_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m13_ns_1_LC_19_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m13_ns_1_LC_19_9_6 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \this_vga_signals.un14_address_if_m13_ns_1_LC_19_9_6  (
            .in0(N__13944),
            .in1(N__17720),
            .in2(N__10298),
            .in3(N__10295),
            .lcout(\this_vga_signals.if_m13_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_3_LC_19_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_3_LC_19_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_3_LC_19_9_7 .LUT_INIT=16'b0111011100010001;
    LogicCell40 \this_vga_signals.un14_address_g1_3_LC_19_9_7  (
            .in0(N__13961),
            .in1(N__14493),
            .in2(_gnd_net_),
            .in3(N__17637),
            .lcout(\this_vga_signals.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_0_2_LC_19_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_0_2_LC_19_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_0_2_LC_19_10_0 .LUT_INIT=16'b0011110001101001;
    LogicCell40 \this_vga_signals.un14_address_g0_0_2_LC_19_10_0  (
            .in0(N__12312),
            .in1(N__11278),
            .in2(N__11294),
            .in3(N__12587),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_0_1_LC_19_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_0_1_LC_19_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_0_1_LC_19_10_1 .LUT_INIT=16'b0000111101111000;
    LogicCell40 \this_vga_signals.un14_address_g0_0_1_LC_19_10_1  (
            .in0(N__14492),
            .in1(N__10342),
            .in2(N__10283),
            .in3(N__11194),
            .lcout(\this_vga_signals.g0_0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_1_1_LC_19_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_1_1_LC_19_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_1_1_LC_19_10_2 .LUT_INIT=16'b1100110010011001;
    LogicCell40 \this_vga_signals.un14_address_g1_1_1_LC_19_10_2  (
            .in0(N__12311),
            .in1(N__12738),
            .in2(_gnd_net_),
            .in3(N__12586),
            .lcout(\this_vga_signals.g3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_39_LC_19_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_39_LC_19_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_39_LC_19_10_3 .LUT_INIT=16'b0100101001011110;
    LogicCell40 \this_vga_signals.un14_address_g0_39_LC_19_10_3  (
            .in0(N__11239),
            .in1(N__13962),
            .in2(N__14515),
            .in3(N__11216),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_LC_19_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_LC_19_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_LC_19_10_4 .LUT_INIT=16'b0001010111101010;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_LC_19_10_4  (
            .in0(N__11195),
            .in1(N__10733),
            .in2(N__14509),
            .in3(N__11279),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m5_0_LC_19_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m5_0_LC_19_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m5_0_LC_19_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vga_signals.un14_address_if_m5_0_LC_19_10_5  (
            .in0(N__12737),
            .in1(N__12718),
            .in2(_gnd_net_),
            .in3(N__12699),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m1_LC_19_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m1_LC_19_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m1_LC_19_10_6 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \this_vga_signals.un14_address_if_m1_LC_19_10_6  (
            .in0(N__12309),
            .in1(N__12412),
            .in2(N__10352),
            .in3(N__12585),
            .lcout(\this_vga_signals.if_m1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_19_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_19_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_19_10_7 .LUT_INIT=16'b0011110001101001;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_19_10_7  (
            .in0(N__12584),
            .in1(N__12454),
            .in2(N__12420),
            .in3(N__12310),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_26_LC_19_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_26_LC_19_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_26_LC_19_11_0 .LUT_INIT=16'b0111011001100100;
    LogicCell40 \this_vga_signals.un14_address_g0_26_LC_19_11_0  (
            .in0(N__14477),
            .in1(N__10732),
            .in2(N__13972),
            .in3(N__11201),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_12_LC_19_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_12_LC_19_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_12_LC_19_11_1 .LUT_INIT=16'b0011011011001001;
    LogicCell40 \this_vga_signals.un14_address_g0_12_LC_19_11_1  (
            .in0(N__12315),
            .in1(N__15090),
            .in2(N__12605),
            .in3(N__15328),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_N_2L1_LC_19_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_N_2L1_LC_19_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_N_2L1_LC_19_11_2 .LUT_INIT=16'b0000000001100101;
    LogicCell40 \this_vga_signals.un14_address_g1_N_2L1_LC_19_11_2  (
            .in0(N__15089),
            .in1(N__12559),
            .in2(N__14510),
            .in3(N__12314),
            .lcout(\this_vga_signals.g1_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_RNI8GTIA1_4_LC_19_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_RNI8GTIA1_4_LC_19_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_RNI8GTIA1_4_LC_19_11_3 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \this_vga_signals.M_vaddress_q_RNI8GTIA1_4_LC_19_11_3  (
            .in0(N__12316),
            .in1(N__15329),
            .in2(N__15120),
            .in3(N__12598),
            .lcout(\this_vga_signals.G_5_0_x2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axb1_LC_19_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axb1_LC_19_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axb1_LC_19_11_4 .LUT_INIT=16'b0001111011100001;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axb1_LC_19_11_4  (
            .in0(N__12288),
            .in1(N__12558),
            .in2(N__15119),
            .in3(N__15322),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g2_3_LC_19_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g2_3_LC_19_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g2_3_LC_19_11_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.un14_address_g2_3_LC_19_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10316),
            .in3(N__14481),
            .lcout(),
            .ltout(\this_vga_signals.g2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_0_1_LC_19_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_0_1_LC_19_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_0_1_LC_19_11_6 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un14_address_g1_0_1_LC_19_11_6  (
            .in0(N__13948),
            .in1(N__11277),
            .in2(N__10313),
            .in3(N__11193),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_0_0_LC_19_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_0_0_LC_19_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_0_0_LC_19_11_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.un14_address_g0_0_0_LC_19_11_7  (
            .in0(N__14032),
            .in1(N__17636),
            .in2(N__10784),
            .in3(N__10781),
            .lcout(\this_vga_signals.g0_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_29_1_LC_19_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_29_1_LC_19_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_29_1_LC_19_12_0 .LUT_INIT=16'b0001000000100011;
    LogicCell40 \this_vga_signals.un14_address_g0_29_1_LC_19_12_0  (
            .in0(N__12607),
            .in1(N__12317),
            .in2(N__14511),
            .in3(N__15093),
            .lcout(\this_vga_signals.g0_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_34_LC_19_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_34_LC_19_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_34_LC_19_12_3 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \this_vga_signals.un14_address_g0_34_LC_19_12_3  (
            .in0(N__12318),
            .in1(N__11501),
            .in2(N__11252),
            .in3(N__12608),
            .lcout(\this_vga_signals.N_3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m12_am_LC_19_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m12_am_LC_19_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m12_am_LC_19_12_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \this_vga_signals.un14_address_if_m12_am_LC_19_12_5  (
            .in0(N__14475),
            .in1(N__10754),
            .in2(_gnd_net_),
            .in3(N__10742),
            .lcout(\this_vga_signals.if_m12_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_2_LC_19_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_2_LC_19_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_2_LC_19_13_2 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_2_LC_19_13_2  (
            .in0(N__10912),
            .in1(N__10369),
            .in2(_gnd_net_),
            .in3(N__10927),
            .lcout(\this_vga_signals.mult1_un40_sum_m_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_19_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_19_13_4 .LUT_INIT=16'b0101111010100001;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_19_13_4  (
            .in0(N__10928),
            .in1(N__10370),
            .in2(N__10916),
            .in3(N__10579),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_0 ),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_i_3_LC_19_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_i_3_LC_19_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_i_3_LC_19_13_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_i_3_LC_19_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10529),
            .in3(N__10526),
            .lcout(this_vga_signals_un6_address_if_generate_plus_mult1_un47_sum_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_1_LC_19_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_1_LC_19_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_1_LC_19_13_6 .LUT_INIT=16'b0001110111100010;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_1_LC_19_13_6  (
            .in0(N__10940),
            .in1(N__10368),
            .in2(N__12833),
            .in3(N__10880),
            .lcout(\this_vga_signals.mult1_un40_sum_m_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_haddress_q_RNID85Q_11_LC_19_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_haddress_q_RNID85Q_11_LC_19_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_haddress_q_RNID85Q_11_LC_19_14_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_haddress_q_RNID85Q_11_LC_19_14_1  (
            .in0(_gnd_net_),
            .in1(N__13497),
            .in2(_gnd_net_),
            .in3(N__13402),
            .lcout(\this_vga_signals.CO1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_c2_LC_19_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_c2_LC_19_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_c2_LC_19_14_2 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_c2_LC_19_14_2  (
            .in0(N__10939),
            .in1(N__11003),
            .in2(_gnd_net_),
            .in3(N__10862),
            .lcout(\this_vga_signals.mult1_un40_sum_1_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc2_0_LC_19_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc2_0_LC_19_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc2_0_LC_19_14_6 .LUT_INIT=16'b1110011110011100;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc2_0_LC_19_14_6  (
            .in0(N__13403),
            .in1(N__13677),
            .in2(N__13514),
            .in3(N__13599),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axbxc2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_LC_19_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_LC_19_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_LC_19_15_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_LC_19_15_0  (
            .in0(N__13651),
            .in1(N__13573),
            .in2(_gnd_net_),
            .in3(N__13382),
            .lcout(),
            .ltout(\this_vga_signals.N_2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_0_LC_19_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_0_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_0_LC_19_15_1 .LUT_INIT=16'b0000111110101111;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_0_LC_19_15_1  (
            .in0(N__10858),
            .in1(_gnd_net_),
            .in2(N__10904),
            .in3(N__13476),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_LC_19_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_LC_19_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_LC_19_15_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_LC_19_15_2  (
            .in0(N__13652),
            .in1(N__10854),
            .in2(N__13502),
            .in3(N__13385),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_1_axbxc3_a4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_LC_19_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_LC_19_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_LC_19_15_3 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_LC_19_15_3  (
            .in0(N__10859),
            .in1(N__13654),
            .in2(N__10901),
            .in3(N__13580),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_19_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_19_15_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_19_15_4  (
            .in0(N__10790),
            .in1(N__10796),
            .in2(N__10898),
            .in3(N__10895),
            .lcout(\this_vga_signals.mult1_un40_sum1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a5_LC_19_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a5_LC_19_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a5_LC_19_15_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a5_LC_19_15_5  (
            .in0(N__13383),
            .in1(N__13475),
            .in2(N__10879),
            .in3(N__13579),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axbxc3_a5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_1_LC_19_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_1_LC_19_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_1_LC_19_15_6 .LUT_INIT=16'b0000010101000010;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_1_LC_19_15_6  (
            .in0(N__13653),
            .in1(N__13574),
            .in2(N__13501),
            .in3(N__13384),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_ac0_2_LC_19_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_ac0_2_LC_19_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_ac0_2_LC_19_15_7 .LUT_INIT=16'b0000000011100101;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_ac0_2_LC_19_15_7  (
            .in0(N__13386),
            .in1(N__13655),
            .in2(N__13507),
            .in3(N__13581),
            .lcout(\this_vga_signals.mult1_un40_sum_1_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_16_LC_19_16_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_16_LC_19_16_0 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_16_LC_19_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_16_LC_19_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10997),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19150),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_18_LC_19_16_4 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_18_LC_19_16_4 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_18_LC_19_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_18_LC_19_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10973),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19150),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_19_LC_19_16_6 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_19_LC_19_16_6 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_19_LC_19_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_19_LC_19_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10985),
            .lcout(M_this_start_data_delay_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19150),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_17_LC_19_16_7 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_17_LC_19_16_7 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_17_LC_19_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_17_LC_19_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10979),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19150),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0_0_LC_19_17_3 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0_0_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0_0_LC_19_17_3 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0_0_LC_19_17_3  (
            .in0(N__13045),
            .in1(N__19471),
            .in2(_gnd_net_),
            .in3(N__13184),
            .lcout(\this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_5_LC_19_17_4.C_ON=1'b0;
    defparam M_state_q_5_LC_19_17_4.SEQ_MODE=4'b1000;
    defparam M_state_q_5_LC_19_17_4.LUT_INIT=16'b0000111110001111;
    LogicCell40 M_state_q_5_LC_19_17_4 (
            .in0(N__11312),
            .in1(N__13046),
            .in2(N__10961),
            .in3(N__11390),
            .lcout(M_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19157),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o4_5_LC_19_17_6 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o4_5_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o4_5_LC_19_17_6 .LUT_INIT=16'b1111111101010001;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o4_5_LC_19_17_6  (
            .in0(N__17160),
            .in1(N__10967),
            .in2(N__13187),
            .in3(N__19531),
            .lcout(\this_start_data_delay.this_edge_detector.N_252_0 ),
            .ltout(\this_start_data_delay.this_edge_detector.N_252_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0_0_LC_19_17_7 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0_0_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0_0_LC_19_17_7 .LUT_INIT=16'b0111000000110000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0_0_LC_19_17_7  (
            .in0(N__13091),
            .in1(N__10952),
            .in2(N__10943),
            .in3(N__11389),
            .lcout(\this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_19_LC_19_18_1 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_19_LC_19_18_1 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_19_LC_19_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_19_LC_19_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11180),
            .lcout(M_this_start_address_delay_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19162),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a2_0_5_LC_19_18_3 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a2_0_5_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a2_0_5_LC_19_18_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a2_0_5_LC_19_18_3  (
            .in0(N__13185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19511),
            .lcout(\this_start_data_delay.this_edge_detector.N_267 ),
            .ltout(\this_start_data_delay.this_edge_detector.N_267_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_4_LC_19_18_4.C_ON=1'b0;
    defparam M_state_q_4_LC_19_18_4.SEQ_MODE=4'b1000;
    defparam M_state_q_4_LC_19_18_4.LUT_INIT=16'b1100000000000000;
    LogicCell40 M_state_q_4_LC_19_18_4 (
            .in0(_gnd_net_),
            .in1(N__13094),
            .in2(N__11174),
            .in3(N__13062),
            .lcout(debug_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19162),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m13_ns_LC_19_31_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m13_ns_LC_19_31_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m13_ns_LC_19_31_1 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_vga_signals.un14_address_if_m13_ns_LC_19_31_1  (
            .in0(N__11171),
            .in1(N__11156),
            .in2(N__13976),
            .in3(N__11135),
            .lcout(if_m13_ns),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_11_LC_20_8_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_11_LC_20_8_2 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_11_LC_20_8_2 .LUT_INIT=16'b1010101010011001;
    LogicCell40 \this_vram.mem_radreg_11_LC_20_8_2  (
            .in0(N__15346),
            .in1(N__12627),
            .in2(_gnd_net_),
            .in3(N__12355),
            .lcout(\this_vram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19113),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_6_3_i_o3_LC_20_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_6_3_i_o3_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_6_3_i_o3_LC_20_9_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un14_address_g0_6_3_i_o3_LC_20_9_1  (
            .in0(N__15046),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15345),
            .lcout(),
            .ltout(\this_vga_signals.N_9_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_4_2_LC_20_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_4_2_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_4_2_LC_20_9_2 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \this_vga_signals.un14_address_g0_4_2_LC_20_9_2  (
            .in0(N__11972),
            .in1(N__12593),
            .in2(N__11018),
            .in3(N__12352),
            .lcout(\this_vga_signals.g0_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_20_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_20_9_4 .LUT_INIT=16'b0111000110001110;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_20_9_4  (
            .in0(N__15205),
            .in1(N__15045),
            .in2(N__16382),
            .in3(N__11897),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_x_LC_20_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_x_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_x_LC_20_9_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_x_LC_20_9_7  (
            .in0(N__15044),
            .in1(N__16378),
            .in2(_gnd_net_),
            .in3(N__15204),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_x ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_44_LC_20_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_44_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_44_LC_20_10_0 .LUT_INIT=16'b0001111011100001;
    LogicCell40 \this_vga_signals.un14_address_g0_44_LC_20_10_0  (
            .in0(N__12556),
            .in1(N__12285),
            .in2(N__15122),
            .in3(N__15297),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_0_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_20_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_20_10_1 .LUT_INIT=16'b1000000000010000;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_20_10_1  (
            .in0(N__16371),
            .in1(N__12804),
            .in2(N__15118),
            .in3(N__15179),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_d ),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_3_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_37_LC_20_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_37_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_37_LC_20_10_2 .LUT_INIT=16'b1111110000000011;
    LogicCell40 \this_vga_signals.un14_address_g0_37_LC_20_10_2  (
            .in0(_gnd_net_),
            .in1(N__12286),
            .in2(N__11225),
            .in3(N__15298),
            .lcout(),
            .ltout(\this_vga_signals.if_N_2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_36_LC_20_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_36_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_36_LC_20_10_3 .LUT_INIT=16'b1110100001010101;
    LogicCell40 \this_vga_signals.un14_address_g0_36_LC_20_10_3  (
            .in0(N__15082),
            .in1(N__14471),
            .in2(N__11222),
            .in3(N__12026),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_42_LC_20_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_42_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_42_LC_20_10_4 .LUT_INIT=16'b1110000100011110;
    LogicCell40 \this_vga_signals.un14_address_g0_42_LC_20_10_4  (
            .in0(N__12557),
            .in1(N__12287),
            .in2(N__11219),
            .in3(N__11903),
            .lcout(\this_vga_signals.N_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_3_0_LC_20_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_3_0_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_3_0_LC_20_10_5 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \this_vga_signals.un14_address_g0_3_0_LC_20_10_5  (
            .in0(N__12284),
            .in1(N__11210),
            .in2(N__11896),
            .in3(N__12555),
            .lcout(),
            .ltout(\this_vga_signals.g0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_18_LC_20_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_18_LC_20_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_18_LC_20_10_6 .LUT_INIT=16'b0001111011010010;
    LogicCell40 \this_vga_signals.un14_address_g0_18_LC_20_10_6  (
            .in0(N__12739),
            .in1(N__12717),
            .in2(N__11204),
            .in3(N__12700),
            .lcout(\this_vga_signals.if_N_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_ac0_2_LC_20_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_ac0_2_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_ac0_2_LC_20_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_ac0_2_LC_20_11_0  (
            .in0(N__15100),
            .in1(N__15299),
            .in2(_gnd_net_),
            .in3(N__12289),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m2_3_LC_20_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m2_3_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m2_3_LC_20_11_1 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \this_vga_signals.un14_address_if_m2_3_LC_20_11_1  (
            .in0(N__14609),
            .in1(N__16347),
            .in2(_gnd_net_),
            .in3(N__15185),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m1_0_LC_20_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m1_0_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m1_0_LC_20_11_2 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \this_vga_signals.un14_address_if_m1_0_LC_20_11_2  (
            .in0(N__15186),
            .in1(N__12554),
            .in2(N__11297),
            .in3(N__12055),
            .lcout(\this_vga_signals.if_m1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m5_0_s_LC_20_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m5_0_s_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m5_0_s_LC_20_11_3 .LUT_INIT=16'b0001001001001000;
    LogicCell40 \this_vga_signals.un14_address_if_m5_0_s_LC_20_11_3  (
            .in0(N__15083),
            .in1(N__16348),
            .in2(N__14508),
            .in3(N__15188),
            .lcout(\this_vga_signals.if_m5_0_s ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_0_4_LC_20_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_0_4_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_0_4_LC_20_11_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un14_address_g0_0_4_LC_20_11_4  (
            .in0(_gnd_net_),
            .in1(N__15085),
            .in2(_gnd_net_),
            .in3(N__15301),
            .lcout(\this_vga_signals.g0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_LC_20_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_LC_20_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_LC_20_11_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_LC_20_11_5  (
            .in0(N__15084),
            .in1(N__16349),
            .in2(_gnd_net_),
            .in3(N__15187),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_2_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_0_LC_20_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_0_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_0_LC_20_11_6 .LUT_INIT=16'b0011110001101001;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_0_LC_20_11_6  (
            .in0(N__12563),
            .in1(N__15300),
            .in2(N__11282),
            .in3(N__12290),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_9_LC_20_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_9_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_9_LC_20_11_7 .LUT_INIT=16'b0011110001101001;
    LogicCell40 \this_vga_signals.un14_address_g0_9_LC_20_11_7  (
            .in0(N__12291),
            .in1(N__15101),
            .in2(N__15333),
            .in3(N__12564),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_c2_LC_20_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_c2_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_c2_LC_20_12_3 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_c2_LC_20_12_3  (
            .in0(N__15091),
            .in1(N__16365),
            .in2(_gnd_net_),
            .in3(N__15200),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_3_1_LC_20_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_3_1_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_3_1_LC_20_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un14_address_g0_3_1_LC_20_12_4  (
            .in0(_gnd_net_),
            .in1(N__12809),
            .in2(N__11255),
            .in3(N__12056),
            .lcout(\this_vga_signals.g0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_19_LC_20_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_19_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_19_LC_20_12_5 .LUT_INIT=16'b1010101010011001;
    LogicCell40 \this_vga_signals.un14_address_g0_19_LC_20_12_5  (
            .in0(N__15314),
            .in1(N__12606),
            .in2(_gnd_net_),
            .in3(N__12313),
            .lcout(),
            .ltout(\this_vga_signals.if_N_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_35_LC_20_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_35_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_35_LC_20_12_6 .LUT_INIT=16'b1110100000110011;
    LogicCell40 \this_vga_signals.un14_address_g0_35_LC_20_12_6  (
            .in0(N__14482),
            .in1(N__15092),
            .in2(N__11243),
            .in3(N__11981),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIMTEJ4_11_LC_20_12_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIMTEJ4_11_LC_20_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIMTEJ4_11_LC_20_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_radreg_RNIMTEJ4_11_LC_20_12_7  (
            .in0(N__16187),
            .in1(N__15628),
            .in2(_gnd_net_),
            .in3(N__16778),
            .lcout(M_this_vram_read_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_20_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_20_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_20_14_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_20_14_2  (
            .in0(N__11438),
            .in1(N__11414),
            .in2(_gnd_net_),
            .in3(N__19908),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o3_5_LC_20_17_3 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o3_5_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o3_5_LC_20_17_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o3_5_LC_20_17_3  (
            .in0(_gnd_net_),
            .in1(N__12645),
            .in2(_gnd_net_),
            .in3(N__13208),
            .lcout(\this_start_data_delay.this_edge_detector.N_253_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_1_3_LC_20_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_1_3_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_1_3_LC_20_17_4 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_1_3_LC_20_17_4  (
            .in0(N__11700),
            .in1(N__19915),
            .in2(N__11378),
            .in3(N__19864),
            .lcout(\this_vga_signals.mult1_un68_sum_i_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_2_LC_20_17_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_2_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_2_LC_20_17_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_2_LC_20_17_5  (
            .in0(N__11849),
            .in1(N__11862),
            .in2(N__11812),
            .in3(N__11764),
            .lcout(),
            .ltout(\this_start_data_delay.this_edge_detector.N_261_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_2_LC_20_17_6.C_ON=1'b0;
    defparam M_state_q_2_LC_20_17_6.SEQ_MODE=4'b1000;
    defparam M_state_q_2_LC_20_17_6.LUT_INIT=16'b1111000011110010;
    LogicCell40 M_state_q_2_LC_20_17_6 (
            .in0(N__12646),
            .in1(N__13052),
            .in2(N__11327),
            .in3(N__19472),
            .lcout(M_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19163),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_0_LC_20_17_7.C_ON=1'b0;
    defparam M_state_q_0_LC_20_17_7.SEQ_MODE=4'b1000;
    defparam M_state_q_0_LC_20_17_7.LUT_INIT=16'b1000000011001100;
    LogicCell40 M_state_q_0_LC_20_17_7 (
            .in0(N__11848),
            .in1(N__11324),
            .in2(N__11811),
            .in3(N__11765),
            .lcout(M_state_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19163),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_0_LC_20_18_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_0_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_0_LC_20_18_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_0_LC_20_18_1  (
            .in0(N__14222),
            .in1(N__11318),
            .in2(N__18848),
            .in3(N__11311),
            .lcout(\this_start_data_delay.this_edge_detector.N_275 ),
            .ltout(\this_start_data_delay.this_edge_detector.N_275_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_1_LC_20_18_2 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_1_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_1_LC_20_18_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_1_LC_20_18_2  (
            .in0(N__11841),
            .in1(N__11807),
            .in2(N__11300),
            .in3(N__11863),
            .lcout(),
            .ltout(\this_start_data_delay.this_edge_detector.N_263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_1_LC_20_18_3.C_ON=1'b0;
    defparam M_state_q_1_LC_20_18_3.SEQ_MODE=4'b1000;
    defparam M_state_q_1_LC_20_18_3.LUT_INIT=16'b1111000011110100;
    LogicCell40 M_state_q_1_LC_20_18_3 (
            .in0(N__13063),
            .in1(N__13213),
            .in2(N__11867),
            .in3(N__19519),
            .lcout(M_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19165),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_3_LC_20_18_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_3_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_3_LC_20_18_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_3_LC_20_18_5  (
            .in0(N__11864),
            .in1(N__11842),
            .in2(N__11813),
            .in3(N__11763),
            .lcout(),
            .ltout(\this_start_data_delay.this_edge_detector.N_259_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_3_LC_20_18_6.C_ON=1'b0;
    defparam M_state_q_3_LC_20_18_6.SEQ_MODE=4'b1000;
    defparam M_state_q_3_LC_20_18_6.LUT_INIT=16'b1111000011110100;
    LogicCell40 M_state_q_3_LC_20_18_6 (
            .in0(N__19518),
            .in1(N__13092),
            .in2(N__11750),
            .in3(N__13064),
            .lcout(M_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19165),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_3_LC_20_31_1 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_3_LC_20_31_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_3_LC_20_31_1 .LUT_INIT=16'b0010101111010100;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_3_LC_20_31_1  (
            .in0(N__11747),
            .in1(N__11726),
            .in2(N__11714),
            .in3(N__11630),
            .lcout(this_vga_signals_un6_address_if_generate_plus_mult1_un68_sum_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_12_LC_21_9_1 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_12_LC_21_9_1 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_12_LC_21_9_1 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \this_vram.mem_radreg_12_LC_21_9_1  (
            .in0(N__12893),
            .in1(N__11995),
            .in2(_gnd_net_),
            .in3(N__15468),
            .lcout(\this_vram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19118),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_14_N_8L16_sx_LC_21_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_14_N_8L16_sx_LC_21_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_14_N_8L16_sx_LC_21_9_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un14_address_g0_14_N_8L16_sx_LC_21_9_2  (
            .in0(_gnd_net_),
            .in1(N__14051),
            .in2(_gnd_net_),
            .in3(N__14031),
            .lcout(\this_vga_signals.g0_14_N_8L16_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_0_LC_21_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_0_LC_21_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_0_LC_21_9_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_0_LC_21_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12994),
            .in3(N__12065),
            .lcout(\this_vga_signals.N_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_21_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_21_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_21_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_21_9_4  (
            .in0(N__12082),
            .in1(N__12044),
            .in2(_gnd_net_),
            .in3(N__12763),
            .lcout(\this_vga_signals.mult1_un40_sum1_3 ),
            .ltout(\this_vga_signals.mult1_un40_sum1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_4_0_LC_21_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_4_0_LC_21_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_4_0_LC_21_9_5 .LUT_INIT=16'b0110011000111100;
    LogicCell40 \this_vga_signals.un14_address_g0_4_0_LC_21_9_5  (
            .in0(N__12892),
            .in1(N__16356),
            .in2(N__11975),
            .in3(N__15467),
            .lcout(\this_vga_signals.g0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIETEJ4_11_LC_21_9_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIETEJ4_11_LC_21_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIETEJ4_11_LC_21_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_radreg_RNIETEJ4_11_LC_21_9_7  (
            .in0(N__15611),
            .in1(N__16418),
            .in2(_gnd_net_),
            .in3(N__15998),
            .lcout(M_this_vram_read_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_1_1_1_LC_21_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_1_1_1_LC_21_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_1_1_1_LC_21_10_0 .LUT_INIT=16'b0110011000001111;
    LogicCell40 \this_vga_signals.un14_address_g0_1_1_1_LC_21_10_0  (
            .in0(N__12935),
            .in1(N__12920),
            .in2(N__12020),
            .in3(N__15459),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_3_2_LC_21_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_3_2_LC_21_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_3_2_LC_21_10_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un14_address_g0_3_2_LC_21_10_1  (
            .in0(N__14749),
            .in1(N__11873),
            .in2(N__11906),
            .in3(N__12861),
            .lcout(\this_vga_signals.g0_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_1_LC_21_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_1_LC_21_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_1_LC_21_10_2 .LUT_INIT=16'b0011110001011010;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_1_LC_21_10_2  (
            .in0(N__12015),
            .in1(N__12919),
            .in2(N__12808),
            .in3(N__15458),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_1_LC_21_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_1_LC_21_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_1_LC_21_10_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_1_LC_21_10_3  (
            .in0(_gnd_net_),
            .in1(N__14707),
            .in2(_gnd_net_),
            .in3(N__12860),
            .lcout(\this_vga_signals.mult1_un40_sum_m_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_6_LC_21_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_6_LC_21_10_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_6_LC_21_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_6_LC_21_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14593),
            .lcout(\this_vga_signals.M_vaddress_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19124),
            .ce(),
            .sr(N__16240));
    defparam \this_vga_signals.M_vaddress_q_fast_6_LC_21_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_fast_6_LC_21_10_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_fast_6_LC_21_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_fast_6_LC_21_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14594),
            .lcout(\this_vga_signals.M_vaddress_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19124),
            .ce(),
            .sr(N__16240));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_3_LC_21_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_3_LC_21_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_3_LC_21_10_7 .LUT_INIT=16'b1111010011111111;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_3_LC_21_10_7  (
            .in0(N__14831),
            .in1(N__12859),
            .in2(N__12782),
            .in3(N__11879),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_3_2_1_LC_21_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_3_2_1_LC_21_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_3_2_1_LC_21_11_0 .LUT_INIT=16'b0011100110011100;
    LogicCell40 \this_vga_signals.un14_address_g0_3_2_1_LC_21_11_0  (
            .in0(N__16363),
            .in1(N__13706),
            .in2(N__15121),
            .in3(N__15189),
            .lcout(\this_vga_signals.g0_3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_x_2_LC_21_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_x_2_LC_21_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_x_2_LC_21_11_1 .LUT_INIT=16'b0001000110001000;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_x_2_LC_21_11_1  (
            .in0(N__13704),
            .in1(N__14753),
            .in2(_gnd_net_),
            .in3(N__12862),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_m_am_x_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_2_LC_21_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_2_LC_21_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_2_LC_21_11_2 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_2_LC_21_11_2  (
            .in0(N__15456),
            .in1(N__13828),
            .in2(N__12059),
            .in3(N__12917),
            .lcout(\this_vga_signals.mult1_un40_sum_m_ns_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_x1_3_LC_21_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_x1_3_LC_21_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_x1_3_LC_21_11_3 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_x1_3_LC_21_11_3  (
            .in0(N__15454),
            .in1(N__12043),
            .in2(N__12764),
            .in3(N__12881),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_m_x1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_3_LC_21_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_3_LC_21_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_3_LC_21_11_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_3_LC_21_11_4  (
            .in0(N__12882),
            .in1(N__15455),
            .in2(N__12032),
            .in3(N__12083),
            .lcout(\this_vga_signals.mult1_un40_sum_m_ns_3 ),
            .ltout(\this_vga_signals.mult1_un40_sum_m_ns_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_21_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_21_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_21_11_5 .LUT_INIT=16'b1010010111000011;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_21_11_5  (
            .in0(N__12918),
            .in1(N__12019),
            .in2(N__12029),
            .in3(N__15457),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_3_i_o3_LC_21_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_3_i_o3_LC_21_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_3_i_o3_LC_21_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un14_address_g1_3_i_o3_LC_21_11_6  (
            .in0(N__16364),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15190),
            .lcout(\this_vga_signals.N_6_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_2_LC_21_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_2_LC_21_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_2_LC_21_11_7 .LUT_INIT=16'b1110000101111000;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_2_LC_21_11_7  (
            .in0(N__13705),
            .in1(N__14754),
            .in2(N__13829),
            .in3(N__12863),
            .lcout(\this_vga_signals.mult1_un40_sum_m_am_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_28_LC_21_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_28_LC_21_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_28_LC_21_12_0 .LUT_INIT=16'b0011110001011010;
    LogicCell40 \this_vga_signals.un14_address_g0_28_LC_21_12_0  (
            .in0(N__11999),
            .in1(N__12886),
            .in2(N__16377),
            .in3(N__15470),
            .lcout(\this_vga_signals.N_6_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_16_LC_21_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_16_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_16_LC_21_12_2 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \this_vga_signals.un14_address_g0_16_LC_21_12_2  (
            .in0(N__15321),
            .in1(N__12621),
            .in2(N__15113),
            .in3(N__12322),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_8_LC_21_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_8_LC_21_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_8_LC_21_12_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vga_signals.un14_address_g0_8_LC_21_12_5  (
            .in0(N__12740),
            .in1(N__12719),
            .in2(_gnd_net_),
            .in3(N__12701),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_5_LC_21_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_5_LC_21_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_5_LC_21_12_6 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \this_vga_signals.un14_address_g0_5_LC_21_12_6  (
            .in0(N__12416),
            .in1(N__12622),
            .in2(N__12683),
            .in3(N__12323),
            .lcout(),
            .ltout(\this_vga_signals.if_N_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_15_LC_21_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_15_LC_21_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_15_LC_21_12_7 .LUT_INIT=16'b0101010111101000;
    LogicCell40 \this_vga_signals.un14_address_g0_15_LC_21_12_7  (
            .in0(N__14448),
            .in1(N__13932),
            .in2(N__12680),
            .in3(N__12673),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_0_LC_21_17_4 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_0_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_0_LC_21_17_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_0_LC_21_17_4  (
            .in0(N__13065),
            .in1(N__12647),
            .in2(N__13186),
            .in3(N__13209),
            .lcout(M_current_address_qZ1Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_i_3_LC_21_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_i_3_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_i_3_LC_21_19_7 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_i_3_LC_21_19_7  (
            .in0(N__12632),
            .in1(N__12467),
            .in2(N__12431),
            .in3(N__12368),
            .lcout(this_vga_signals_un14_address_if_generate_plus_mult1_un54_sum_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_4_LC_22_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_4_LC_22_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_4_LC_22_9_0 .LUT_INIT=16'b1111111101001111;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_4_LC_22_9_0  (
            .in0(N__13816),
            .in1(N__13748),
            .in2(N__12749),
            .in3(N__14672),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_7_rep1_LC_22_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_7_rep1_LC_22_9_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_7_rep1_LC_22_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_7_rep1_LC_22_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14566),
            .lcout(\this_vga_signals.M_vaddress_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19125),
            .ce(),
            .sr(N__16241));
    defparam \this_vga_signals.M_vaddress_q_fast_7_LC_22_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_fast_7_LC_22_9_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_fast_7_LC_22_9_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vaddress_q_fast_7_LC_22_9_2  (
            .in0(N__14567),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vaddress_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19125),
            .ce(),
            .sr(N__16241));
    defparam \this_vga_signals.M_vaddress_q_fast_9_LC_22_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_fast_9_LC_22_9_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_fast_9_LC_22_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_fast_9_LC_22_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14543),
            .lcout(\this_vga_signals.M_vaddress_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19125),
            .ce(),
            .sr(N__16241));
    defparam \this_vga_signals.M_vaddress_q_7_LC_22_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_7_LC_22_9_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_7_LC_22_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_7_LC_22_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14565),
            .lcout(\this_vga_signals.M_vaddress_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19125),
            .ce(),
            .sr(N__16241));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_axb1_LC_22_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_axb1_LC_22_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_axb1_LC_22_9_7 .LUT_INIT=16'b1100001001101101;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_axb1_LC_22_9_7  (
            .in0(N__13682),
            .in1(N__13604),
            .in2(N__13520),
            .in3(N__13409),
            .lcout(\this_vga_signals.mult1_un40_sum_0_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_fast_RNI08841_0_8_LC_22_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_fast_RNI08841_0_8_LC_22_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_fast_RNI08841_0_8_LC_22_10_0 .LUT_INIT=16'b0110010001100001;
    LogicCell40 \this_vga_signals.M_vaddress_q_fast_RNI08841_0_8_LC_22_10_0  (
            .in0(N__12961),
            .in1(N__12990),
            .in2(N__13761),
            .in3(N__13811),
            .lcout(\this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8 ),
            .ltout(\this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_LC_22_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_LC_22_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_LC_22_10_1 .LUT_INIT=16'b1001011010011001;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_LC_22_10_1  (
            .in0(N__12818),
            .in1(N__13703),
            .in2(N__12812),
            .in3(N__15453),
            .lcout(\this_vga_signals.mult1_un40_sum_m_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_0_LC_22_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_0_LC_22_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_0_LC_22_10_2 .LUT_INIT=16'b0010001000000111;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_0_LC_22_10_2  (
            .in0(N__12778),
            .in1(N__13004),
            .in2(N__12965),
            .in3(N__12989),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_LC_22_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_LC_22_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_LC_22_10_3 .LUT_INIT=16'b1000101011011011;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_LC_22_10_3  (
            .in0(N__13747),
            .in1(N__13810),
            .in2(N__12767),
            .in3(N__15452),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axbxc3_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_fast_RNIHLHA_8_LC_22_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_fast_RNIHLHA_8_LC_22_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_fast_RNIHLHA_8_LC_22_10_4 .LUT_INIT=16'b0000110000001100;
    LogicCell40 \this_vga_signals.M_vaddress_q_fast_RNIHLHA_8_LC_22_10_4  (
            .in0(_gnd_net_),
            .in1(N__12988),
            .in2(N__12964),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.CO1_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_fast_8_LC_22_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_fast_8_LC_22_10_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_fast_8_LC_22_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_fast_8_LC_22_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14528),
            .lcout(\this_vga_signals.M_vaddress_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19128),
            .ce(),
            .sr(N__16238));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_1_0_LC_22_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_1_0_LC_22_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_1_0_LC_22_10_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_1_0_LC_22_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12963),
            .in3(N__13003),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axbxc3_a4_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_fast_5_LC_22_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_fast_5_LC_22_10_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_fast_5_LC_22_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_fast_5_LC_22_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16401),
            .lcout(\this_vga_signals.M_vaddress_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19128),
            .ce(),
            .sr(N__16238));
    defparam \this_vga_signals.M_vaddress_q_fast_RNI08841_8_LC_22_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_fast_RNI08841_8_LC_22_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_fast_RNI08841_8_LC_22_11_0 .LUT_INIT=16'b0011100111000011;
    LogicCell40 \this_vga_signals.M_vaddress_q_fast_RNI08841_8_LC_22_11_0  (
            .in0(N__12995),
            .in1(N__13804),
            .in2(N__13763),
            .in3(N__12962),
            .lcout(\this_vga_signals.N_353_0 ),
            .ltout(\this_vga_signals.N_353_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_bm_2_LC_22_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_bm_2_LC_22_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_bm_2_LC_22_11_1 .LUT_INIT=16'b0001111010000111;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_bm_2_LC_22_11_1  (
            .in0(N__12858),
            .in1(N__12934),
            .in2(N__12923),
            .in3(N__14723),
            .lcout(\this_vga_signals.mult1_un40_sum_m_bm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_6_rep1_LC_22_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_6_rep1_LC_22_11_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_6_rep1_LC_22_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_6_rep1_LC_22_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14592),
            .lcout(\this_vga_signals.M_vaddress_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19136),
            .ce(),
            .sr(N__16236));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_3_LC_22_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_3_LC_22_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_3_LC_22_11_3 .LUT_INIT=16'b1101110011100011;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_3_LC_22_11_3  (
            .in0(N__14800),
            .in1(N__14656),
            .in2(N__13815),
            .in3(N__13752),
            .lcout(\this_vga_signals.mult1_un40_sum_0_axbxc3_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_1_0_LC_22_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_1_0_LC_22_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_1_0_LC_22_11_4 .LUT_INIT=16'b0011000001011100;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_1_0_LC_22_11_4  (
            .in0(N__13809),
            .in1(N__14664),
            .in2(N__13762),
            .in3(N__12857),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_0_axbxc3_5_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_LC_22_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_LC_22_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_LC_22_11_5 .LUT_INIT=16'b1011110100000000;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_LC_22_11_5  (
            .in0(N__14871),
            .in1(N__14828),
            .in2(N__12902),
            .in3(N__12899),
            .lcout(\this_vga_signals.mult1_un40_sum0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_9_LC_22_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_9_LC_22_11_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_9_LC_22_11_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_vaddress_q_9_LC_22_11_6  (
            .in0(_gnd_net_),
            .in1(N__14539),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19136),
            .ce(),
            .sr(N__16236));
    defparam \this_vga_signals.M_vaddress_q_5_rep1_LC_22_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_5_rep1_LC_22_11_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_5_rep1_LC_22_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_5_rep1_LC_22_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16406),
            .lcout(\this_vga_signals.M_vaddress_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19136),
            .ce(),
            .sr(N__16236));
    defparam \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_LC_22_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_LC_22_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_LC_22_12_0 .LUT_INIT=16'b1001011001001011;
    LogicCell40 \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_LC_22_12_0  (
            .in0(N__14825),
            .in1(N__14660),
            .in2(N__13817),
            .in3(N__13760),
            .lcout(\this_vga_signals.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_0_LC_22_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_0_LC_22_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_0_LC_22_12_1 .LUT_INIT=16'b0100110111000011;
    LogicCell40 \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_0_LC_22_12_1  (
            .in0(N__13805),
            .in1(N__14824),
            .in2(N__14671),
            .in3(N__13759),
            .lcout(\this_vga_signals.N_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_RNIA1HT_1_7_LC_22_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_RNIA1HT_1_7_LC_22_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_RNIA1HT_1_7_LC_22_12_3 .LUT_INIT=16'b0011001010001001;
    LogicCell40 \this_vga_signals.M_vaddress_q_RNIA1HT_1_7_LC_22_12_3  (
            .in0(N__14872),
            .in1(N__14826),
            .in2(N__14756),
            .in3(N__14665),
            .lcout(\this_vga_signals.N_355_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_31_LC_22_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_31_LC_22_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_31_LC_22_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un14_address_g0_31_LC_22_12_4  (
            .in0(N__15000),
            .in1(N__16346),
            .in2(_gnd_net_),
            .in3(N__15191),
            .lcout(\this_vga_signals.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_RNIA1HT_0_7_LC_22_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_RNIA1HT_0_7_LC_22_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_RNIA1HT_0_7_LC_22_12_5 .LUT_INIT=16'b0100110010011011;
    LogicCell40 \this_vga_signals.M_vaddress_q_RNIA1HT_0_7_LC_22_12_5  (
            .in0(N__14873),
            .in1(N__14827),
            .in2(N__14755),
            .in3(N__14666),
            .lcout(\this_vga_signals.N_15_0_0 ),
            .ltout(\this_vga_signals.N_15_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_1_N_2L1_LC_22_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_1_N_2L1_LC_22_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_1_N_2L1_LC_22_12_6 .LUT_INIT=16'b0110100101011010;
    LogicCell40 \this_vga_signals.un14_address_g0_1_N_2L1_LC_22_12_6  (
            .in0(N__14765),
            .in1(N__14894),
            .in2(N__13685),
            .in3(N__15469),
            .lcout(\this_vga_signals.g0_1_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_haddress_q_RNI8ARU_11_LC_22_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_haddress_q_RNI8ARU_11_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_haddress_q_RNI8ARU_11_LC_22_16_1 .LUT_INIT=16'b1000111001011000;
    LogicCell40 \this_vga_signals.M_haddress_q_RNI8ARU_11_LC_22_16_1  (
            .in0(N__13678),
            .in1(N__13600),
            .in2(N__13516),
            .in3(N__13405),
            .lcout(M_haddress_q_RNI8ARU_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_RNI4EAV_1_LC_22_17_6.C_ON=1'b0;
    defparam M_state_q_RNI4EAV_1_LC_22_17_6.SEQ_MODE=4'b0000;
    defparam M_state_q_RNI4EAV_1_LC_22_17_6.LUT_INIT=16'b1100111011001100;
    LogicCell40 M_state_q_RNI4EAV_1_LC_22_17_6 (
            .in0(N__13066),
            .in1(N__17816),
            .in2(N__13180),
            .in3(N__13217),
            .lcout(M_current_address_q_0_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_data_d_0_sqmuxa_0_a4_LC_22_18_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_data_d_0_sqmuxa_0_a4_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_data_d_0_sqmuxa_0_a4_LC_22_18_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_data_d_0_sqmuxa_0_a4_LC_22_18_1  (
            .in0(N__13165),
            .in1(N__13093),
            .in2(_gnd_net_),
            .in3(N__13067),
            .lcout(M_current_data_d_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_22_18_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_22_18_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vram.mem_mem_6_0_wclke_3_LC_22_18_2  (
            .in0(N__17348),
            .in1(N__16972),
            .in2(N__17297),
            .in3(N__17178),
            .lcout(\this_vram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3_0_LC_22_21_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3_0_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3_0_LC_22_21_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3_0_LC_22_21_5  (
            .in0(N__14261),
            .in1(N__14249),
            .in2(_gnd_net_),
            .in3(N__14237),
            .lcout(\this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_data_q_1_LC_22_28_3.C_ON=1'b0;
    defparam M_current_data_q_1_LC_22_28_3.SEQ_MODE=4'b1000;
    defparam M_current_data_q_1_LC_22_28_3.LUT_INIT=16'b0000000011100010;
    LogicCell40 M_current_data_q_1_LC_22_28_3 (
            .in0(N__14126),
            .in1(N__19601),
            .in2(N__18032),
            .in3(N__19505),
            .lcout(M_current_data_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19187),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_0_LC_23_9_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vaddress_q_0_LC_23_9_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_0_LC_23_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vaddress_q_0_LC_23_9_0  (
            .in0(_gnd_net_),
            .in1(N__14050),
            .in2(N__14111),
            .in3(N__14110),
            .lcout(\this_vga_signals.M_vaddress_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_23_9_0_),
            .carryout(\this_vga_signals.un1_M_vaddress_q_cry_0 ),
            .clk(N__19129),
            .ce(),
            .sr(N__16239));
    defparam \this_vga_signals.M_vaddress_q_1_LC_23_9_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vaddress_q_1_LC_23_9_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_1_LC_23_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vaddress_q_1_LC_23_9_1  (
            .in0(_gnd_net_),
            .in1(N__14020),
            .in2(_gnd_net_),
            .in3(N__13979),
            .lcout(\this_vga_signals.M_vaddress_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vaddress_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vaddress_q_cry_1 ),
            .clk(N__19129),
            .ce(),
            .sr(N__16239));
    defparam \this_vga_signals.M_vaddress_q_2_LC_23_9_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vaddress_q_2_LC_23_9_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_2_LC_23_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vaddress_q_2_LC_23_9_2  (
            .in0(_gnd_net_),
            .in1(N__13878),
            .in2(_gnd_net_),
            .in3(N__13838),
            .lcout(\this_vga_signals.M_vaddress_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vaddress_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vaddress_q_cry_2 ),
            .clk(N__19129),
            .ce(),
            .sr(N__16239));
    defparam \this_vga_signals.M_vaddress_q_3_LC_23_9_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vaddress_q_3_LC_23_9_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_3_LC_23_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vaddress_q_3_LC_23_9_3  (
            .in0(_gnd_net_),
            .in1(N__14339),
            .in2(_gnd_net_),
            .in3(N__13835),
            .lcout(\this_vga_signals.M_vaddress_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vaddress_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vaddress_q_cry_3 ),
            .clk(N__19129),
            .ce(),
            .sr(N__16239));
    defparam \this_vga_signals.M_vaddress_q_4_LC_23_9_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_vaddress_q_4_LC_23_9_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_4_LC_23_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vaddress_q_4_LC_23_9_4  (
            .in0(_gnd_net_),
            .in1(N__14999),
            .in2(_gnd_net_),
            .in3(N__13832),
            .lcout(\this_vga_signals.M_vaddress_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vaddress_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vaddress_q_cry_4 ),
            .clk(N__19129),
            .ce(),
            .sr(N__16239));
    defparam \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKME_LC_23_9_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKME_LC_23_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKME_LC_23_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKME_LC_23_9_5  (
            .in0(_gnd_net_),
            .in1(N__16345),
            .in2(_gnd_net_),
            .in3(N__14597),
            .lcout(\this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKMEZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vaddress_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vaddress_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNE_LC_23_9_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNE_LC_23_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNE_LC_23_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNE_LC_23_9_6  (
            .in0(_gnd_net_),
            .in1(N__14766),
            .in2(_gnd_net_),
            .in3(N__14570),
            .lcout(\this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNEZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vaddress_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vaddress_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOE_LC_23_9_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOE_LC_23_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOE_LC_23_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOE_LC_23_9_7  (
            .in0(_gnd_net_),
            .in1(N__14870),
            .in2(_gnd_net_),
            .in3(N__14552),
            .lcout(\this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOEZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vaddress_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vaddress_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPE_LC_23_10_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPE_LC_23_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPE_LC_23_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPE_LC_23_10_0  (
            .in0(_gnd_net_),
            .in1(N__14823),
            .in2(_gnd_net_),
            .in3(N__14549),
            .lcout(\this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPEZ0 ),
            .ltout(),
            .carryin(bfn_23_10_0_),
            .carryout(\this_vga_signals.un1_M_vaddress_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01RE_LC_23_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01RE_LC_23_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01RE_LC_23_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01RE_LC_23_10_1  (
            .in0(_gnd_net_),
            .in1(N__14670),
            .in2(_gnd_net_),
            .in3(N__14546),
            .lcout(\this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01REZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_8_LC_23_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_8_LC_23_10_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_8_LC_23_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_8_LC_23_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14527),
            .lcout(\this_vga_signals.M_vaddress_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19137),
            .ce(),
            .sr(N__16237));
    defparam \this_vga_signals.un14_address_g0_i_0_LC_23_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_i_0_LC_23_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_i_0_LC_23_11_0 .LUT_INIT=16'b0001010000101000;
    LogicCell40 \this_vga_signals.un14_address_g0_i_0_LC_23_11_0  (
            .in0(N__16309),
            .in1(N__15001),
            .in2(N__14436),
            .in3(N__15206),
            .lcout(\this_vga_signals.N_1253_0 ),
            .ltout(\this_vga_signals.N_1253_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_1_N_5L7_x1_LC_23_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_1_N_5L7_x1_LC_23_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_1_N_5L7_x1_LC_23_11_1 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un14_address_g0_1_N_5L7_x1_LC_23_11_1  (
            .in0(N__15397),
            .in1(N__15404),
            .in2(N__14288),
            .in3(N__15361),
            .lcout(\this_vga_signals.g0_1_N_5L7_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_RNIHQ4M_7_LC_23_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_RNIHQ4M_7_LC_23_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vaddress_q_RNIHQ4M_7_LC_23_11_2 .LUT_INIT=16'b0110011011011101;
    LogicCell40 \this_vga_signals.M_vaddress_q_RNIHQ4M_7_LC_23_11_2  (
            .in0(N__14876),
            .in1(N__14822),
            .in2(_gnd_net_),
            .in3(N__14669),
            .lcout(),
            .ltout(\this_vga_signals.g1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_2_LC_23_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_2_LC_23_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_2_LC_23_11_3 .LUT_INIT=16'b0111100000011110;
    LogicCell40 \this_vga_signals.un14_address_g0_2_LC_23_11_3  (
            .in0(N__14757),
            .in1(N__16308),
            .in2(N__15488),
            .in3(N__15485),
            .lcout(),
            .ltout(\this_vga_signals.N_3520_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_7_LC_23_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_7_LC_23_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_7_LC_23_11_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \this_vga_signals.un14_address_g0_7_LC_23_11_4  (
            .in0(N__15479),
            .in1(N__14882),
            .in2(N__15473),
            .in3(N__15466),
            .lcout(\this_vga_signals.mult1_un40_sum_0_2 ),
            .ltout(\this_vga_signals.mult1_un40_sum_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_1_N_5L7_x0_LC_23_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_1_N_5L7_x0_LC_23_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_1_N_5L7_x0_LC_23_11_5 .LUT_INIT=16'b0110100101011010;
    LogicCell40 \this_vga_signals.un14_address_g0_1_N_5L7_x0_LC_23_11_5  (
            .in0(N__15398),
            .in1(N__15376),
            .in2(N__15365),
            .in3(N__15362),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_N_5L7_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_1_N_5L7_ns_LC_23_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_1_N_5L7_ns_LC_23_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_1_N_5L7_ns_LC_23_11_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un14_address_g0_1_N_5L7_ns_LC_23_11_6  (
            .in0(_gnd_net_),
            .in1(N__15334),
            .in2(N__15224),
            .in3(N__15221),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_N_5L7_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g0_1_1_0_LC_23_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g0_1_1_0_LC_23_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g0_1_1_0_LC_23_11_7 .LUT_INIT=16'b0111100011100001;
    LogicCell40 \this_vga_signals.un14_address_g0_1_1_0_LC_23_11_7  (
            .in0(N__15207),
            .in1(N__15064),
            .in2(N__14909),
            .in3(N__16310),
            .lcout(\this_vga_signals.g0_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_13_LC_23_12_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_13_LC_23_12_2 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_13_LC_23_12_2 .LUT_INIT=16'b1001000111101000;
    LogicCell40 \this_vram.mem_radreg_13_LC_23_12_2  (
            .in0(N__14668),
            .in1(N__14875),
            .in2(N__14767),
            .in3(N__14830),
            .lcout(\this_vram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19151),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_g1_0_LC_23_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_g1_0_LC_23_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_g1_0_LC_23_12_5 .LUT_INIT=16'b1101110110111011;
    LogicCell40 \this_vga_signals.un14_address_g1_0_LC_23_12_5  (
            .in0(N__16293),
            .in1(N__14758),
            .in2(_gnd_net_),
            .in3(N__14893),
            .lcout(\this_vga_signals.g1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un14_address_if_m6_LC_23_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_m6_LC_23_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_m6_LC_23_12_7 .LUT_INIT=16'b0100001010010100;
    LogicCell40 \this_vga_signals.un14_address_if_m6_LC_23_12_7  (
            .in0(N__14874),
            .in1(N__14829),
            .in2(N__14768),
            .in3(N__14667),
            .lcout(\this_vga_signals.if_i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_13_1 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_13_1  (
            .in0(N__15632),
            .in1(N__16685),
            .in2(_gnd_net_),
            .in3(N__15926),
            .lcout(M_this_vram_read_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_23_17_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_23_17_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vram.mem_mem_4_0_wclke_3_LC_23_17_4  (
            .in0(N__17330),
            .in1(N__16968),
            .in2(N__17284),
            .in3(N__17194),
            .lcout(\this_vram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_RNIBHE21_3_LC_23_17_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_RNIBHE21_3_LC_23_17_7 .SEQ_MODE=4'b0000;
    defparam \this_reset_cond.M_stage_q_RNIBHE21_3_LC_23_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_reset_cond.M_stage_q_RNIBHE21_3_LC_23_17_7  (
            .in0(_gnd_net_),
            .in1(N__15779),
            .in2(_gnd_net_),
            .in3(N__17815),
            .lcout(M_current_address_q_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_esr_0_LC_23_27_7.C_ON=1'b0;
    defparam M_current_address_q_esr_0_LC_23_27_7.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_0_LC_23_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_current_address_q_esr_0_LC_23_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18156),
            .lcout(M_current_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19188),
            .ce(N__18325),
            .sr(N__17792));
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_7_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_7_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_1_0_RNISSK11_LC_24_7_0  (
            .in0(N__16519),
            .in1(N__15662),
            .in2(_gnd_net_),
            .in3(N__15644),
            .lcout(\this_vram.mem_mem_1_0_RNISSKZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5OL72_0_12_LC_24_8_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5OL72_0_12_LC_24_8_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5OL72_0_12_LC_24_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_radreg_RNI5OL72_0_12_LC_24_8_2  (
            .in0(N__16652),
            .in1(N__15638),
            .in2(_gnd_net_),
            .in3(N__16731),
            .lcout(),
            .ltout(\this_vram.mem_N_109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIETEJ4_0_11_LC_24_8_3 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIETEJ4_0_11_LC_24_8_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIETEJ4_0_11_LC_24_8_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vram.mem_radreg_RNIETEJ4_0_11_LC_24_8_3  (
            .in0(N__15621),
            .in1(_gnd_net_),
            .in2(N__15593),
            .in3(N__15494),
            .lcout(M_this_vram_read_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_8_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_8_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_0_0_RNIQOI11_LC_24_8_5  (
            .in0(N__15524),
            .in1(N__15512),
            .in2(_gnd_net_),
            .in3(N__16520),
            .lcout(),
            .ltout(\this_vram.mem_mem_0_0_RNIQOIZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_8_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_8_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_8_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_8_6  (
            .in0(_gnd_net_),
            .in1(N__16034),
            .in2(N__15497),
            .in3(N__16730),
            .lcout(\this_vram.mem_N_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_9_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_9_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vram.mem_mem_2_0_RNIU0N11_LC_24_9_1  (
            .in0(N__16513),
            .in1(_gnd_net_),
            .in2(N__16061),
            .in3(N__16052),
            .lcout(\this_vram.mem_mem_2_0_RNIU0NZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_9_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_9_5  (
            .in0(N__16512),
            .in1(N__16028),
            .in2(_gnd_net_),
            .in3(N__16016),
            .lcout(),
            .ltout(\this_vram.mem_mem_1_0_RNISSK11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5OL72_12_LC_24_9_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5OL72_12_LC_24_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5OL72_12_LC_24_9_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \this_vram.mem_radreg_RNI5OL72_12_LC_24_9_6  (
            .in0(N__16097),
            .in1(_gnd_net_),
            .in2(N__16001),
            .in3(N__16711),
            .lcout(\this_vram.mem_N_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_10_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_0_1_RNISOI11_LC_24_10_0  (
            .in0(N__15989),
            .in1(N__15974),
            .in2(_gnd_net_),
            .in3(N__16506),
            .lcout(\this_vram.mem_mem_0_1_RNISOIZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_10_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_2_1_RNI01N11_LC_24_10_1  (
            .in0(N__16508),
            .in1(N__15962),
            .in2(_gnd_net_),
            .in3(N__15944),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_10_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_10_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_10_2  (
            .in0(_gnd_net_),
            .in1(N__15935),
            .in2(N__15929),
            .in3(N__16733),
            .lcout(\this_vram.mem_N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_10_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_10_4  (
            .in0(N__15917),
            .in1(N__15902),
            .in2(_gnd_net_),
            .in3(N__16507),
            .lcout(\this_vram.mem_mem_2_0_RNIU0N11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_10_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_10_6  (
            .in0(N__15896),
            .in1(N__15884),
            .in2(_gnd_net_),
            .in3(N__16505),
            .lcout(),
            .ltout(\this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI1GH72_12_LC_24_10_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI1GH72_12_LC_24_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI1GH72_12_LC_24_10_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vram.mem_radreg_RNI1GH72_12_LC_24_10_7  (
            .in0(N__16732),
            .in1(_gnd_net_),
            .in2(N__16427),
            .in3(N__16424),
            .lcout(\this_vram.mem_N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vaddress_q_5_LC_24_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vaddress_q_5_LC_24_11_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vaddress_q_5_LC_24_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vaddress_q_5_LC_24_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16405),
            .lcout(\this_vga_signals.M_vaddress_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19152),
            .ce(),
            .sr(N__16235));
    defparam \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_12_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_12_4  (
            .in0(N__16475),
            .in1(N__16214),
            .in2(_gnd_net_),
            .in3(N__16196),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5GH72_12_LC_24_12_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5GH72_12_LC_24_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5GH72_12_LC_24_12_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vram.mem_radreg_RNI5GH72_12_LC_24_12_5  (
            .in0(N__16734),
            .in1(_gnd_net_),
            .in2(N__16190),
            .in3(N__16148),
            .lcout(\this_vram.mem_N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_12_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_12_7  (
            .in0(N__16175),
            .in1(N__16160),
            .in2(_gnd_net_),
            .in3(N__16474),
            .lcout(\this_vram.mem_mem_0_1_RNISOI11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_24_13_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_24_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_24_13_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vram.mem_mem_1_0_wclke_3_LC_24_13_1  (
            .in0(N__17347),
            .in1(N__16973),
            .in2(N__17291),
            .in3(N__17218),
            .lcout(\this_vram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_2  (
            .in0(N__16478),
            .in1(N__16121),
            .in2(_gnd_net_),
            .in3(N__16103),
            .lcout(\this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_13_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_13_3  (
            .in0(N__16088),
            .in1(N__16073),
            .in2(_gnd_net_),
            .in3(N__16476),
            .lcout(),
            .ltout(\this_vram.mem_mem_1_1_RNIUSK11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI9OL72_12_LC_24_13_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI9OL72_12_LC_24_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI9OL72_12_LC_24_13_4 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \this_vram.mem_radreg_RNI9OL72_12_LC_24_13_4  (
            .in0(N__16736),
            .in1(N__16553),
            .in2(N__16781),
            .in3(_gnd_net_),
            .lcout(\this_vram.mem_N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_13_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_1_1_RNIUSK11_LC_24_13_5  (
            .in0(N__16766),
            .in1(N__16751),
            .in2(_gnd_net_),
            .in3(N__16477),
            .lcout(),
            .ltout(\this_vram.mem_mem_1_1_RNIUSKZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_13_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_13_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_13_6  (
            .in0(N__16735),
            .in1(_gnd_net_),
            .in2(N__16688),
            .in3(N__16436),
            .lcout(\this_vram.mem_N_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_13_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_3_0_RNI05P11_LC_24_13_7  (
            .in0(N__16679),
            .in1(N__16667),
            .in2(_gnd_net_),
            .in3(N__16479),
            .lcout(\this_vram.mem_mem_3_0_RNI05PZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_24_14_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_24_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_24_14_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vram.mem_mem_2_0_wclke_3_LC_24_14_0  (
            .in0(N__17345),
            .in1(N__16966),
            .in2(N__17289),
            .in3(N__17214),
            .lcout(\this_vram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_24_14_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_24_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_24_14_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vram.mem_mem_3_0_wclke_3_LC_24_14_2  (
            .in0(N__17346),
            .in1(N__16967),
            .in2(N__17290),
            .in3(N__17215),
            .lcout(\this_vram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_24_14_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_24_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_24_14_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vram.mem_mem_0_0_wclke_3_LC_24_14_4  (
            .in0(N__17344),
            .in1(N__16965),
            .in2(N__17288),
            .in3(N__17213),
            .lcout(\this_vram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_0  (
            .in0(N__16577),
            .in1(N__16559),
            .in2(_gnd_net_),
            .in3(N__16514),
            .lcout(\this_vram.mem_mem_3_1_RNI25P11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6  (
            .in0(N__16544),
            .in1(N__16538),
            .in2(_gnd_net_),
            .in3(N__16515),
            .lcout(\this_vram.mem_mem_3_1_RNI25PZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_esr_13_LC_24_16_7.C_ON=1'b0;
    defparam M_current_address_q_esr_13_LC_24_16_7.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_13_LC_24_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_current_address_q_esr_13_LC_24_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17491),
            .lcout(M_current_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19169),
            .ce(N__17868),
            .sr(N__17808));
    defparam M_current_address_q_esr_6_LC_24_18_7.C_ON=1'b0;
    defparam M_current_address_q_esr_6_LC_24_18_7.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_6_LC_24_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_current_address_q_esr_6_LC_24_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17492),
            .lcout(M_current_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19172),
            .ce(N__18301),
            .sr(N__17807));
    defparam M_current_address_q_esr_12_LC_24_19_7.C_ON=1'b0;
    defparam M_current_address_q_esr_12_LC_24_19_7.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_12_LC_24_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_current_address_q_esr_12_LC_24_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17101),
            .lcout(M_current_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19175),
            .ce(N__17869),
            .sr(N__17806));
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_20_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_20_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vram.mem_mem_5_0_wclke_3_LC_24_20_5  (
            .in0(N__17317),
            .in1(N__16954),
            .in2(N__17292),
            .in3(N__17216),
            .lcout(\this_vram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_20_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_20_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vram.mem_mem_7_0_wclke_3_LC_24_20_7  (
            .in0(N__17318),
            .in1(N__16955),
            .in2(N__17293),
            .in3(N__17217),
            .lcout(\this_vram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_esr_5_LC_24_21_0.C_ON=1'b0;
    defparam M_current_address_q_esr_5_LC_24_21_0.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_5_LC_24_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_current_address_q_esr_5_LC_24_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17108),
            .lcout(M_current_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19178),
            .ce(N__18316),
            .sr(N__17805));
    defparam M_current_address_q_esr_11_LC_24_22_3.C_ON=1'b0;
    defparam M_current_address_q_esr_11_LC_24_22_3.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_11_LC_24_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_current_address_q_esr_11_LC_24_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16916),
            .lcout(M_current_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19179),
            .ce(N__17880),
            .sr(N__17804));
    defparam M_current_address_q_esr_4_LC_24_23_6.C_ON=1'b0;
    defparam M_current_address_q_esr_4_LC_24_23_6.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_4_LC_24_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_current_address_q_esr_4_LC_24_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16912),
            .lcout(M_current_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19182),
            .ce(N__18317),
            .sr(N__17802));
    defparam M_current_address_q_esr_2_LC_24_24_6.C_ON=1'b0;
    defparam M_current_address_q_esr_2_LC_24_24_6.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_2_LC_24_24_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_current_address_q_esr_2_LC_24_24_6 (
            .in0(N__19730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_current_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19183),
            .ce(N__18318),
            .sr(N__17799));
    defparam M_current_address_q_esr_9_LC_24_25_0.C_ON=1'b0;
    defparam M_current_address_q_esr_9_LC_24_25_0.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_9_LC_24_25_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_current_address_q_esr_9_LC_24_25_0 (
            .in0(N__19723),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_current_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19186),
            .ce(N__17881),
            .sr(N__17797));
    defparam M_current_data_q_0_LC_24_26_4.C_ON=1'b0;
    defparam M_current_data_q_0_LC_24_26_4.SEQ_MODE=4'b1000;
    defparam M_current_data_q_0_LC_24_26_4.LUT_INIT=16'b0000000011100010;
    LogicCell40 M_current_data_q_0_LC_24_26_4 (
            .in0(N__18554),
            .in1(N__19609),
            .in2(N__18173),
            .in3(N__19532),
            .lcout(M_current_data_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19189),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_esr_1_LC_24_27_2.C_ON=1'b0;
    defparam M_current_address_q_esr_1_LC_24_27_2.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_1_LC_24_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_current_address_q_esr_1_LC_24_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18021),
            .lcout(M_current_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19193),
            .ce(N__18326),
            .sr(N__17794));
    defparam M_current_address_q_esr_3_LC_24_27_4.C_ON=1'b0;
    defparam M_current_address_q_esr_3_LC_24_27_4.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_3_LC_24_27_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_current_address_q_esr_3_LC_24_27_4 (
            .in0(N__19566),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_current_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19193),
            .ce(N__18326),
            .sr(N__17794));
    defparam M_current_address_q_esr_10_LC_24_28_6.C_ON=1'b0;
    defparam M_current_address_q_esr_10_LC_24_28_6.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_10_LC_24_28_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_current_address_q_esr_10_LC_24_28_6 (
            .in0(N__19571),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_current_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19194),
            .ce(N__17879),
            .sr(N__17793));
    defparam M_current_address_q_esr_7_LC_24_28_7.C_ON=1'b0;
    defparam M_current_address_q_esr_7_LC_24_28_7.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_7_LC_24_28_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_current_address_q_esr_7_LC_24_28_7 (
            .in0(N__18169),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_current_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19194),
            .ce(N__17879),
            .sr(N__17793));
    defparam M_current_address_q_esr_8_LC_24_29_2.C_ON=1'b0;
    defparam M_current_address_q_esr_8_LC_24_29_2.SEQ_MODE=4'b1000;
    defparam M_current_address_q_esr_8_LC_24_29_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_current_address_q_esr_8_LC_24_29_2 (
            .in0(N__18031),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_current_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19197),
            .ce(N__17885),
            .sr(N__17791));
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_i_3_LC_24_30_2 .C_ON=1'b0;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_i_3_LC_24_30_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_i_3_LC_24_30_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_i_3_LC_24_30_2  (
            .in0(N__17738),
            .in1(N__17699),
            .in2(_gnd_net_),
            .in3(N__17672),
            .lcout(this_vga_signals_un14_address_if_generate_plus_mult1_un61_sum_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_24_31_5 .C_ON=1'b0;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_24_31_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_24_31_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_24_31_5  (
            .in0(_gnd_net_),
            .in1(N__19922),
            .in2(_gnd_net_),
            .in3(N__19880),
            .lcout(this_vga_signals_un6_address_if_generate_plus_mult1_un61_sum_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_data_q_2_LC_26_24_1.C_ON=1'b0;
    defparam M_current_data_q_2_LC_26_24_1.SEQ_MODE=4'b1000;
    defparam M_current_data_q_2_LC_26_24_1.LUT_INIT=16'b0000111000000010;
    LogicCell40 M_current_data_q_2_LC_26_24_1 (
            .in0(N__19639),
            .in1(N__19613),
            .in2(N__19523),
            .in3(N__19722),
            .lcout(M_current_data_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19192),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_data_q_3_LC_26_27_6.C_ON=1'b0;
    defparam M_current_data_q_3_LC_26_27_6.SEQ_MODE=4'b1000;
    defparam M_current_data_q_3_LC_26_27_6.LUT_INIT=16'b0000000011100010;
    LogicCell40 M_current_data_q_3_LC_26_27_6 (
            .in0(N__19220),
            .in1(N__19608),
            .in2(N__19570),
            .in3(N__19504),
            .lcout(M_current_data_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19198),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4_0_LC_32_21_4 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4_0_LC_32_21_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4_0_LC_32_21_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4_0_LC_32_21_4  (
            .in0(N__18917),
            .in1(N__18905),
            .in2(N__18884),
            .in3(N__18869),
            .lcout(\this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
