// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 23 2022 02:01:14

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    led,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output [7:0] led;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__34843;
    wire N__34842;
    wire N__34841;
    wire N__34832;
    wire N__34831;
    wire N__34830;
    wire N__34823;
    wire N__34822;
    wire N__34821;
    wire N__34814;
    wire N__34813;
    wire N__34812;
    wire N__34805;
    wire N__34804;
    wire N__34803;
    wire N__34796;
    wire N__34795;
    wire N__34794;
    wire N__34787;
    wire N__34786;
    wire N__34785;
    wire N__34778;
    wire N__34777;
    wire N__34776;
    wire N__34769;
    wire N__34768;
    wire N__34767;
    wire N__34760;
    wire N__34759;
    wire N__34758;
    wire N__34751;
    wire N__34750;
    wire N__34749;
    wire N__34742;
    wire N__34741;
    wire N__34740;
    wire N__34733;
    wire N__34732;
    wire N__34731;
    wire N__34724;
    wire N__34723;
    wire N__34722;
    wire N__34715;
    wire N__34714;
    wire N__34713;
    wire N__34706;
    wire N__34705;
    wire N__34704;
    wire N__34697;
    wire N__34696;
    wire N__34695;
    wire N__34688;
    wire N__34687;
    wire N__34686;
    wire N__34679;
    wire N__34678;
    wire N__34677;
    wire N__34670;
    wire N__34669;
    wire N__34668;
    wire N__34661;
    wire N__34660;
    wire N__34659;
    wire N__34652;
    wire N__34651;
    wire N__34650;
    wire N__34643;
    wire N__34642;
    wire N__34641;
    wire N__34634;
    wire N__34633;
    wire N__34632;
    wire N__34625;
    wire N__34624;
    wire N__34623;
    wire N__34616;
    wire N__34615;
    wire N__34614;
    wire N__34607;
    wire N__34606;
    wire N__34605;
    wire N__34598;
    wire N__34597;
    wire N__34596;
    wire N__34589;
    wire N__34588;
    wire N__34587;
    wire N__34580;
    wire N__34579;
    wire N__34578;
    wire N__34571;
    wire N__34570;
    wire N__34569;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34553;
    wire N__34552;
    wire N__34551;
    wire N__34544;
    wire N__34543;
    wire N__34542;
    wire N__34535;
    wire N__34534;
    wire N__34533;
    wire N__34526;
    wire N__34525;
    wire N__34524;
    wire N__34517;
    wire N__34516;
    wire N__34515;
    wire N__34508;
    wire N__34507;
    wire N__34506;
    wire N__34499;
    wire N__34498;
    wire N__34497;
    wire N__34490;
    wire N__34489;
    wire N__34488;
    wire N__34481;
    wire N__34480;
    wire N__34479;
    wire N__34472;
    wire N__34471;
    wire N__34470;
    wire N__34463;
    wire N__34462;
    wire N__34461;
    wire N__34454;
    wire N__34453;
    wire N__34452;
    wire N__34445;
    wire N__34444;
    wire N__34443;
    wire N__34436;
    wire N__34435;
    wire N__34434;
    wire N__34427;
    wire N__34426;
    wire N__34425;
    wire N__34418;
    wire N__34417;
    wire N__34416;
    wire N__34409;
    wire N__34408;
    wire N__34407;
    wire N__34400;
    wire N__34399;
    wire N__34398;
    wire N__34391;
    wire N__34390;
    wire N__34389;
    wire N__34382;
    wire N__34381;
    wire N__34380;
    wire N__34363;
    wire N__34362;
    wire N__34359;
    wire N__34358;
    wire N__34357;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34347;
    wire N__34344;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34333;
    wire N__34332;
    wire N__34331;
    wire N__34328;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34318;
    wire N__34313;
    wire N__34310;
    wire N__34307;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34274;
    wire N__34271;
    wire N__34266;
    wire N__34261;
    wire N__34258;
    wire N__34251;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34222;
    wire N__34221;
    wire N__34220;
    wire N__34217;
    wire N__34214;
    wire N__34213;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34202;
    wire N__34199;
    wire N__34196;
    wire N__34193;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34155;
    wire N__34152;
    wire N__34151;
    wire N__34150;
    wire N__34145;
    wire N__34144;
    wire N__34141;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34129;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34100;
    wire N__34097;
    wire N__34092;
    wire N__34087;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34059;
    wire N__34058;
    wire N__34057;
    wire N__34054;
    wire N__34051;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34012;
    wire N__34009;
    wire N__34000;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33992;
    wire N__33991;
    wire N__33990;
    wire N__33989;
    wire N__33986;
    wire N__33983;
    wire N__33982;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33971;
    wire N__33970;
    wire N__33967;
    wire N__33966;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33945;
    wire N__33940;
    wire N__33937;
    wire N__33934;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33885;
    wire N__33882;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33837;
    wire N__33836;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33828;
    wire N__33827;
    wire N__33824;
    wire N__33823;
    wire N__33822;
    wire N__33819;
    wire N__33818;
    wire N__33815;
    wire N__33814;
    wire N__33813;
    wire N__33808;
    wire N__33803;
    wire N__33798;
    wire N__33795;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33730;
    wire N__33725;
    wire N__33720;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33704;
    wire N__33697;
    wire N__33694;
    wire N__33693;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33651;
    wire N__33646;
    wire N__33643;
    wire N__33642;
    wire N__33641;
    wire N__33638;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33614;
    wire N__33613;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33582;
    wire N__33579;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33551;
    wire N__33548;
    wire N__33543;
    wire N__33538;
    wire N__33537;
    wire N__33536;
    wire N__33533;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33512;
    wire N__33509;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33497;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33460;
    wire N__33457;
    wire N__33452;
    wire N__33447;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33427;
    wire N__33426;
    wire N__33423;
    wire N__33422;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33412;
    wire N__33407;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33390;
    wire N__33389;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33365;
    wire N__33362;
    wire N__33357;
    wire N__33354;
    wire N__33351;
    wire N__33348;
    wire N__33345;
    wire N__33340;
    wire N__33337;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33329;
    wire N__33328;
    wire N__33327;
    wire N__33326;
    wire N__33323;
    wire N__33320;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33312;
    wire N__33311;
    wire N__33308;
    wire N__33305;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33270;
    wire N__33267;
    wire N__33266;
    wire N__33263;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33248;
    wire N__33245;
    wire N__33242;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33206;
    wire N__33199;
    wire N__33198;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33126;
    wire N__33125;
    wire N__33122;
    wire N__33117;
    wire N__33116;
    wire N__33115;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33049;
    wire N__33046;
    wire N__33045;
    wire N__33044;
    wire N__33043;
    wire N__33040;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33025;
    wire N__33024;
    wire N__33023;
    wire N__33022;
    wire N__33019;
    wire N__33012;
    wire N__33007;
    wire N__33006;
    wire N__33005;
    wire N__33002;
    wire N__33001;
    wire N__32994;
    wire N__32989;
    wire N__32986;
    wire N__32985;
    wire N__32984;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32967;
    wire N__32960;
    wire N__32957;
    wire N__32952;
    wire N__32947;
    wire N__32944;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32931;
    wire N__32930;
    wire N__32929;
    wire N__32926;
    wire N__32925;
    wire N__32924;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32872;
    wire N__32861;
    wire N__32854;
    wire N__32853;
    wire N__32852;
    wire N__32851;
    wire N__32850;
    wire N__32849;
    wire N__32848;
    wire N__32847;
    wire N__32846;
    wire N__32845;
    wire N__32844;
    wire N__32843;
    wire N__32840;
    wire N__32835;
    wire N__32834;
    wire N__32831;
    wire N__32830;
    wire N__32829;
    wire N__32828;
    wire N__32827;
    wire N__32826;
    wire N__32825;
    wire N__32824;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32805;
    wire N__32800;
    wire N__32795;
    wire N__32792;
    wire N__32791;
    wire N__32790;
    wire N__32789;
    wire N__32788;
    wire N__32787;
    wire N__32786;
    wire N__32785;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32777;
    wire N__32776;
    wire N__32775;
    wire N__32774;
    wire N__32773;
    wire N__32772;
    wire N__32771;
    wire N__32770;
    wire N__32765;
    wire N__32762;
    wire N__32761;
    wire N__32760;
    wire N__32759;
    wire N__32758;
    wire N__32757;
    wire N__32756;
    wire N__32755;
    wire N__32754;
    wire N__32753;
    wire N__32752;
    wire N__32751;
    wire N__32750;
    wire N__32747;
    wire N__32746;
    wire N__32743;
    wire N__32740;
    wire N__32735;
    wire N__32732;
    wire N__32727;
    wire N__32724;
    wire N__32723;
    wire N__32716;
    wire N__32713;
    wire N__32710;
    wire N__32707;
    wire N__32704;
    wire N__32699;
    wire N__32696;
    wire N__32691;
    wire N__32688;
    wire N__32685;
    wire N__32682;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32664;
    wire N__32659;
    wire N__32650;
    wire N__32645;
    wire N__32640;
    wire N__32639;
    wire N__32638;
    wire N__32637;
    wire N__32634;
    wire N__32629;
    wire N__32626;
    wire N__32625;
    wire N__32624;
    wire N__32623;
    wire N__32622;
    wire N__32621;
    wire N__32620;
    wire N__32617;
    wire N__32616;
    wire N__32613;
    wire N__32600;
    wire N__32597;
    wire N__32590;
    wire N__32589;
    wire N__32588;
    wire N__32585;
    wire N__32582;
    wire N__32577;
    wire N__32574;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32502;
    wire N__32499;
    wire N__32494;
    wire N__32487;
    wire N__32476;
    wire N__32471;
    wire N__32464;
    wire N__32437;
    wire N__32436;
    wire N__32435;
    wire N__32434;
    wire N__32433;
    wire N__32432;
    wire N__32431;
    wire N__32430;
    wire N__32429;
    wire N__32428;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32393;
    wire N__32392;
    wire N__32391;
    wire N__32390;
    wire N__32389;
    wire N__32388;
    wire N__32387;
    wire N__32386;
    wire N__32385;
    wire N__32384;
    wire N__32383;
    wire N__32382;
    wire N__32381;
    wire N__32380;
    wire N__32379;
    wire N__32378;
    wire N__32377;
    wire N__32376;
    wire N__32375;
    wire N__32374;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32257;
    wire N__32254;
    wire N__32253;
    wire N__32252;
    wire N__32251;
    wire N__32250;
    wire N__32249;
    wire N__32242;
    wire N__32241;
    wire N__32240;
    wire N__32239;
    wire N__32238;
    wire N__32237;
    wire N__32236;
    wire N__32235;
    wire N__32234;
    wire N__32227;
    wire N__32224;
    wire N__32219;
    wire N__32214;
    wire N__32205;
    wire N__32204;
    wire N__32203;
    wire N__32200;
    wire N__32193;
    wire N__32190;
    wire N__32185;
    wire N__32176;
    wire N__32173;
    wire N__32170;
    wire N__32167;
    wire N__32166;
    wire N__32165;
    wire N__32164;
    wire N__32163;
    wire N__32162;
    wire N__32161;
    wire N__32160;
    wire N__32159;
    wire N__32158;
    wire N__32157;
    wire N__32156;
    wire N__32155;
    wire N__32154;
    wire N__32147;
    wire N__32138;
    wire N__32137;
    wire N__32136;
    wire N__32127;
    wire N__32120;
    wire N__32115;
    wire N__32110;
    wire N__32107;
    wire N__32104;
    wire N__32099;
    wire N__32092;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32077;
    wire N__32074;
    wire N__32071;
    wire N__32062;
    wire N__32061;
    wire N__32060;
    wire N__32059;
    wire N__32058;
    wire N__32057;
    wire N__32056;
    wire N__32055;
    wire N__32054;
    wire N__32053;
    wire N__32052;
    wire N__32051;
    wire N__32050;
    wire N__32049;
    wire N__32048;
    wire N__32047;
    wire N__32046;
    wire N__32045;
    wire N__32044;
    wire N__32043;
    wire N__32042;
    wire N__32041;
    wire N__32040;
    wire N__32039;
    wire N__32038;
    wire N__32037;
    wire N__32036;
    wire N__32035;
    wire N__32034;
    wire N__32033;
    wire N__32032;
    wire N__32031;
    wire N__32030;
    wire N__32029;
    wire N__32028;
    wire N__32027;
    wire N__32026;
    wire N__32025;
    wire N__32024;
    wire N__32023;
    wire N__32022;
    wire N__32021;
    wire N__32020;
    wire N__32019;
    wire N__32018;
    wire N__32017;
    wire N__32016;
    wire N__32015;
    wire N__32014;
    wire N__32013;
    wire N__32012;
    wire N__32011;
    wire N__32010;
    wire N__32009;
    wire N__32008;
    wire N__32007;
    wire N__32006;
    wire N__32005;
    wire N__32004;
    wire N__32003;
    wire N__32002;
    wire N__32001;
    wire N__32000;
    wire N__31999;
    wire N__31998;
    wire N__31997;
    wire N__31996;
    wire N__31995;
    wire N__31994;
    wire N__31993;
    wire N__31992;
    wire N__31991;
    wire N__31990;
    wire N__31989;
    wire N__31988;
    wire N__31987;
    wire N__31986;
    wire N__31985;
    wire N__31984;
    wire N__31983;
    wire N__31982;
    wire N__31981;
    wire N__31980;
    wire N__31979;
    wire N__31978;
    wire N__31977;
    wire N__31976;
    wire N__31975;
    wire N__31974;
    wire N__31973;
    wire N__31972;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31968;
    wire N__31967;
    wire N__31966;
    wire N__31965;
    wire N__31964;
    wire N__31963;
    wire N__31962;
    wire N__31961;
    wire N__31960;
    wire N__31959;
    wire N__31958;
    wire N__31957;
    wire N__31956;
    wire N__31955;
    wire N__31954;
    wire N__31953;
    wire N__31952;
    wire N__31951;
    wire N__31950;
    wire N__31949;
    wire N__31948;
    wire N__31947;
    wire N__31946;
    wire N__31945;
    wire N__31944;
    wire N__31943;
    wire N__31942;
    wire N__31941;
    wire N__31940;
    wire N__31939;
    wire N__31938;
    wire N__31937;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31677;
    wire N__31676;
    wire N__31673;
    wire N__31670;
    wire N__31669;
    wire N__31668;
    wire N__31665;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31643;
    wire N__31636;
    wire N__31635;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31615;
    wire N__31612;
    wire N__31611;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31591;
    wire N__31590;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31567;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31552;
    wire N__31549;
    wire N__31546;
    wire N__31545;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31537;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31516;
    wire N__31515;
    wire N__31514;
    wire N__31509;
    wire N__31508;
    wire N__31507;
    wire N__31506;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31490;
    wire N__31487;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31441;
    wire N__31438;
    wire N__31437;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31404;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31368;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31323;
    wire N__31320;
    wire N__31319;
    wire N__31318;
    wire N__31317;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31296;
    wire N__31295;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31267;
    wire N__31258;
    wire N__31255;
    wire N__31254;
    wire N__31253;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31232;
    wire N__31231;
    wire N__31228;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31203;
    wire N__31202;
    wire N__31201;
    wire N__31200;
    wire N__31199;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31171;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31150;
    wire N__31149;
    wire N__31148;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31129;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31117;
    wire N__31116;
    wire N__31115;
    wire N__31108;
    wire N__31107;
    wire N__31104;
    wire N__31103;
    wire N__31102;
    wire N__31101;
    wire N__31100;
    wire N__31097;
    wire N__31094;
    wire N__31091;
    wire N__31088;
    wire N__31083;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31053;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30991;
    wire N__30988;
    wire N__30985;
    wire N__30982;
    wire N__30979;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30971;
    wire N__30966;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30949;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30936;
    wire N__30933;
    wire N__30932;
    wire N__30929;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30891;
    wire N__30888;
    wire N__30887;
    wire N__30884;
    wire N__30883;
    wire N__30880;
    wire N__30877;
    wire N__30874;
    wire N__30871;
    wire N__30862;
    wire N__30861;
    wire N__30860;
    wire N__30859;
    wire N__30858;
    wire N__30857;
    wire N__30856;
    wire N__30853;
    wire N__30852;
    wire N__30849;
    wire N__30848;
    wire N__30847;
    wire N__30844;
    wire N__30843;
    wire N__30842;
    wire N__30841;
    wire N__30840;
    wire N__30839;
    wire N__30838;
    wire N__30835;
    wire N__30828;
    wire N__30823;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30809;
    wire N__30806;
    wire N__30801;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30785;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30760;
    wire N__30757;
    wire N__30756;
    wire N__30755;
    wire N__30754;
    wire N__30745;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30725;
    wire N__30720;
    wire N__30715;
    wire N__30706;
    wire N__30703;
    wire N__30700;
    wire N__30699;
    wire N__30698;
    wire N__30697;
    wire N__30696;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30685;
    wire N__30684;
    wire N__30683;
    wire N__30682;
    wire N__30677;
    wire N__30676;
    wire N__30675;
    wire N__30672;
    wire N__30671;
    wire N__30670;
    wire N__30669;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30648;
    wire N__30645;
    wire N__30640;
    wire N__30637;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30618;
    wire N__30613;
    wire N__30610;
    wire N__30609;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30597;
    wire N__30592;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30578;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30528;
    wire N__30527;
    wire N__30526;
    wire N__30525;
    wire N__30524;
    wire N__30523;
    wire N__30522;
    wire N__30521;
    wire N__30520;
    wire N__30519;
    wire N__30518;
    wire N__30515;
    wire N__30510;
    wire N__30503;
    wire N__30496;
    wire N__30489;
    wire N__30488;
    wire N__30487;
    wire N__30476;
    wire N__30471;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30410;
    wire N__30407;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30364;
    wire N__30363;
    wire N__30362;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30292;
    wire N__30289;
    wire N__30284;
    wire N__30281;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30237;
    wire N__30236;
    wire N__30233;
    wire N__30228;
    wire N__30227;
    wire N__30222;
    wire N__30219;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30195;
    wire N__30194;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30182;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30156;
    wire N__30155;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30145;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30124;
    wire N__30119;
    wire N__30118;
    wire N__30117;
    wire N__30116;
    wire N__30115;
    wire N__30112;
    wire N__30107;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30093;
    wire N__30092;
    wire N__30091;
    wire N__30090;
    wire N__30089;
    wire N__30086;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30078;
    wire N__30077;
    wire N__30076;
    wire N__30075;
    wire N__30074;
    wire N__30073;
    wire N__30072;
    wire N__30071;
    wire N__30066;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30044;
    wire N__30043;
    wire N__30042;
    wire N__30041;
    wire N__30040;
    wire N__30039;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30031;
    wire N__30030;
    wire N__30025;
    wire N__30022;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30014;
    wire N__30013;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30005;
    wire N__30002;
    wire N__30001;
    wire N__29998;
    wire N__29997;
    wire N__29994;
    wire N__29985;
    wire N__29982;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29967;
    wire N__29966;
    wire N__29963;
    wire N__29962;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29948;
    wire N__29947;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29935;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29913;
    wire N__29898;
    wire N__29895;
    wire N__29892;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29848;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29836;
    wire N__29833;
    wire N__29828;
    wire N__29827;
    wire N__29822;
    wire N__29811;
    wire N__29808;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29786;
    wire N__29783;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29751;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29704;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29673;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29646;
    wire N__29645;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29620;
    wire N__29619;
    wire N__29618;
    wire N__29617;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29596;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29586;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29567;
    wire N__29564;
    wire N__29561;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29538;
    wire N__29537;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29521;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29508;
    wire N__29505;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29478;
    wire N__29477;
    wire N__29474;
    wire N__29469;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29448;
    wire N__29447;
    wire N__29444;
    wire N__29439;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29395;
    wire N__29392;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29382;
    wire N__29379;
    wire N__29378;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29356;
    wire N__29355;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29326;
    wire N__29325;
    wire N__29322;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29295;
    wire N__29292;
    wire N__29291;
    wire N__29290;
    wire N__29287;
    wire N__29284;
    wire N__29279;
    wire N__29276;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29238;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29219;
    wire N__29216;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29191;
    wire N__29190;
    wire N__29189;
    wire N__29188;
    wire N__29187;
    wire N__29182;
    wire N__29181;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29164;
    wire N__29163;
    wire N__29162;
    wire N__29161;
    wire N__29160;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29114;
    wire N__29111;
    wire N__29102;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29082;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29021;
    wire N__29020;
    wire N__29017;
    wire N__29012;
    wire N__29009;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28971;
    wire N__28968;
    wire N__28967;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28955;
    wire N__28952;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28877;
    wire N__28876;
    wire N__28871;
    wire N__28866;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28842;
    wire N__28839;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28785;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28749;
    wire N__28748;
    wire N__28745;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28698;
    wire N__28695;
    wire N__28694;
    wire N__28691;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28578;
    wire N__28575;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28561;
    wire N__28560;
    wire N__28559;
    wire N__28556;
    wire N__28551;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28535;
    wire N__28528;
    wire N__28525;
    wire N__28524;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28509;
    wire N__28506;
    wire N__28505;
    wire N__28504;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28483;
    wire N__28482;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28471;
    wire N__28470;
    wire N__28469;
    wire N__28468;
    wire N__28467;
    wire N__28466;
    wire N__28465;
    wire N__28462;
    wire N__28457;
    wire N__28452;
    wire N__28445;
    wire N__28440;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28266;
    wire N__28263;
    wire N__28262;
    wire N__28259;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28238;
    wire N__28233;
    wire N__28228;
    wire N__28227;
    wire N__28226;
    wire N__28223;
    wire N__28222;
    wire N__28221;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28213;
    wire N__28212;
    wire N__28211;
    wire N__28208;
    wire N__28207;
    wire N__28204;
    wire N__28203;
    wire N__28200;
    wire N__28199;
    wire N__28198;
    wire N__28195;
    wire N__28190;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28171;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28163;
    wire N__28162;
    wire N__28161;
    wire N__28160;
    wire N__28157;
    wire N__28150;
    wire N__28145;
    wire N__28140;
    wire N__28137;
    wire N__28132;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28116;
    wire N__28111;
    wire N__28104;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28077;
    wire N__28076;
    wire N__28075;
    wire N__28074;
    wire N__28069;
    wire N__28064;
    wire N__28061;
    wire N__28056;
    wire N__28053;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28041;
    wire N__28040;
    wire N__28037;
    wire N__28036;
    wire N__28035;
    wire N__28032;
    wire N__28031;
    wire N__28028;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28006;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27994;
    wire N__27991;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27961;
    wire N__27960;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27946;
    wire N__27945;
    wire N__27944;
    wire N__27941;
    wire N__27940;
    wire N__27937;
    wire N__27936;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27925;
    wire N__27924;
    wire N__27921;
    wire N__27916;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27902;
    wire N__27899;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27878;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27825;
    wire N__27824;
    wire N__27823;
    wire N__27822;
    wire N__27821;
    wire N__27820;
    wire N__27819;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27805;
    wire N__27804;
    wire N__27803;
    wire N__27802;
    wire N__27801;
    wire N__27800;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27781;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27763;
    wire N__27762;
    wire N__27759;
    wire N__27754;
    wire N__27747;
    wire N__27744;
    wire N__27737;
    wire N__27734;
    wire N__27729;
    wire N__27724;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27676;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27657;
    wire N__27656;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27631;
    wire N__27628;
    wire N__27627;
    wire N__27626;
    wire N__27625;
    wire N__27624;
    wire N__27623;
    wire N__27622;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27611;
    wire N__27608;
    wire N__27607;
    wire N__27604;
    wire N__27603;
    wire N__27600;
    wire N__27599;
    wire N__27598;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27586;
    wire N__27583;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27558;
    wire N__27555;
    wire N__27554;
    wire N__27545;
    wire N__27542;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27518;
    wire N__27511;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27501;
    wire N__27498;
    wire N__27497;
    wire N__27496;
    wire N__27495;
    wire N__27494;
    wire N__27493;
    wire N__27490;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27482;
    wire N__27481;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27461;
    wire N__27460;
    wire N__27459;
    wire N__27454;
    wire N__27453;
    wire N__27452;
    wire N__27451;
    wire N__27450;
    wire N__27445;
    wire N__27442;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27426;
    wire N__27419;
    wire N__27416;
    wire N__27409;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27383;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27351;
    wire N__27348;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27313;
    wire N__27310;
    wire N__27309;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27291;
    wire N__27290;
    wire N__27289;
    wire N__27288;
    wire N__27287;
    wire N__27286;
    wire N__27285;
    wire N__27284;
    wire N__27283;
    wire N__27282;
    wire N__27281;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27235;
    wire N__27232;
    wire N__27231;
    wire N__27228;
    wire N__27227;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27216;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27208;
    wire N__27207;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27195;
    wire N__27190;
    wire N__27185;
    wire N__27182;
    wire N__27169;
    wire N__27168;
    wire N__27167;
    wire N__27162;
    wire N__27161;
    wire N__27160;
    wire N__27159;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27127;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27118;
    wire N__27115;
    wire N__27112;
    wire N__27107;
    wire N__27104;
    wire N__27099;
    wire N__27098;
    wire N__27097;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27087;
    wire N__27086;
    wire N__27083;
    wire N__27080;
    wire N__27075;
    wire N__27070;
    wire N__27065;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27051;
    wire N__27046;
    wire N__27045;
    wire N__27044;
    wire N__27043;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27031;
    wire N__27030;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27018;
    wire N__27013;
    wire N__27004;
    wire N__27003;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26995;
    wire N__26992;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26978;
    wire N__26975;
    wire N__26974;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26953;
    wire N__26948;
    wire N__26947;
    wire N__26944;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26900;
    wire N__26895;
    wire N__26890;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26882;
    wire N__26879;
    wire N__26878;
    wire N__26877;
    wire N__26874;
    wire N__26873;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26856;
    wire N__26853;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26826;
    wire N__26823;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26807;
    wire N__26800;
    wire N__26797;
    wire N__26796;
    wire N__26793;
    wire N__26792;
    wire N__26791;
    wire N__26790;
    wire N__26787;
    wire N__26786;
    wire N__26783;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26769;
    wire N__26766;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26737;
    wire N__26734;
    wire N__26733;
    wire N__26732;
    wire N__26725;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26717;
    wire N__26716;
    wire N__26715;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26696;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26628;
    wire N__26627;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26574;
    wire N__26573;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26499;
    wire N__26498;
    wire N__26497;
    wire N__26494;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26476;
    wire N__26475;
    wire N__26474;
    wire N__26473;
    wire N__26472;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26464;
    wire N__26463;
    wire N__26462;
    wire N__26459;
    wire N__26454;
    wire N__26453;
    wire N__26450;
    wire N__26445;
    wire N__26442;
    wire N__26437;
    wire N__26436;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26426;
    wire N__26425;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26404;
    wire N__26401;
    wire N__26400;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26386;
    wire N__26381;
    wire N__26378;
    wire N__26373;
    wire N__26362;
    wire N__26361;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26340;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26328;
    wire N__26327;
    wire N__26326;
    wire N__26325;
    wire N__26324;
    wire N__26317;
    wire N__26310;
    wire N__26309;
    wire N__26308;
    wire N__26307;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26290;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26166;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26140;
    wire N__26135;
    wire N__26132;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26100;
    wire N__26097;
    wire N__26096;
    wire N__26093;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26077;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26047;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25962;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25951;
    wire N__25948;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25929;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25902;
    wire N__25899;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25882;
    wire N__25881;
    wire N__25878;
    wire N__25877;
    wire N__25876;
    wire N__25873;
    wire N__25866;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25851;
    wire N__25850;
    wire N__25843;
    wire N__25840;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25816;
    wire N__25813;
    wire N__25812;
    wire N__25811;
    wire N__25810;
    wire N__25809;
    wire N__25804;
    wire N__25801;
    wire N__25796;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25747;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25728;
    wire N__25727;
    wire N__25726;
    wire N__25725;
    wire N__25724;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25716;
    wire N__25709;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25683;
    wire N__25680;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25663;
    wire N__25660;
    wire N__25655;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25518;
    wire N__25515;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25447;
    wire N__25446;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25428;
    wire N__25425;
    wire N__25424;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25412;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25392;
    wire N__25391;
    wire N__25390;
    wire N__25387;
    wire N__25384;
    wire N__25383;
    wire N__25382;
    wire N__25381;
    wire N__25380;
    wire N__25379;
    wire N__25374;
    wire N__25369;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25348;
    wire N__25345;
    wire N__25336;
    wire N__25333;
    wire N__25332;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25291;
    wire N__25288;
    wire N__25287;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25270;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25218;
    wire N__25215;
    wire N__25214;
    wire N__25211;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25161;
    wire N__25158;
    wire N__25157;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25097;
    wire N__25094;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25066;
    wire N__25063;
    wire N__25058;
    wire N__25051;
    wire N__25050;
    wire N__25049;
    wire N__25046;
    wire N__25041;
    wire N__25036;
    wire N__25035;
    wire N__25034;
    wire N__25031;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24859;
    wire N__24856;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24842;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24786;
    wire N__24785;
    wire N__24784;
    wire N__24781;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24732;
    wire N__24731;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24678;
    wire N__24677;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24577;
    wire N__24576;
    wire N__24575;
    wire N__24572;
    wire N__24569;
    wire N__24568;
    wire N__24567;
    wire N__24566;
    wire N__24563;
    wire N__24562;
    wire N__24561;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24525;
    wire N__24524;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24480;
    wire N__24477;
    wire N__24476;
    wire N__24475;
    wire N__24474;
    wire N__24473;
    wire N__24470;
    wire N__24469;
    wire N__24468;
    wire N__24467;
    wire N__24466;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24455;
    wire N__24454;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24436;
    wire N__24435;
    wire N__24432;
    wire N__24431;
    wire N__24428;
    wire N__24423;
    wire N__24420;
    wire N__24419;
    wire N__24414;
    wire N__24407;
    wire N__24404;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24390;
    wire N__24387;
    wire N__24382;
    wire N__24379;
    wire N__24372;
    wire N__24369;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24328;
    wire N__24325;
    wire N__24322;
    wire N__24319;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24307;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24241;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24233;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24221;
    wire N__24218;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24180;
    wire N__24179;
    wire N__24176;
    wire N__24175;
    wire N__24174;
    wire N__24173;
    wire N__24172;
    wire N__24171;
    wire N__24170;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24152;
    wire N__24151;
    wire N__24150;
    wire N__24149;
    wire N__24144;
    wire N__24143;
    wire N__24142;
    wire N__24139;
    wire N__24132;
    wire N__24129;
    wire N__24124;
    wire N__24121;
    wire N__24116;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24096;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24076;
    wire N__24073;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23982;
    wire N__23977;
    wire N__23976;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23959;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23920;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23908;
    wire N__23905;
    wire N__23900;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23886;
    wire N__23885;
    wire N__23882;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23713;
    wire N__23712;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23695;
    wire N__23692;
    wire N__23689;
    wire N__23686;
    wire N__23683;
    wire N__23678;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23570;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23552;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23454;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23428;
    wire N__23427;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23349;
    wire N__23348;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23340;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23323;
    wire N__23320;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23293;
    wire N__23290;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23272;
    wire N__23271;
    wire N__23268;
    wire N__23263;
    wire N__23260;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23199;
    wire N__23198;
    wire N__23197;
    wire N__23196;
    wire N__23193;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23185;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23161;
    wire N__23154;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23132;
    wire N__23129;
    wire N__23124;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23010;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22985;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22860;
    wire N__22859;
    wire N__22856;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22836;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22719;
    wire N__22716;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22691;
    wire N__22688;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22655;
    wire N__22654;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22640;
    wire N__22637;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22515;
    wire N__22512;
    wire N__22509;
    wire N__22508;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22496;
    wire N__22493;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22252;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22237;
    wire N__22232;
    wire N__22225;
    wire N__22224;
    wire N__22221;
    wire N__22220;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22027;
    wire N__22026;
    wire N__22025;
    wire N__22024;
    wire N__22023;
    wire N__22022;
    wire N__22017;
    wire N__22012;
    wire N__22011;
    wire N__22010;
    wire N__22009;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21994;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21988;
    wire N__21987;
    wire N__21984;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21972;
    wire N__21969;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21948;
    wire N__21945;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21929;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21867;
    wire N__21866;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21858;
    wire N__21855;
    wire N__21854;
    wire N__21853;
    wire N__21852;
    wire N__21849;
    wire N__21848;
    wire N__21843;
    wire N__21840;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21826;
    wire N__21823;
    wire N__21822;
    wire N__21819;
    wire N__21814;
    wire N__21811;
    wire N__21810;
    wire N__21809;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21775;
    wire N__21768;
    wire N__21763;
    wire N__21760;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21744;
    wire N__21743;
    wire N__21740;
    wire N__21735;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21708;
    wire N__21705;
    wire N__21700;
    wire N__21695;
    wire N__21690;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21642;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21555;
    wire N__21552;
    wire N__21551;
    wire N__21548;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21523;
    wire N__21522;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21505;
    wire N__21504;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21493;
    wire N__21492;
    wire N__21489;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21471;
    wire N__21468;
    wire N__21467;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21445;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21387;
    wire N__21384;
    wire N__21383;
    wire N__21380;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21355;
    wire N__21350;
    wire N__21347;
    wire N__21346;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21330;
    wire N__21327;
    wire N__21322;
    wire N__21319;
    wire N__21314;
    wire N__21309;
    wire N__21306;
    wire N__21301;
    wire N__21298;
    wire N__21297;
    wire N__21294;
    wire N__21293;
    wire N__21290;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21275;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21253;
    wire N__21252;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21237;
    wire N__21232;
    wire N__21227;
    wire N__21224;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21198;
    wire N__21197;
    wire N__21196;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21182;
    wire N__21181;
    wire N__21178;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21126;
    wire N__21121;
    wire N__21116;
    wire N__21109;
    wire N__21106;
    wire N__21105;
    wire N__21104;
    wire N__21101;
    wire N__21096;
    wire N__21091;
    wire N__21090;
    wire N__21089;
    wire N__21086;
    wire N__21085;
    wire N__21082;
    wire N__21081;
    wire N__21078;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21053;
    wire N__21050;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21038;
    wire N__21033;
    wire N__21030;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21013;
    wire N__21006;
    wire N__21001;
    wire N__21000;
    wire N__20999;
    wire N__20998;
    wire N__20995;
    wire N__20992;
    wire N__20991;
    wire N__20988;
    wire N__20983;
    wire N__20982;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20964;
    wire N__20963;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20913;
    wire N__20912;
    wire N__20911;
    wire N__20908;
    wire N__20903;
    wire N__20900;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20801;
    wire N__20800;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20788;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20771;
    wire N__20770;
    wire N__20769;
    wire N__20764;
    wire N__20757;
    wire N__20752;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20613;
    wire N__20612;
    wire N__20609;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20590;
    wire N__20587;
    wire N__20578;
    wire N__20577;
    wire N__20576;
    wire N__20573;
    wire N__20568;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20556;
    wire N__20553;
    wire N__20550;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20529;
    wire N__20526;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20511;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20483;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20357;
    wire N__20356;
    wire N__20353;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20315;
    wire N__20312;
    wire N__20305;
    wire N__20304;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20242;
    wire N__20239;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20177;
    wire N__20176;
    wire N__20175;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20160;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20145;
    wire N__20142;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20107;
    wire N__20106;
    wire N__20101;
    wire N__20100;
    wire N__20099;
    wire N__20098;
    wire N__20097;
    wire N__20096;
    wire N__20095;
    wire N__20094;
    wire N__20093;
    wire N__20092;
    wire N__20091;
    wire N__20088;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20041;
    wire N__20040;
    wire N__20037;
    wire N__20032;
    wire N__20029;
    wire N__20028;
    wire N__20027;
    wire N__20026;
    wire N__20025;
    wire N__20024;
    wire N__20023;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20006;
    wire N__20001;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19834;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19813;
    wire N__19812;
    wire N__19809;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19752;
    wire N__19751;
    wire N__19750;
    wire N__19747;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19714;
    wire N__19711;
    wire N__19710;
    wire N__19709;
    wire N__19708;
    wire N__19707;
    wire N__19706;
    wire N__19705;
    wire N__19704;
    wire N__19703;
    wire N__19702;
    wire N__19701;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19693;
    wire N__19692;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19680;
    wire N__19677;
    wire N__19676;
    wire N__19675;
    wire N__19672;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19664;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19652;
    wire N__19649;
    wire N__19648;
    wire N__19645;
    wire N__19644;
    wire N__19643;
    wire N__19642;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19630;
    wire N__19625;
    wire N__19618;
    wire N__19617;
    wire N__19616;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19604;
    wire N__19601;
    wire N__19594;
    wire N__19587;
    wire N__19584;
    wire N__19579;
    wire N__19574;
    wire N__19567;
    wire N__19562;
    wire N__19559;
    wire N__19546;
    wire N__19541;
    wire N__19528;
    wire N__19527;
    wire N__19526;
    wire N__19525;
    wire N__19524;
    wire N__19523;
    wire N__19522;
    wire N__19521;
    wire N__19520;
    wire N__19519;
    wire N__19518;
    wire N__19517;
    wire N__19514;
    wire N__19513;
    wire N__19512;
    wire N__19509;
    wire N__19508;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19492;
    wire N__19489;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19475;
    wire N__19474;
    wire N__19473;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19463;
    wire N__19462;
    wire N__19459;
    wire N__19458;
    wire N__19457;
    wire N__19456;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19444;
    wire N__19439;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19423;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19403;
    wire N__19396;
    wire N__19387;
    wire N__19380;
    wire N__19375;
    wire N__19360;
    wire N__19357;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19257;
    wire N__19256;
    wire N__19255;
    wire N__19254;
    wire N__19253;
    wire N__19250;
    wire N__19249;
    wire N__19248;
    wire N__19247;
    wire N__19246;
    wire N__19243;
    wire N__19242;
    wire N__19241;
    wire N__19238;
    wire N__19237;
    wire N__19234;
    wire N__19233;
    wire N__19232;
    wire N__19231;
    wire N__19230;
    wire N__19229;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19221;
    wire N__19218;
    wire N__19217;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19203;
    wire N__19202;
    wire N__19201;
    wire N__19198;
    wire N__19193;
    wire N__19190;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19139;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19131;
    wire N__19130;
    wire N__19125;
    wire N__19122;
    wire N__19115;
    wire N__19112;
    wire N__19107;
    wire N__19104;
    wire N__19099;
    wire N__19094;
    wire N__19089;
    wire N__19082;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19053;
    wire N__19048;
    wire N__19035;
    wire N__19018;
    wire N__19015;
    wire N__19014;
    wire N__19013;
    wire N__19012;
    wire N__19011;
    wire N__19010;
    wire N__19009;
    wire N__19008;
    wire N__19007;
    wire N__19006;
    wire N__19005;
    wire N__19004;
    wire N__19001;
    wire N__19000;
    wire N__18997;
    wire N__18996;
    wire N__18995;
    wire N__18992;
    wire N__18991;
    wire N__18986;
    wire N__18979;
    wire N__18978;
    wire N__18977;
    wire N__18976;
    wire N__18973;
    wire N__18972;
    wire N__18969;
    wire N__18966;
    wire N__18965;
    wire N__18964;
    wire N__18961;
    wire N__18960;
    wire N__18957;
    wire N__18952;
    wire N__18945;
    wire N__18942;
    wire N__18937;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18914;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18872;
    wire N__18865;
    wire N__18858;
    wire N__18855;
    wire N__18844;
    wire N__18843;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18835;
    wire N__18834;
    wire N__18831;
    wire N__18830;
    wire N__18827;
    wire N__18822;
    wire N__18817;
    wire N__18814;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18735;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18580;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18572;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18549;
    wire N__18548;
    wire N__18545;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18535;
    wire N__18528;
    wire N__18527;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18513;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18396;
    wire N__18395;
    wire N__18394;
    wire N__18393;
    wire N__18392;
    wire N__18391;
    wire N__18390;
    wire N__18389;
    wire N__18386;
    wire N__18381;
    wire N__18378;
    wire N__18373;
    wire N__18372;
    wire N__18371;
    wire N__18370;
    wire N__18369;
    wire N__18368;
    wire N__18363;
    wire N__18362;
    wire N__18361;
    wire N__18360;
    wire N__18357;
    wire N__18356;
    wire N__18355;
    wire N__18354;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18340;
    wire N__18331;
    wire N__18330;
    wire N__18329;
    wire N__18328;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18316;
    wire N__18311;
    wire N__18306;
    wire N__18295;
    wire N__18288;
    wire N__18285;
    wire N__18268;
    wire N__18267;
    wire N__18266;
    wire N__18265;
    wire N__18264;
    wire N__18263;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18251;
    wire N__18248;
    wire N__18243;
    wire N__18232;
    wire N__18231;
    wire N__18230;
    wire N__18229;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18221;
    wire N__18220;
    wire N__18219;
    wire N__18218;
    wire N__18217;
    wire N__18214;
    wire N__18209;
    wire N__18204;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18145;
    wire N__18142;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18130;
    wire N__18129;
    wire N__18128;
    wire N__18127;
    wire N__18124;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18116;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18105;
    wire N__18104;
    wire N__18103;
    wire N__18102;
    wire N__18101;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18091;
    wire N__18090;
    wire N__18089;
    wire N__18088;
    wire N__18085;
    wire N__18084;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18060;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18043;
    wire N__18042;
    wire N__18039;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18031;
    wire N__18028;
    wire N__18027;
    wire N__18026;
    wire N__18019;
    wire N__18014;
    wire N__18009;
    wire N__18006;
    wire N__17997;
    wire N__17994;
    wire N__17989;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17973;
    wire N__17968;
    wire N__17963;
    wire N__17944;
    wire N__17943;
    wire N__17942;
    wire N__17941;
    wire N__17940;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17929;
    wire N__17922;
    wire N__17921;
    wire N__17920;
    wire N__17919;
    wire N__17918;
    wire N__17917;
    wire N__17916;
    wire N__17915;
    wire N__17912;
    wire N__17907;
    wire N__17904;
    wire N__17903;
    wire N__17902;
    wire N__17901;
    wire N__17898;
    wire N__17891;
    wire N__17888;
    wire N__17887;
    wire N__17884;
    wire N__17883;
    wire N__17880;
    wire N__17877;
    wire N__17870;
    wire N__17863;
    wire N__17856;
    wire N__17849;
    wire N__17836;
    wire N__17833;
    wire N__17830;
    wire N__17827;
    wire N__17824;
    wire N__17821;
    wire N__17818;
    wire N__17817;
    wire N__17814;
    wire N__17813;
    wire N__17812;
    wire N__17811;
    wire N__17808;
    wire N__17807;
    wire N__17806;
    wire N__17805;
    wire N__17804;
    wire N__17803;
    wire N__17802;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17790;
    wire N__17789;
    wire N__17786;
    wire N__17781;
    wire N__17778;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17758;
    wire N__17755;
    wire N__17748;
    wire N__17739;
    wire N__17734;
    wire N__17727;
    wire N__17722;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17679;
    wire N__17678;
    wire N__17677;
    wire N__17676;
    wire N__17675;
    wire N__17674;
    wire N__17673;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17659;
    wire N__17658;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17650;
    wire N__17649;
    wire N__17648;
    wire N__17647;
    wire N__17646;
    wire N__17641;
    wire N__17634;
    wire N__17629;
    wire N__17624;
    wire N__17621;
    wire N__17612;
    wire N__17599;
    wire N__17596;
    wire N__17595;
    wire N__17594;
    wire N__17593;
    wire N__17590;
    wire N__17589;
    wire N__17586;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17508;
    wire N__17505;
    wire N__17502;
    wire N__17499;
    wire N__17496;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17466;
    wire N__17465;
    wire N__17462;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17404;
    wire N__17403;
    wire N__17400;
    wire N__17397;
    wire N__17394;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17382;
    wire N__17379;
    wire N__17376;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17343;
    wire N__17342;
    wire N__17341;
    wire N__17340;
    wire N__17339;
    wire N__17338;
    wire N__17337;
    wire N__17336;
    wire N__17335;
    wire N__17332;
    wire N__17331;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17319;
    wire N__17314;
    wire N__17307;
    wire N__17306;
    wire N__17305;
    wire N__17304;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17280;
    wire N__17275;
    wire N__17270;
    wire N__17267;
    wire N__17260;
    wire N__17257;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17235;
    wire N__17234;
    wire N__17233;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17225;
    wire N__17224;
    wire N__17221;
    wire N__17220;
    wire N__17219;
    wire N__17218;
    wire N__17217;
    wire N__17212;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17204;
    wire N__17201;
    wire N__17200;
    wire N__17199;
    wire N__17196;
    wire N__17193;
    wire N__17190;
    wire N__17183;
    wire N__17180;
    wire N__17179;
    wire N__17178;
    wire N__17177;
    wire N__17176;
    wire N__17175;
    wire N__17174;
    wire N__17173;
    wire N__17172;
    wire N__17171;
    wire N__17170;
    wire N__17167;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17151;
    wire N__17140;
    wire N__17137;
    wire N__17132;
    wire N__17127;
    wire N__17116;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17028;
    wire N__17025;
    wire N__17022;
    wire N__17019;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16972;
    wire N__16971;
    wire N__16968;
    wire N__16965;
    wire N__16962;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16950;
    wire N__16947;
    wire N__16944;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16869;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16855;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16840;
    wire N__16837;
    wire N__16832;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16816;
    wire N__16815;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16804;
    wire N__16803;
    wire N__16800;
    wire N__16795;
    wire N__16792;
    wire N__16791;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16777;
    wire N__16774;
    wire N__16769;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16753;
    wire N__16752;
    wire N__16751;
    wire N__16748;
    wire N__16747;
    wire N__16744;
    wire N__16743;
    wire N__16740;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16728;
    wire N__16725;
    wire N__16722;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16706;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16689;
    wire N__16686;
    wire N__16683;
    wire N__16678;
    wire N__16675;
    wire N__16674;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16657;
    wire N__16654;
    wire N__16651;
    wire N__16646;
    wire N__16645;
    wire N__16644;
    wire N__16641;
    wire N__16636;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16602;
    wire N__16599;
    wire N__16594;
    wire N__16591;
    wire N__16588;
    wire N__16587;
    wire N__16586;
    wire N__16585;
    wire N__16584;
    wire N__16579;
    wire N__16578;
    wire N__16575;
    wire N__16572;
    wire N__16571;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16540;
    wire N__16539;
    wire N__16538;
    wire N__16535;
    wire N__16530;
    wire N__16525;
    wire N__16520;
    wire N__16515;
    wire N__16504;
    wire N__16503;
    wire N__16502;
    wire N__16501;
    wire N__16500;
    wire N__16499;
    wire N__16498;
    wire N__16495;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16470;
    wire N__16469;
    wire N__16468;
    wire N__16467;
    wire N__16464;
    wire N__16461;
    wire N__16456;
    wire N__16449;
    wire N__16446;
    wire N__16443;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16425;
    wire N__16420;
    wire N__16415;
    wire N__16402;
    wire N__16399;
    wire N__16396;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16311;
    wire N__16310;
    wire N__16309;
    wire N__16308;
    wire N__16303;
    wire N__16298;
    wire N__16295;
    wire N__16288;
    wire N__16285;
    wire N__16282;
    wire N__16281;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16179;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16168;
    wire N__16167;
    wire N__16166;
    wire N__16163;
    wire N__16158;
    wire N__16155;
    wire N__16150;
    wire N__16141;
    wire N__16140;
    wire N__16139;
    wire N__16138;
    wire N__16137;
    wire N__16136;
    wire N__16135;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16123;
    wire N__16118;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16099;
    wire N__16092;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16036;
    wire N__16033;
    wire N__16032;
    wire N__16031;
    wire N__16026;
    wire N__16023;
    wire N__16018;
    wire N__16017;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16000;
    wire N__15999;
    wire N__15998;
    wire N__15997;
    wire N__15996;
    wire N__15995;
    wire N__15994;
    wire N__15991;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15981;
    wire N__15976;
    wire N__15975;
    wire N__15972;
    wire N__15969;
    wire N__15966;
    wire N__15965;
    wire N__15964;
    wire N__15961;
    wire N__15960;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15942;
    wire N__15939;
    wire N__15938;
    wire N__15937;
    wire N__15936;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15921;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15903;
    wire N__15886;
    wire N__15885;
    wire N__15882;
    wire N__15879;
    wire N__15876;
    wire N__15875;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15863;
    wire N__15862;
    wire N__15861;
    wire N__15858;
    wire N__15853;
    wire N__15848;
    wire N__15841;
    wire N__15838;
    wire N__15835;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15817;
    wire N__15816;
    wire N__15811;
    wire N__15808;
    wire N__15807;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15793;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15685;
    wire N__15682;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15659;
    wire N__15656;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15648;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15630;
    wire N__15627;
    wire N__15622;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15517;
    wire N__15514;
    wire N__15513;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15505;
    wire N__15502;
    wire N__15499;
    wire N__15496;
    wire N__15493;
    wire N__15488;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15402;
    wire N__15399;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15379;
    wire N__15376;
    wire N__15373;
    wire N__15370;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15360;
    wire N__15357;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15343;
    wire N__15340;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15328;
    wire N__15325;
    wire N__15324;
    wire N__15323;
    wire N__15322;
    wire N__15319;
    wire N__15314;
    wire N__15311;
    wire N__15310;
    wire N__15309;
    wire N__15308;
    wire N__15305;
    wire N__15300;
    wire N__15297;
    wire N__15292;
    wire N__15291;
    wire N__15290;
    wire N__15285;
    wire N__15280;
    wire N__15275;
    wire N__15268;
    wire N__15265;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15238;
    wire N__15235;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15183;
    wire N__15182;
    wire N__15179;
    wire N__15174;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15159;
    wire N__15158;
    wire N__15155;
    wire N__15150;
    wire N__15145;
    wire N__15144;
    wire N__15143;
    wire N__15142;
    wire N__15141;
    wire N__15140;
    wire N__15139;
    wire N__15138;
    wire N__15121;
    wire N__15118;
    wire N__15115;
    wire N__15114;
    wire N__15113;
    wire N__15112;
    wire N__15111;
    wire N__15110;
    wire N__15109;
    wire N__15108;
    wire N__15107;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15081;
    wire N__15078;
    wire N__15077;
    wire N__15076;
    wire N__15073;
    wire N__15072;
    wire N__15067;
    wire N__15066;
    wire N__15065;
    wire N__15064;
    wire N__15061;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15040;
    wire N__15039;
    wire N__15036;
    wire N__15031;
    wire N__15022;
    wire N__15017;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14995;
    wire N__14994;
    wire N__14993;
    wire N__14992;
    wire N__14991;
    wire N__14988;
    wire N__14983;
    wire N__14978;
    wire N__14971;
    wire N__14968;
    wire N__14967;
    wire N__14966;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14954;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14940;
    wire N__14939;
    wire N__14938;
    wire N__14937;
    wire N__14934;
    wire N__14931;
    wire N__14928;
    wire N__14923;
    wire N__14920;
    wire N__14911;
    wire N__14910;
    wire N__14909;
    wire N__14904;
    wire N__14901;
    wire N__14898;
    wire N__14893;
    wire N__14892;
    wire N__14891;
    wire N__14890;
    wire N__14887;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14872;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14835;
    wire N__14834;
    wire N__14833;
    wire N__14830;
    wire N__14825;
    wire N__14822;
    wire N__14817;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14805;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14788;
    wire N__14787;
    wire N__14782;
    wire N__14779;
    wire N__14778;
    wire N__14775;
    wire N__14772;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14752;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14737;
    wire N__14736;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14719;
    wire N__14718;
    wire N__14717;
    wire N__14716;
    wire N__14715;
    wire N__14714;
    wire N__14711;
    wire N__14710;
    wire N__14707;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14695;
    wire N__14694;
    wire N__14693;
    wire N__14692;
    wire N__14691;
    wire N__14690;
    wire N__14689;
    wire N__14684;
    wire N__14679;
    wire N__14676;
    wire N__14673;
    wire N__14670;
    wire N__14665;
    wire N__14664;
    wire N__14659;
    wire N__14654;
    wire N__14651;
    wire N__14650;
    wire N__14645;
    wire N__14642;
    wire N__14637;
    wire N__14636;
    wire N__14633;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14604;
    wire N__14593;
    wire N__14590;
    wire N__14589;
    wire N__14586;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14574;
    wire N__14569;
    wire N__14566;
    wire N__14565;
    wire N__14564;
    wire N__14563;
    wire N__14558;
    wire N__14553;
    wire N__14548;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14536;
    wire N__14535;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14529;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14505;
    wire N__14504;
    wire N__14501;
    wire N__14498;
    wire N__14493;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14475;
    wire N__14472;
    wire N__14469;
    wire N__14464;
    wire N__14461;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire N__14436;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14415;
    wire N__14412;
    wire N__14409;
    wire N__14404;
    wire N__14401;
    wire N__14400;
    wire N__14397;
    wire N__14396;
    wire N__14393;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14381;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14367;
    wire N__14366;
    wire N__14363;
    wire N__14358;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14304;
    wire N__14303;
    wire N__14302;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14290;
    wire N__14287;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14259;
    wire N__14256;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14136;
    wire N__14133;
    wire N__14130;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14013;
    wire N__14012;
    wire N__14011;
    wire N__14010;
    wire N__14007;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13994;
    wire N__13993;
    wire N__13990;
    wire N__13985;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13914;
    wire N__13913;
    wire N__13910;
    wire N__13905;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13876;
    wire N__13873;
    wire N__13870;
    wire N__13867;
    wire N__13866;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13849;
    wire N__13848;
    wire N__13847;
    wire N__13846;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13834;
    wire N__13831;
    wire N__13826;
    wire N__13825;
    wire N__13822;
    wire N__13817;
    wire N__13814;
    wire N__13813;
    wire N__13806;
    wire N__13803;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13743;
    wire N__13740;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13681;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13657;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13645;
    wire N__13642;
    wire N__13639;
    wire N__13636;
    wire N__13633;
    wire N__13630;
    wire N__13627;
    wire N__13626;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13618;
    wire N__13615;
    wire N__13614;
    wire N__13613;
    wire N__13612;
    wire N__13609;
    wire N__13608;
    wire N__13605;
    wire N__13600;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13581;
    wire N__13570;
    wire N__13567;
    wire N__13564;
    wire N__13563;
    wire N__13560;
    wire N__13557;
    wire N__13552;
    wire N__13549;
    wire N__13546;
    wire N__13545;
    wire N__13542;
    wire N__13539;
    wire N__13534;
    wire N__13533;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13525;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13509;
    wire N__13508;
    wire N__13507;
    wire N__13506;
    wire N__13503;
    wire N__13496;
    wire N__13493;
    wire N__13486;
    wire N__13477;
    wire N__13476;
    wire N__13473;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13455;
    wire N__13452;
    wire N__13449;
    wire N__13444;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13436;
    wire N__13433;
    wire N__13432;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13404;
    wire N__13401;
    wire N__13398;
    wire N__13387;
    wire N__13384;
    wire N__13381;
    wire N__13380;
    wire N__13379;
    wire N__13378;
    wire N__13375;
    wire N__13370;
    wire N__13367;
    wire N__13360;
    wire N__13359;
    wire N__13356;
    wire N__13353;
    wire N__13348;
    wire N__13345;
    wire N__13342;
    wire N__13341;
    wire N__13338;
    wire N__13335;
    wire N__13330;
    wire N__13329;
    wire N__13328;
    wire N__13325;
    wire N__13320;
    wire N__13319;
    wire N__13318;
    wire N__13317;
    wire N__13316;
    wire N__13315;
    wire N__13314;
    wire N__13311;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13299;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13273;
    wire N__13270;
    wire N__13269;
    wire N__13266;
    wire N__13265;
    wire N__13264;
    wire N__13263;
    wire N__13260;
    wire N__13259;
    wire N__13256;
    wire N__13251;
    wire N__13248;
    wire N__13243;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13224;
    wire N__13223;
    wire N__13222;
    wire N__13219;
    wire N__13218;
    wire N__13217;
    wire N__13214;
    wire N__13213;
    wire N__13210;
    wire N__13209;
    wire N__13208;
    wire N__13207;
    wire N__13204;
    wire N__13201;
    wire N__13196;
    wire N__13195;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13181;
    wire N__13178;
    wire N__13177;
    wire N__13170;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13154;
    wire N__13151;
    wire N__13146;
    wire N__13135;
    wire N__13132;
    wire N__13131;
    wire N__13130;
    wire N__13129;
    wire N__13128;
    wire N__13127;
    wire N__13126;
    wire N__13123;
    wire N__13120;
    wire N__13119;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13111;
    wire N__13110;
    wire N__13107;
    wire N__13106;
    wire N__13105;
    wire N__13104;
    wire N__13101;
    wire N__13094;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13068;
    wire N__13067;
    wire N__13066;
    wire N__13063;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13042;
    wire N__13039;
    wire N__13036;
    wire N__13031;
    wire N__13028;
    wire N__13023;
    wire N__13012;
    wire N__13009;
    wire N__13006;
    wire N__13005;
    wire N__13004;
    wire N__13003;
    wire N__13002;
    wire N__13001;
    wire N__13000;
    wire N__12999;
    wire N__12998;
    wire N__12997;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12981;
    wire N__12978;
    wire N__12973;
    wire N__12972;
    wire N__12971;
    wire N__12970;
    wire N__12967;
    wire N__12962;
    wire N__12953;
    wire N__12952;
    wire N__12951;
    wire N__12950;
    wire N__12943;
    wire N__12936;
    wire N__12933;
    wire N__12928;
    wire N__12919;
    wire N__12916;
    wire N__12915;
    wire N__12914;
    wire N__12913;
    wire N__12912;
    wire N__12907;
    wire N__12904;
    wire N__12899;
    wire N__12898;
    wire N__12897;
    wire N__12890;
    wire N__12887;
    wire N__12886;
    wire N__12885;
    wire N__12884;
    wire N__12883;
    wire N__12882;
    wire N__12881;
    wire N__12880;
    wire N__12879;
    wire N__12878;
    wire N__12875;
    wire N__12870;
    wire N__12861;
    wire N__12856;
    wire N__12849;
    wire N__12838;
    wire N__12835;
    wire N__12834;
    wire N__12833;
    wire N__12832;
    wire N__12827;
    wire N__12826;
    wire N__12825;
    wire N__12824;
    wire N__12823;
    wire N__12818;
    wire N__12817;
    wire N__12814;
    wire N__12813;
    wire N__12810;
    wire N__12805;
    wire N__12802;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12794;
    wire N__12793;
    wire N__12792;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12774;
    wire N__12771;
    wire N__12766;
    wire N__12759;
    wire N__12742;
    wire N__12741;
    wire N__12736;
    wire N__12733;
    wire N__12730;
    wire N__12727;
    wire N__12726;
    wire N__12725;
    wire N__12722;
    wire N__12721;
    wire N__12720;
    wire N__12719;
    wire N__12718;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12696;
    wire N__12685;
    wire N__12682;
    wire N__12679;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12667;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12657;
    wire N__12656;
    wire N__12653;
    wire N__12648;
    wire N__12643;
    wire N__12640;
    wire N__12637;
    wire N__12634;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12604;
    wire N__12601;
    wire N__12598;
    wire N__12595;
    wire N__12592;
    wire N__12589;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12579;
    wire N__12576;
    wire N__12575;
    wire N__12574;
    wire N__12573;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12557;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12532;
    wire N__12529;
    wire N__12528;
    wire N__12525;
    wire N__12524;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12511;
    wire N__12502;
    wire N__12499;
    wire N__12496;
    wire N__12493;
    wire N__12490;
    wire N__12487;
    wire N__12484;
    wire N__12481;
    wire N__12478;
    wire N__12475;
    wire N__12472;
    wire N__12469;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12457;
    wire N__12454;
    wire N__12451;
    wire N__12448;
    wire N__12447;
    wire N__12446;
    wire N__12445;
    wire N__12444;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12420;
    wire N__12417;
    wire N__12414;
    wire N__12409;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12349;
    wire N__12346;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12338;
    wire N__12333;
    wire N__12330;
    wire N__12325;
    wire N__12324;
    wire N__12321;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12301;
    wire N__12296;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12241;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12136;
    wire N__12133;
    wire N__12130;
    wire N__12127;
    wire N__12124;
    wire N__12121;
    wire N__12118;
    wire N__12115;
    wire N__12114;
    wire N__12109;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12061;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12040;
    wire N__12037;
    wire N__12034;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12016;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__12001;
    wire N__11998;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11983;
    wire N__11982;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11953;
    wire N__11950;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11863;
    wire N__11860;
    wire N__11857;
    wire N__11854;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11767;
    wire N__11764;
    wire N__11761;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11689;
    wire N__11686;
    wire N__11683;
    wire N__11680;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire M_this_map_ram_read_data_4;
    wire M_this_ppu_sprites_addr_9;
    wire M_this_ppu_sprites_addr_8;
    wire M_this_ppu_sprites_addr_7;
    wire M_this_ppu_sprites_addr_6;
    wire VCCG0;
    wire GNDG0;
    wire port_nmib_0_i;
    wire port_clk_c;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire rgb_c_5;
    wire port_data_rw_0_i;
    wire rgb_c_0;
    wire rgb_c_1;
    wire rgb_c_3;
    wire rgb_c_4;
    wire \this_vga_ramdac.N_2870_reto ;
    wire rgb_c_2;
    wire \this_vga_ramdac.i2_mux_0 ;
    wire \this_vga_ramdac.N_2875_reto ;
    wire \this_vga_signals.un4_hsynclto7_0_cascade_ ;
    wire this_vga_signals_hsync_1_i;
    wire \this_vga_signals.un2_hsynclt7_cascade_ ;
    wire \this_vga_signals.hsync_1_0 ;
    wire this_vga_signals_hvisibility_i;
    wire \this_vga_signals.if_N_8_i_0_cascade_ ;
    wire \this_vga_signals.if_N_9_0_0_cascade_ ;
    wire \this_pixel_clk.M_counter_q_i_1 ;
    wire \this_pixel_clk.M_counter_qZ0Z_0 ;
    wire \this_vga_signals.mult1_un61_sum_0_3_cascade_ ;
    wire \this_vga_signals.N_614_1 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_0 ;
    wire \this_vga_signals.g0_i_x4_0_cascade_ ;
    wire \this_vga_signals.g0_i_x4_2 ;
    wire \this_vga_signals.N_931_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_esr_RNI0JBR6Z0Z_9 ;
    wire \this_vga_signals.un4_hsynclto3_0 ;
    wire \this_vga_signals.un2_hsynclt6_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_ ;
    wire \this_vga_signals.M_hcounter_d7lt7_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_d7lto7_1 ;
    wire this_vga_signals_vvisibility_i;
    wire \this_vga_signals.N_5_i_5 ;
    wire \this_vga_signals.mult1_un82_sum_c3_0 ;
    wire \this_vga_signals.g0_4_cascade_ ;
    wire \this_vga_signals.g0_7_0_cascade_ ;
    wire M_this_vga_signals_address_1;
    wire \this_vga_ramdac.N_24_mux ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1 ;
    wire \this_vga_signals.g1 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_3_0_0 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_3_0_0_cascade_ ;
    wire \this_vga_signals.g2_0_0 ;
    wire \this_vga_signals.if_N_9_0_0 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb1 ;
    wire \this_vga_signals.mult1_un61_sum_axb1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb2_1 ;
    wire \this_vga_signals.N_236_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_3_0 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_ ;
    wire \this_vga_signals.N_3_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1 ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_9 ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.SUM_3_i_0_0_3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ;
    wire \this_vga_signals.N_236 ;
    wire \this_vga_signals.SUM_3_i_0_0_3 ;
    wire \this_vga_signals.g0_1 ;
    wire \this_vga_signals.un6_vvisibilitylt8_cascade_ ;
    wire \this_vga_signals.vvisibility_1_cascade_ ;
    wire \this_vga_signals.vsync_1_3 ;
    wire \this_vga_signals.vsync_1_2_cascade_ ;
    wire this_vga_signals_vsync_1_i;
    wire \this_vga_signals.if_m7_0_x4_0_cascade_ ;
    wire \this_vga_signals.if_N_9_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_c2_0 ;
    wire \this_vga_signals.mult1_un82_sum_c3 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_c3 ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.d_N_12 ;
    wire \this_vga_signals.d_N_11 ;
    wire \this_vga_signals.M_hcounter_q_RNIUAKU9Z0Z_4 ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3 ;
    wire \this_vga_signals.N_2_7_0 ;
    wire \this_vga_signals.mult1_un75_sum_axb2 ;
    wire \this_vga_signals.mult1_un75_sum_axb1 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_3_d ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_hcounter_d7lt4 ;
    wire bfn_7_19_0_;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_7_20_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.N_614_0 ;
    wire \this_vga_signals.N_931_1 ;
    wire \this_vga_signals.vaddress_0_5_cascade_ ;
    wire \this_vga_signals.g0_31_N_4L6 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_4_cascade_ ;
    wire \this_vga_signals.g0_31_N_3L3 ;
    wire \this_vga_signals.g3_3_0 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_2_cascade_ ;
    wire \this_vga_signals.g0_8_0_cascade_ ;
    wire \this_vga_signals.vaddress_2_5_cascade_ ;
    wire \this_vga_signals.vaddress_3_0_6_cascade_ ;
    wire \this_vga_signals.g2_3_cascade_ ;
    wire \this_vga_signals.g1_1_1_cascade_ ;
    wire \this_vga_signals.g0_i_x4_0_2_cascade_ ;
    wire \this_vga_signals.vaddress_6_5 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_1_0_0 ;
    wire \this_vga_signals.vaddress_3_0_6 ;
    wire \this_vga_signals.vaddress_3_5_cascade_ ;
    wire \this_vga_signals.vaddress_3_6_cascade_ ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ;
    wire M_this_ppu_vram_data_3;
    wire \this_sprites_ram.mem_out_bus6_3 ;
    wire \this_sprites_ram.mem_out_bus2_3 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus4_3 ;
    wire \this_sprites_ram.mem_out_bus0_3 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus5_3 ;
    wire \this_sprites_ram.mem_out_bus1_3 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2 ;
    wire M_this_vga_signals_address_4;
    wire \this_sprites_ram.mem_out_bus7_0 ;
    wire \this_sprites_ram.mem_out_bus3_0 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3 ;
    wire M_this_vga_signals_address_2;
    wire \this_vga_ramdac.m19 ;
    wire \this_vga_ramdac.N_2874_reto ;
    wire \this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ;
    wire \this_sprites_ram.mem_out_bus7_3 ;
    wire \this_sprites_ram.mem_out_bus3_3 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ;
    wire bfn_10_11_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_10_12_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.vaddress_c2 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_cascade_ ;
    wire \this_vga_signals.g1_0_1 ;
    wire \this_vga_signals.g0_31_N_5L8 ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_0 ;
    wire \this_vga_signals.m9_1_cascade_ ;
    wire \this_vga_signals.g2_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_1_0 ;
    wire \this_vga_signals.g1_0_0_1_cascade_ ;
    wire \this_vga_signals.g2_0_1_cascade_ ;
    wire \this_vga_signals.vaddress_6_6 ;
    wire \this_vga_signals.N_4_1_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_ ;
    wire \this_vga_signals.g0_i_x4_0_0 ;
    wire \this_vga_signals.g1_4_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_1_0_0_1 ;
    wire \this_vga_signals.g0_2_0_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_0_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_3_2 ;
    wire M_this_vga_signals_address_3;
    wire \this_sprites_ram.mem_WE_6 ;
    wire \this_vga_signals.N_3_2_1 ;
    wire M_this_vga_signals_address_6;
    wire \this_vga_signals.M_vcounter_d7lto8_1 ;
    wire \this_vga_signals.M_lcounter_d_0_sqmuxa ;
    wire \this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_ ;
    wire N_2_0_cascade_;
    wire \this_vga_signals.M_pcounter_qZ0Z_0 ;
    wire M_counter_q_RNILQS8_1;
    wire \this_vga_signals.M_pcounter_q_3_1_cascade_ ;
    wire \this_vga_signals.M_pcounter_qZ0Z_1 ;
    wire N_3_0_cascade_;
    wire \this_vga_signals.M_pcounter_q_i_5_1 ;
    wire \this_vga_signals.M_pcounter_q_i_5_0 ;
    wire \this_vga_signals.M_hcounter_d7_0 ;
    wire \this_vga_signals.M_pcounter_q_3_0 ;
    wire \this_sprites_ram.mem_WE_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.N_1_4_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_axb1_0 ;
    wire \this_vga_signals.SUM_2_i_1_2_3_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ;
    wire \this_vga_signals.M_vcounter_q_8_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_q_7_repZ0Z1 ;
    wire \this_vga_signals.SUM_2_i_1_0_3 ;
    wire \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5Z0Z_0 ;
    wire \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJHZ0Z5 ;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i_cascade_;
    wire \this_vga_signals.N_50 ;
    wire \this_vga_signals.vaddress_1_6_cascade_ ;
    wire \this_vga_signals.if_m8_0_a3_1_1_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire \this_vga_signals.N_614_1_g ;
    wire \this_vga_signals.N_931_g ;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_1_cascade_ ;
    wire \this_vga_signals.if_N_5_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.vaddress_5_cascade_ ;
    wire \this_vga_signals.g1_0_0_0 ;
    wire \this_vga_signals.g0_1_2_0_1 ;
    wire \this_vga_signals.g0_1_2_cascade_ ;
    wire \this_vga_signals.g1_0_1_0_0 ;
    wire \this_vga_signals.g2_0 ;
    wire \this_vga_signals.g1_1_1 ;
    wire \this_vga_signals.N_5_i_0 ;
    wire \this_vga_signals.g0_2_0_2_x1 ;
    wire \this_vga_signals.g0_2_0_2_x0_cascade_ ;
    wire \this_vga_signals.g0_2_0_2_cascade_ ;
    wire \this_sprites_ram.mem_out_bus7_2 ;
    wire \this_sprites_ram.mem_out_bus3_2 ;
    wire \this_sprites_ram.mem_out_bus5_0 ;
    wire \this_sprites_ram.mem_out_bus1_0 ;
    wire \this_sprites_ram.mem_WE_8 ;
    wire \this_vga_ramdac.m6 ;
    wire \this_vga_ramdac.N_2871_reto ;
    wire G_384_cascade_;
    wire \this_vga_ramdac.N_2872_reto ;
    wire \this_vga_signals.M_lcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_lcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire G_384;
    wire \this_vga_ramdac.N_2873_reto ;
    wire N_3_0;
    wire N_2_0;
    wire M_this_vga_signals_pixel_clk_0_0;
    wire \this_sprites_ram.mem_WE_2 ;
    wire M_this_ppu_vram_addr_7;
    wire M_this_ppu_sprites_addr_4;
    wire \this_vga_signals.vaddress_4_5 ;
    wire \this_vga_signals.vaddress_5 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_0 ;
    wire \this_vga_signals.mult1_un47_sum_c3_cascade_ ;
    wire \this_vga_signals.N_5_i_0_0 ;
    wire \this_vga_signals.i2_mux ;
    wire \this_vga_signals.i2_mux_cascade_ ;
    wire \this_vga_signals.if_i2_mux_cascade_ ;
    wire \this_vga_signals.vaddress_0_6 ;
    wire \this_vga_signals.g2_2 ;
    wire m18x_N_3LZ0Z3;
    wire \this_vga_signals.M_vcounter_q_esr_RNI5BS7NZ0Z_5 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_0_0 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_0_x0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1_0_x1 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0 ;
    wire \this_vga_signals.g0_2_0_2 ;
    wire \this_vga_signals.g1_0_0_0_1 ;
    wire \this_vga_signals.N_51 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0 ;
    wire \this_vga_signals.g2_1 ;
    wire \this_vga_signals.g1_0 ;
    wire \this_vga_signals.g1_N_4L5_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5EZ0Z1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2 ;
    wire \this_vga_signals.g0_1_1 ;
    wire \this_vga_signals.d_N_3_0_i ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_x0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_cascade_ ;
    wire \this_vga_signals.g0_7 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_0 ;
    wire this_vga_signals_un5_vaddress_g1_1_0;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_0 ;
    wire \this_vga_signals.g1_2 ;
    wire \this_vga_signals.m21_0_1_1 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ;
    wire M_this_ppu_vram_data_0;
    wire \this_vga_ramdac.m16 ;
    wire M_this_vram_read_data_2;
    wire M_this_vram_read_data_1;
    wire M_this_vram_read_data_0;
    wire M_this_vram_read_data_3;
    wire \this_vga_ramdac.i2_mux ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.line_clk_1 ;
    wire M_this_vga_signals_line_clk_0_cascade_;
    wire \this_ppu.M_state_d_0_sqmuxa_cascade_ ;
    wire \this_sprites_ram.mem_out_bus5_2 ;
    wire \this_sprites_ram.mem_out_bus1_2 ;
    wire \this_sprites_ram.mem_out_bus7_1 ;
    wire \this_sprites_ram.mem_out_bus3_1 ;
    wire this_vga_signals_vvisibility;
    wire \this_vga_signals.vaddress_2_5 ;
    wire \this_vga_signals.g1_1_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_0_0 ;
    wire \this_vga_signals.g1_2_0_0 ;
    wire \this_vga_signals.if_i2_mux ;
    wire \this_vga_signals.M_vcounter_d7lt3 ;
    wire \this_vga_signals.M_vcounter_d7lt9_1 ;
    wire \this_vga_signals.M_vcounter_d7lt9_1_cascade_ ;
    wire \this_vga_signals.un4_lvisibility_1 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_0 ;
    wire \this_vga_signals.g0_0 ;
    wire \this_vga_signals.vaddress_1_5_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_0_1 ;
    wire \this_vga_signals.M_vcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.vaddress_1_5 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire \this_vga_signals.vaddress_2_6_cascade_ ;
    wire \this_vga_signals.g1_2_0 ;
    wire \this_vga_signals.M_vcounter_q_RNITP439_0Z0Z_2_cascade_ ;
    wire \this_vga_signals.m16_0_1 ;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0;
    wire \this_vga_signals.mult1_un54_sum_c3_1_cascade_ ;
    wire \this_vga_signals.g0_12 ;
    wire \this_vga_signals.M_vcounter_q_RNITP439Z0Z_2 ;
    wire \this_vga_signals.g2_1_1 ;
    wire \this_vga_signals.g1_1_1_0 ;
    wire \this_vga_signals.if_N_5_1 ;
    wire \this_vga_signals.g0_5_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2_0 ;
    wire \this_vga_signals.g0_1_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3 ;
    wire \this_vga_signals.g0_1_2_0_cascade_ ;
    wire \this_vga_signals.g1_3 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0_2_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1 ;
    wire if_generate_plus_mult1_un68_sum_axb1_520;
    wire \this_vga_signals.mult1_un61_sum_c3 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_i ;
    wire \this_vga_signals.g2_0_0_0 ;
    wire \this_vga_signals.g1_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i ;
    wire \this_vga_signals.g1_0_2 ;
    wire \this_vga_signals.g0_0_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_0_0_0 ;
    wire \this_vga_signals.m21_0_1 ;
    wire \this_vga_signals.i14_mux_i ;
    wire \this_vga_signals.N_25_0_0_cascade_ ;
    wire \this_vga_signals.i13_mux_0_i ;
    wire \this_vga_signals.if_i1_mux ;
    wire \this_vga_signals.g1_0_0_cascade_ ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_N_4L5_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_N_4L5_cascade_ ;
    wire \this_vga_signals.N_5_i ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire \this_ppu.un1_M_count_q_1_cry_0_0_c_RNOZ0 ;
    wire bfn_13_18_0_;
    wire \this_ppu.M_count_q_RNO_0Z0Z_1 ;
    wire \this_ppu.un1_M_count_q_1_cry_0 ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_2 ;
    wire \this_ppu.un1_M_count_q_1_cry_1 ;
    wire \this_ppu.un1_M_count_q_1_cry_2 ;
    wire \this_ppu.M_last_q_RNIMRAD5_4 ;
    wire \this_ppu.un1_M_count_q_1_cry_3 ;
    wire \this_ppu.un1_M_count_q_1_cry_4 ;
    wire \this_ppu.M_last_q_RNIMRAD5_5 ;
    wire \this_ppu.un1_M_count_q_1_cry_5 ;
    wire \this_ppu.un1_M_count_q_1_cry_6 ;
    wire \this_ppu.M_last_q_RNIMRAD5_1 ;
    wire \this_ppu.M_last_q_RNIMRAD5_0 ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_4 ;
    wire \this_ppu.un1_M_count_q_1_axb_0_cascade_ ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_6 ;
    wire \this_ppu.line_clk.M_last_qZ0 ;
    wire M_this_vga_signals_line_clk_0;
    wire \this_ppu.N_82_i_cascade_ ;
    wire \this_ppu.M_last_q_RNIMRAD5_3 ;
    wire \this_reset_cond.M_stage_qZ0Z_3 ;
    wire \this_sprites_ram.mem_out_bus4_0 ;
    wire \this_sprites_ram.mem_out_bus0_0 ;
    wire \this_sprites_ram.mem_out_bus6_0 ;
    wire \this_sprites_ram.mem_out_bus2_0 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z2 ;
    wire \this_vga_signals.if_N_5_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_4 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_5 ;
    wire \this_sprites_ram.mem_out_bus4_1 ;
    wire \this_sprites_ram.mem_out_bus0_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.mult1_un54_sum_c3_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0 ;
    wire \this_sprites_ram.mem_out_bus4_2 ;
    wire \this_sprites_ram.mem_out_bus0_2 ;
    wire \this_sprites_ram.mem_out_bus6_2 ;
    wire \this_sprites_ram.mem_out_bus2_2 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_ ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0 ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ;
    wire M_this_ppu_vram_data_1;
    wire \this_sprites_ram.mem_out_bus5_1 ;
    wire \this_sprites_ram.mem_out_bus1_1 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ;
    wire \this_ppu.N_91_cascade_ ;
    wire \this_ppu.M_count_qZ1Z_1 ;
    wire \this_ppu.M_count_qZ1Z_2 ;
    wire \this_ppu.M_count_qZ1Z_0 ;
    wire \this_ppu.M_state_q_i_1_cascade_ ;
    wire \this_ppu.M_last_q_RNIMRAD5_2 ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_3 ;
    wire \this_ppu.M_count_qZ1Z_3 ;
    wire \this_ppu.M_count_qZ1Z_4 ;
    wire \this_ppu.M_count_qZ0Z_6 ;
    wire \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4 ;
    wire \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_5 ;
    wire \this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4_cascade_ ;
    wire \this_ppu.M_state_d_0_sqmuxa_1 ;
    wire \this_ppu.M_state_d_0_sqmuxa_1_cascade_ ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_5 ;
    wire \this_ppu.M_count_qZ1Z_5 ;
    wire \this_ppu.M_state_q_i_1 ;
    wire \this_ppu.M_count_qZ0Z_7 ;
    wire \this_ppu.N_82_i ;
    wire \this_ppu.un1_M_count_q_1_axb_7 ;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire \this_sprites_ram.mem_out_bus6_1 ;
    wire \this_sprites_ram.mem_out_bus2_1 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2 ;
    wire M_this_ppu_vram_data_2;
    wire \this_ppu.M_state_qZ0Z_0 ;
    wire \this_ppu.M_state_qZ0Z_1 ;
    wire \this_sprites_ram.mem_WE_0 ;
    wire M_this_ppu_map_addr_6;
    wire M_this_ppu_map_addr_5;
    wire M_this_ppu_sprites_addr_5;
    wire \this_ppu.un1_M_vaddress_q_c2 ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire \this_sprites_ram.mem_WE_14 ;
    wire \this_sprites_ram.mem_WE_12 ;
    wire M_this_sprites_ram_write_en_0;
    wire \this_sprites_ram.mem_WE_10 ;
    wire M_this_sprites_ram_write_data_0;
    wire M_this_sprites_ram_write_data_1;
    wire \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux_cascade_ ;
    wire M_this_sprites_ram_write_data_2;
    wire \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ;
    wire M_this_sprites_ram_write_data_3;
    wire M_this_vga_ramdac_en_0;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire M_this_vga_signals_address_5;
    wire M_this_ppu_map_addr_7;
    wire \this_ppu.un1_M_vaddress_q_c5 ;
    wire \this_ppu.M_last_q_RNIQKTIG ;
    wire \this_ppu.M_vaddress_qZ0Z_7 ;
    wire M_this_ppu_map_addr_9;
    wire GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_8 ;
    wire \this_vga_signals.un23_i_a2_x1Z0Z_0_cascade_ ;
    wire dma_ac0Z0Z_5;
    wire this_vga_signals_un23_i_a2_1_3;
    wire this_vga_signals_un23_i_a2_4_2;
    wire this_vga_signals_un23_i_a2_3_2_cascade_;
    wire dma_c3_0;
    wire dma_axb0;
    wire M_this_state_q_RNI2S2SZ0Z_13;
    wire M_this_state_q_RNITS9I4Z0Z_7_cascade_;
    wire dma_ac0_5_i;
    wire dma_ac0_5_i_cascade_;
    wire dma_ac0_5_i_i;
    wire \this_vga_signals.un23_i_a2_4Z0Z_0 ;
    wire M_this_state_q_RNI6Q0SZ0Z_7;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8 ;
    wire \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_3 ;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10 ;
    wire M_this_ppu_vram_addr_0;
    wire M_this_ppu_vram_en_0;
    wire M_this_ppu_vram_addr_1;
    wire \this_ppu.M_state_d_0_sqmuxa ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_1 ;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_9 ;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2_cascade_ ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_2 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_3 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_10 ;
    wire M_this_state_q_RNIMJ231Z0Z_8;
    wire \this_vga_signals.M_this_state_q_ns_15 ;
    wire bfn_18_17_0_;
    wire un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0;
    wire un1_M_this_sprites_address_q_cry_0;
    wire M_this_sprites_address_qZ0Z_2;
    wire un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0;
    wire un1_M_this_sprites_address_q_cry_1;
    wire un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0;
    wire un1_M_this_sprites_address_q_cry_2;
    wire un1_M_this_sprites_address_q_cry_3;
    wire un1_M_this_sprites_address_q_cry_4;
    wire un1_M_this_sprites_address_q_cry_5;
    wire un1_M_this_sprites_address_q_cry_6;
    wire un1_M_this_sprites_address_q_cry_7;
    wire M_this_sprites_address_qZ0Z_8;
    wire un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0;
    wire bfn_18_18_0_;
    wire M_this_sprites_address_qZ0Z_9;
    wire un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0;
    wire un1_M_this_sprites_address_q_cry_8;
    wire M_this_sprites_address_qZ0Z_10;
    wire un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0;
    wire un1_M_this_sprites_address_q_cry_9;
    wire un1_M_this_sprites_address_q_cry_10;
    wire un1_M_this_sprites_address_q_cry_11;
    wire un1_M_this_sprites_address_q_cry_12;
    wire un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12 ;
    wire un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_13 ;
    wire un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0;
    wire M_this_sprites_address_qZ0Z_13;
    wire \this_vga_signals.M_this_state_q_ns_0_o2_0_0_0 ;
    wire \this_vga_signals.M_this_state_q_ns_0_o2_0_1Z0Z_0_cascade_ ;
    wire M_this_sprites_address_q_RNI1DGI7Z0Z_0;
    wire M_this_map_ram_read_data_5;
    wire \this_sprites_ram.mem_radregZ0Z_11 ;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_2_cascade_ ;
    wire \this_vga_signals.M_this_map_address_d_8_mZ0Z_2 ;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_9 ;
    wire \this_vga_signals.M_this_map_address_d_5_mZ0Z_9 ;
    wire M_this_ppu_map_addr_1;
    wire M_this_ppu_vram_addr_2;
    wire \this_ppu.un1_M_haddress_q_c2 ;
    wire M_this_ppu_map_addr_0;
    wire \this_ppu.M_vaddress_qZ0Z_6 ;
    wire this_ppu_M_vaddress_q_i_6;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_6 ;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6_cascade_ ;
    wire un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0;
    wire M_this_sprites_address_qZ0Z_6;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_0 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_5 ;
    wire un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0;
    wire \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_6 ;
    wire \this_vga_signals.N_294_cascade_ ;
    wire \this_vga_signals.un1_M_this_state_q_14Z0Z_1_cascade_ ;
    wire un1_M_this_state_q_14_0;
    wire this_vga_signals_un23_i_a2_1_1;
    wire un23_i_a2_1;
    wire \this_vga_signals.N_486 ;
    wire \this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_5 ;
    wire \this_vga_signals.N_486_cascade_ ;
    wire \this_vga_signals.N_438_1 ;
    wire this_vga_signals_M_this_state_q_ns_i_o2_0_12;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_11 ;
    wire \this_vga_signals.N_446_1 ;
    wire M_this_sprites_address_qZ0Z_11;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11 ;
    wire M_this_state_qZ0Z_1;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_ ;
    wire un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0;
    wire M_this_sprites_address_qZ0Z_7;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_7 ;
    wire un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_4 ;
    wire \this_vga_signals.un1_M_this_state_q_19_0 ;
    wire \this_vga_signals.M_this_state_d_1_sqmuxaZ0_cascade_ ;
    wire \this_vga_signals.N_399_0 ;
    wire \this_vga_signals.M_this_map_address_d_5_mZ0Z_5 ;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_5_cascade_ ;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_0 ;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_6 ;
    wire \this_vga_signals.M_this_map_address_d_5_mZ0Z_6_cascade_ ;
    wire M_this_map_address_q_RNICF7V6Z0Z_0;
    wire bfn_19_22_0_;
    wire un1_M_this_map_address_q_cry_0;
    wire M_this_map_address_qZ0Z_2;
    wire un1_M_this_map_address_q_cry_1_c_RNI8JSRZ0;
    wire un1_M_this_map_address_q_cry_1;
    wire un1_M_this_map_address_q_cry_2;
    wire un1_M_this_map_address_q_cry_3;
    wire M_this_map_address_qZ0Z_5;
    wire un1_M_this_map_address_q_cry_4_c_RNIESVRZ0;
    wire un1_M_this_map_address_q_cry_4;
    wire M_this_map_address_qZ0Z_6;
    wire un1_M_this_map_address_q_cry_5_c_RNIGV0SZ0;
    wire un1_M_this_map_address_q_cry_5;
    wire un1_M_this_map_address_q_cry_6_c_RNII22SZ0;
    wire un1_M_this_map_address_q_cry_6;
    wire un1_M_this_map_address_q_cry_7;
    wire bfn_19_23_0_;
    wire M_this_map_address_qZ0Z_9;
    wire un1_M_this_map_address_q_cry_8;
    wire un1_M_this_map_address_q_cry_8_c_RNIM84SZ0;
    wire \this_vga_signals.M_this_map_address_d_5_mZ0Z_7 ;
    wire M_this_map_address_qZ0Z_7;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_7 ;
    wire M_this_ppu_map_addr_2;
    wire \this_ppu.un1_M_haddress_q_c5 ;
    wire \this_ppu.M_last_q_RNI21NK5 ;
    wire \this_reset_cond.M_stage_qZ0Z_6 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire M_this_sprites_address_qZ0Z_5;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5 ;
    wire M_this_sprites_address_qZ0Z_1;
    wire N_389_0_cascade_;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1 ;
    wire M_this_state_q_fastZ0Z_15;
    wire N_297;
    wire \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_9 ;
    wire M_this_state_qZ0Z_9;
    wire \this_vga_signals.M_this_state_q_ns_0_a3_sxZ0Z_9_cascade_ ;
    wire port_address_in_4;
    wire port_rw_in;
    wire port_address_in_7;
    wire \this_vga_signals.N_291 ;
    wire \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1 ;
    wire port_address_in_5;
    wire port_address_in_6;
    wire \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_4_cascade_ ;
    wire \this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0 ;
    wire \this_vga_signals.N_444_1 ;
    wire this_vga_signals_M_this_state_q_ns_i_o2_0_14;
    wire M_this_state_q_fastZ0Z_14;
    wire M_this_sprites_address_qZ0Z_12;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_12 ;
    wire \this_vga_signals.M_this_external_address_d_5Z0Z_14 ;
    wire \this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_14 ;
    wire M_this_sprites_address_qZ0Z_4;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4 ;
    wire M_this_map_address_qZ0Z_0;
    wire \this_vga_signals.M_this_map_address_d_8_mZ0Z_0 ;
    wire M_this_sprites_address_qZ0Z_0;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0 ;
    wire \this_vga_signals.M_this_map_address_d_8_mZ0Z_1 ;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_1_cascade_ ;
    wire un1_M_this_map_address_q_cry_0_c_RNI6GRRZ0;
    wire M_this_map_address_qZ0Z_1;
    wire \this_vga_signals.M_this_map_address_d_8_mZ0Z_3_cascade_ ;
    wire un1_M_this_map_address_q_cry_2_c_RNIAMTRZ0;
    wire M_this_map_address_qZ0Z_3;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_3 ;
    wire \this_vga_signals.M_this_map_address_d_8_mZ0Z_4 ;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_4 ;
    wire un1_M_this_map_address_q_cry_3_c_RNICPURZ0;
    wire M_this_map_address_qZ0Z_4;
    wire M_this_state_qZ0Z_3;
    wire un1_M_this_state_q_12_0;
    wire \this_vga_signals.M_this_map_address_d_5_mZ0Z_8 ;
    wire \this_vga_signals.un1_M_this_map_ram_write_en_0 ;
    wire un1_M_this_map_address_q_cry_7_c_RNIK53SZ0;
    wire N_989_g;
    wire \this_vga_signals.N_469 ;
    wire M_this_state_qZ0Z_14;
    wire this_start_data_delay_M_last_q;
    wire port_enb_c;
    wire M_this_delay_clk_out_0;
    wire port_address_in_2;
    wire port_address_in_0;
    wire port_address_in_3;
    wire port_address_in_1;
    wire \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_10 ;
    wire \this_vga_signals.M_this_external_address_d_5Z0Z_13_cascade_ ;
    wire \this_vga_signals.M_this_state_d_1_sqmuxaZ0 ;
    wire \this_vga_signals.M_this_state_d_0_sqmuxaZ0Z_1 ;
    wire \this_vga_signals.un1_M_this_state_q_21_0_cascade_ ;
    wire \this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_13 ;
    wire M_this_state_qZ0Z_12;
    wire \this_vga_signals.N_293_1 ;
    wire M_this_state_qZ0Z_15;
    wire \this_vga_signals.M_this_map_ram_write_data_1_sqmuxa ;
    wire \this_vga_signals.N_293_cascade_ ;
    wire M_this_map_ram_read_data_7;
    wire \this_sprites_ram.mem_radregZ0Z_13 ;
    wire \this_vga_signals.M_this_external_address_d_8_mZ0Z_5 ;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_5 ;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_6 ;
    wire \this_vga_signals.M_this_external_address_d_8_mZ0Z_6_cascade_ ;
    wire M_this_map_address_qZ0Z_8;
    wire M_this_state_qZ0Z_4;
    wire \this_vga_signals.M_this_map_address_q_mZ0Z_8 ;
    wire M_this_reset_cond_out_0;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_7 ;
    wire \this_reset_cond.M_stage_qZ0Z_8 ;
    wire M_this_sprites_address_qZ0Z_3;
    wire M_this_state_qZ0Z_2;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3 ;
    wire M_this_state_d88_1_cascade_;
    wire \this_vga_signals.N_390_0 ;
    wire M_this_state_d88_12_cascade_;
    wire N_507_cascade_;
    wire N_508_cascade_;
    wire M_this_state_d88_11;
    wire M_this_state_d88_11_cascade_;
    wire M_this_state_d88_12;
    wire N_436;
    wire N_465;
    wire N_435;
    wire M_this_state_qsr_0_cascade_;
    wire N_466;
    wire led_c_1;
    wire M_this_state_d88;
    wire un1_M_this_state_q_16_0;
    wire bfn_22_20_0_;
    wire un1_M_this_external_address_q_cry_0;
    wire un1_M_this_external_address_q_cry_1;
    wire un1_M_this_external_address_q_cry_2;
    wire un1_M_this_external_address_q_cry_3;
    wire M_this_external_address_qZ0Z_5;
    wire un1_M_this_external_address_q_cry_4_c_RNIOSKBZ0;
    wire un1_M_this_external_address_q_cry_4;
    wire M_this_external_address_qZ0Z_6;
    wire un1_M_this_external_address_q_cry_5_c_RNIQVLBZ0;
    wire un1_M_this_external_address_q_cry_5;
    wire un1_M_this_external_address_q_cry_6;
    wire un1_M_this_external_address_q_cry_7;
    wire bfn_22_21_0_;
    wire un1_M_this_external_address_q_cry_8;
    wire un1_M_this_external_address_q_cry_9;
    wire un1_M_this_external_address_q_cry_10;
    wire un1_M_this_external_address_q_cry_11;
    wire M_this_external_address_qZ0Z_13;
    wire un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0;
    wire un1_M_this_external_address_q_cry_12;
    wire M_this_external_address_qZ0Z_14;
    wire un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0;
    wire un1_M_this_external_address_q_cry_13;
    wire un1_M_this_external_address_q_cry_14;
    wire un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_8_cascade_ ;
    wire M_this_external_address_qZ0Z_8;
    wire \this_vga_signals.M_this_external_address_d_5_mZ0Z_8 ;
    wire \this_vga_signals.M_this_external_address_d_8_mZ0Z_0_cascade_ ;
    wire M_this_external_address_q_RNIE44V9Z0Z_0;
    wire M_this_external_address_qZ0Z_0;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_0 ;
    wire \this_vga_signals.M_this_external_address_d_5_mZ0Z_9 ;
    wire un1_M_this_external_address_q_cry_8_c_RNI09PBZ0;
    wire \this_vga_signals.M_this_external_address_d_5_mZ0Z_11_cascade_ ;
    wire un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0;
    wire M_this_external_address_qZ0Z_11;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_11 ;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_3_cascade_ ;
    wire un1_M_this_external_address_q_cry_2_c_RNIKMIBZ0;
    wire M_this_external_address_qZ0Z_3;
    wire \this_vga_signals.M_this_external_address_d_8_mZ0Z_3 ;
    wire M_this_data_count_q_s_0;
    wire M_this_state_qZ0Z_10;
    wire \this_vga_signals.N_292_cascade_ ;
    wire \this_vga_signals.M_this_external_address_d_2_sqmuxaZ0 ;
    wire M_this_state_d88_9;
    wire N_506;
    wire N_509;
    wire N_510_cascade_;
    wire N_511;
    wire N_512;
    wire M_this_data_count_qZ0Z_0;
    wire bfn_23_17_0_;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_data_count_q_s_1;
    wire M_this_data_count_q_cry_0;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_q_s_2;
    wire M_this_data_count_q_cry_1;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_q_s_3;
    wire M_this_data_count_q_cry_2;
    wire M_this_data_count_qZ0Z_4;
    wire M_this_data_count_q_s_4;
    wire M_this_data_count_q_cry_3;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_q_s_5;
    wire M_this_data_count_q_cry_4;
    wire M_this_data_count_qZ0Z_6;
    wire M_this_data_count_q_s_6;
    wire M_this_data_count_q_cry_5;
    wire M_this_data_count_q_cry_6;
    wire M_this_data_count_q_cry_7;
    wire bfn_23_18_0_;
    wire M_this_data_count_q_cry_8;
    wire M_this_data_count_q_cry_9;
    wire M_this_data_count_q_cry_10;
    wire M_this_data_count_q_cry_11;
    wire M_this_data_count_q_cry_12;
    wire CONSTANT_ONE_NET;
    wire M_this_data_count_q_cry_13;
    wire M_this_data_count_q_cry_14;
    wire M_this_map_ram_read_data_6;
    wire \this_sprites_ram.mem_radregZ0Z_12 ;
    wire M_this_state_qZ0Z_7;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_1 ;
    wire \this_vga_signals.M_this_external_address_d_8_mZ0Z_1_cascade_ ;
    wire un1_M_this_external_address_q_cry_0_c_RNIGGGBZ0;
    wire M_this_external_address_qZ0Z_1;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_2 ;
    wire \this_vga_signals.M_this_external_address_d_8_mZ0Z_2_cascade_ ;
    wire un1_M_this_external_address_q_cry_1_c_RNIIJHBZ0;
    wire M_this_external_address_qZ0Z_2;
    wire \this_vga_signals.M_this_external_address_d_8_mZ0Z_4 ;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_4 ;
    wire un1_M_this_external_address_q_cry_3_c_RNIMPJBZ0;
    wire M_this_external_address_qZ0Z_4;
    wire \this_vga_signals.M_this_external_address_d_5_i_mZ0Z_15_cascade_ ;
    wire un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0;
    wire M_this_external_address_qZ0Z_15;
    wire \this_vga_signals.M_this_external_address_q_i_mZ0Z_15 ;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_7 ;
    wire \this_vga_signals.M_this_external_address_d_8_mZ0Z_7_cascade_ ;
    wire un1_M_this_external_address_q_cry_6_c_RNIS2NBZ0;
    wire M_this_external_address_qZ0Z_7;
    wire \this_vga_signals.M_this_external_address_d_5_mZ0Z_10_cascade_ ;
    wire un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0;
    wire M_this_external_address_qZ0Z_10;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_10 ;
    wire M_this_external_address_qZ0Z_9;
    wire M_this_state_qZ0Z_6;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_9 ;
    wire M_this_state_qZ0Z_5;
    wire \this_vga_signals.M_this_external_address_d_5_mZ0Z_12 ;
    wire \this_vga_signals.un1_M_this_state_q_21_0 ;
    wire \this_vga_signals.M_this_external_address_q_mZ0Z_12 ;
    wire un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0;
    wire M_this_external_address_qZ0Z_12;
    wire M_this_map_ram_write_data_3;
    wire M_this_state_qZ0Z_13;
    wire N_391_0;
    wire \this_vga_signals.un1_M_this_state_q_18Z0Z_1 ;
    wire M_this_state_qZ0Z_11;
    wire \this_vga_signals.N_387_0 ;
    wire \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0 ;
    wire N_513;
    wire M_this_data_count_q_s_7;
    wire M_this_data_count_qZ0Z_7;
    wire M_this_data_count_q_s_8;
    wire N_514_cascade_;
    wire M_this_data_count_q_s_9;
    wire N_515_cascade_;
    wire M_this_data_count_q_s_11;
    wire M_this_data_count_q_s_12;
    wire N_518_cascade_;
    wire M_this_data_count_qZ0Z_12;
    wire M_this_data_count_q_s_14;
    wire N_520_cascade_;
    wire M_this_data_count_qZ0Z_14;
    wire M_this_data_count_q_s_15;
    wire N_521_cascade_;
    wire M_this_data_count_qZ0Z_15;
    wire N_517;
    wire \this_vga_signals.M_this_data_count_q_3_bmZ0Z_10 ;
    wire M_this_data_count_q_cry_9_THRU_CO;
    wire M_this_data_count_q_3_10_cascade_;
    wire M_this_state_qZ0Z_8;
    wire N_389_0;
    wire M_this_reset_cond_out_g_0;
    wire \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8_cascade_ ;
    wire \this_vga_signals.M_this_data_count_q_3_bmZ0Z_13 ;
    wire \this_vga_signals.M_this_data_count_q_3_amZ0Z_13_cascade_ ;
    wire M_this_data_count_q_3_sn_N_2;
    wire M_this_data_count_q_cry_12_THRU_CO;
    wire M_this_data_count_q_3_13_cascade_;
    wire N_570_0_i;
    wire M_this_data_count_qZ0Z_13;
    wire clk_0_c_g;
    wire M_this_data_count_qe_0_i;
    wire M_this_data_count_qZ0Z_9;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_qZ0Z_8;
    wire M_this_state_d88_10;
    wire M_this_data_count_qZ0Z_10;
    wire \this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8 ;
    wire \this_vga_signals.M_this_data_count_q_3_amZ0Z_10 ;
    wire M_this_map_ram_write_data_6;
    wire M_this_map_ram_write_data_7;
    wire \this_ppu.M_haddress_qZ0Z_7 ;
    wire M_this_ppu_map_addr_4;
    wire M_this_ppu_vram_addr_6;
    wire M_this_ppu_vram_addr_i_6;
    wire M_this_map_ram_write_data_2;
    wire M_this_map_ram_write_data_1;
    wire M_this_map_ram_write_data_0;
    wire M_this_map_ram_write_data_5;
    wire M_this_map_ram_write_en_0;
    wire M_this_map_ram_write_data_4;
    wire port_data_c_3;
    wire port_data_c_2;
    wire \this_vga_signals.M_this_external_address_d21Z0Z_2_cascade_ ;
    wire \this_vga_signals.M_this_external_address_dZ0Z21 ;
    wire port_data_c_1;
    wire \this_vga_signals.M_this_external_address_d21Z0Z_2 ;
    wire port_data_c_0;
    wire \this_vga_signals.M_this_external_address_dZ0Z22 ;
    wire port_data_c_5;
    wire port_data_c_6;
    wire port_data_c_7;
    wire port_data_c_4;
    wire \this_vga_signals.M_this_external_address_d21Z0Z_6 ;
    wire _gnd_net_;

    defparam \this_map_ram.mem_mem_0_0_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_0_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,M_this_ppu_sprites_addr_9,dangling_wire_2,dangling_wire_3,dangling_wire_4,M_this_ppu_sprites_addr_8,dangling_wire_5,dangling_wire_6,dangling_wire_7,M_this_ppu_sprites_addr_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,M_this_ppu_sprites_addr_6,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__21433,N__23860,N__21574,N__20539,N__20506,N__33160,N__33094,N__25120,N__23595,N__23959}),
            .WADDR({dangling_wire_13,N__25234,N__27676,N__25171,N__24697,N__24748,N__26518,N__26593,N__24808,N__26647,N__26119}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__30400,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__33073,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__33067,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__33058,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__32057),
            .RE(N__30145),
            .WCLKE(N__33044),
            .WCLK(N__32058),
            .WE(N__30156));
    defparam \this_map_ram.mem_mem_0_1_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_1_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_42,dangling_wire_43,M_this_map_ram_read_data_7,dangling_wire_44,dangling_wire_45,dangling_wire_46,M_this_map_ram_read_data_6,dangling_wire_47,dangling_wire_48,dangling_wire_49,M_this_map_ram_read_data_5,dangling_wire_50,dangling_wire_51,dangling_wire_52,M_this_map_ram_read_data_4,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__21427,N__23854,N__21568,N__20533,N__20500,N__33154,N__33088,N__25113,N__23583,N__23949}),
            .WADDR({dangling_wire_55,N__25228,N__27670,N__25165,N__24691,N__24742,N__26512,N__26587,N__24802,N__26641,N__26113}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__33187,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__31471,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__33052,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__32947,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__32061),
            .RE(N__30160),
            .WCLKE(N__33045),
            .WCLK(N__32062),
            .WE(N__30155));
    defparam \this_sprites_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,\this_sprites_ram.mem_out_bus0_1 ,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,\this_sprites_ram.mem_out_bus0_0 ,dangling_wire_95,dangling_wire_96,dangling_wire_97}),
            .RADDR({N__11326,N__11773,N__11665,N__11551,N__11437,N__20455,N__15613,N__15763,N__23545,N__22177,N__22372}),
            .WADDR({N__22819,N__22966,N__23113,N__24340,N__23812,N__24973,N__26263,N__28366,N__22618,N__25618,N__26062}),
            .MASK({dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113}),
            .WDATA({dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,N__21297,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,N__21388,dangling_wire_125,dangling_wire_126,dangling_wire_127}),
            .RCLKE(),
            .RCLK(N__31937),
            .RE(N__30039),
            .WCLKE(N__20866),
            .WCLK(N__31938),
            .WE(N__30041));
    defparam \this_sprites_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,\this_sprites_ram.mem_out_bus0_3 ,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,\this_sprites_ram.mem_out_bus0_2 ,dangling_wire_139,dangling_wire_140,dangling_wire_141}),
            .RADDR({N__11320,N__11767,N__11659,N__11545,N__11431,N__20449,N__15607,N__15757,N__23539,N__22171,N__22366}),
            .WADDR({N__22813,N__22960,N__23107,N__24334,N__23806,N__24967,N__26257,N__28360,N__22612,N__25612,N__26056}),
            .MASK({dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157}),
            .WDATA({dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,N__21089,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,N__21195,dangling_wire_169,dangling_wire_170,dangling_wire_171}),
            .RCLKE(),
            .RCLK(N__31939),
            .RE(N__30038),
            .WCLKE(N__20862),
            .WCLK(N__31940),
            .WE(N__30040));
    defparam \this_sprites_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,\this_sprites_ram.mem_out_bus1_1 ,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,\this_sprites_ram.mem_out_bus1_0 ,dangling_wire_183,dangling_wire_184,dangling_wire_185}),
            .RADDR({N__11314,N__11761,N__11653,N__11539,N__11425,N__20443,N__15601,N__15751,N__23533,N__22165,N__22360}),
            .WADDR({N__22807,N__22954,N__23101,N__24328,N__23800,N__24961,N__26251,N__28354,N__22606,N__25606,N__26050}),
            .MASK({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .WDATA({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,N__21289,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,N__21383,dangling_wire_213,dangling_wire_214,dangling_wire_215}),
            .RCLKE(),
            .RCLK(N__31942),
            .RE(N__29948),
            .WCLKE(N__20836),
            .WCLK(N__31943),
            .WE(N__30042));
    defparam \this_sprites_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,\this_sprites_ram.mem_out_bus1_3 ,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,\this_sprites_ram.mem_out_bus1_2 ,dangling_wire_227,dangling_wire_228,dangling_wire_229}),
            .RADDR({N__11308,N__11755,N__11647,N__11533,N__11419,N__20437,N__15595,N__15745,N__23527,N__22159,N__22354}),
            .WADDR({N__22801,N__22948,N__23095,N__24322,N__23794,N__24955,N__26245,N__28348,N__22600,N__25600,N__26044}),
            .MASK({dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245}),
            .WDATA({dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,N__21077,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,N__21182,dangling_wire_257,dangling_wire_258,dangling_wire_259}),
            .RCLKE(),
            .RCLK(N__31947),
            .RE(N__29947),
            .WCLKE(N__20832),
            .WCLK(N__31948),
            .WE(N__29961));
    defparam \this_sprites_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,\this_sprites_ram.mem_out_bus2_1 ,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,\this_sprites_ram.mem_out_bus2_0 ,dangling_wire_271,dangling_wire_272,dangling_wire_273}),
            .RADDR({N__11302,N__11749,N__11641,N__11527,N__11413,N__20431,N__15589,N__15739,N__23521,N__22153,N__22348}),
            .WADDR({N__22795,N__22942,N__23089,N__24316,N__23788,N__24949,N__26239,N__28342,N__22594,N__25594,N__26038}),
            .MASK({dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289}),
            .WDATA({dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,N__21275,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,N__21372,dangling_wire_301,dangling_wire_302,dangling_wire_303}),
            .RCLKE(),
            .RCLK(N__31960),
            .RE(N__29848),
            .WCLKE(N__20752),
            .WCLK(N__31959),
            .WE(N__29962));
    defparam \this_sprites_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,\this_sprites_ram.mem_out_bus2_3 ,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,\this_sprites_ram.mem_out_bus2_2 ,dangling_wire_315,dangling_wire_316,dangling_wire_317}),
            .RADDR({N__11296,N__11743,N__11635,N__11521,N__11407,N__20425,N__15583,N__15733,N__23515,N__22147,N__22342}),
            .WADDR({N__22789,N__22936,N__23083,N__24310,N__23782,N__24943,N__26233,N__28336,N__22588,N__25588,N__26032}),
            .MASK({dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333}),
            .WDATA({dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,N__21090,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,N__21196,dangling_wire_345,dangling_wire_346,dangling_wire_347}),
            .RCLKE(),
            .RCLK(N__31970),
            .RE(N__29836),
            .WCLKE(N__20751),
            .WCLK(N__31971),
            .WE(N__29766));
    defparam \this_sprites_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,\this_sprites_ram.mem_out_bus3_1 ,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,\this_sprites_ram.mem_out_bus3_0 ,dangling_wire_359,dangling_wire_360,dangling_wire_361}),
            .RADDR({N__11290,N__11737,N__11629,N__11515,N__11401,N__20419,N__15577,N__15727,N__23509,N__22141,N__22336}),
            .WADDR({N__22783,N__22930,N__23077,N__24304,N__23776,N__24937,N__26227,N__28330,N__22582,N__25582,N__26026}),
            .MASK({dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377}),
            .WDATA({dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,N__21252,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,N__21355,dangling_wire_389,dangling_wire_390,dangling_wire_391}),
            .RCLKE(),
            .RCLK(N__31985),
            .RE(N__29869),
            .WCLKE(N__15403),
            .WCLK(N__31986),
            .WE(N__29935));
    defparam \this_sprites_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,\this_sprites_ram.mem_out_bus3_3 ,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,\this_sprites_ram.mem_out_bus3_2 ,dangling_wire_403,dangling_wire_404,dangling_wire_405}),
            .RADDR({N__11284,N__11731,N__11623,N__11509,N__11395,N__20413,N__15571,N__15721,N__23503,N__22135,N__22330}),
            .WADDR({N__22777,N__22924,N__23071,N__24298,N__23770,N__24931,N__26221,N__28324,N__22576,N__25576,N__26020}),
            .MASK({dangling_wire_406,dangling_wire_407,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421}),
            .WDATA({dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,N__21081,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,N__21177,dangling_wire_433,dangling_wire_434,dangling_wire_435}),
            .RCLKE(),
            .RCLK(N__31999),
            .RE(N__29876),
            .WCLKE(N__15402),
            .WCLK(N__32000),
            .WE(N__30030));
    defparam \this_sprites_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,\this_sprites_ram.mem_out_bus4_1 ,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,\this_sprites_ram.mem_out_bus4_0 ,dangling_wire_447,dangling_wire_448,dangling_wire_449}),
            .RADDR({N__11278,N__11725,N__11617,N__11503,N__11389,N__20407,N__15565,N__15715,N__23497,N__22129,N__22324}),
            .WADDR({N__22771,N__22918,N__23065,N__24292,N__23764,N__24925,N__26215,N__28318,N__22570,N__25570,N__26014}),
            .MASK({dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465}),
            .WDATA({dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,N__21237,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,N__21346,dangling_wire_477,dangling_wire_478,dangling_wire_479}),
            .RCLKE(),
            .RCLK(N__32013),
            .RE(N__29966),
            .WCLKE(N__14334),
            .WCLK(N__32014),
            .WE(N__30031));
    defparam \this_sprites_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,\this_sprites_ram.mem_out_bus4_3 ,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,\this_sprites_ram.mem_out_bus4_2 ,dangling_wire_491,dangling_wire_492,dangling_wire_493}),
            .RADDR({N__11272,N__11719,N__11611,N__11497,N__11383,N__20401,N__15559,N__15709,N__23491,N__22123,N__22318}),
            .WADDR({N__22765,N__22912,N__23059,N__24286,N__23758,N__24919,N__26209,N__28312,N__22564,N__25564,N__26008}),
            .MASK({dangling_wire_494,dangling_wire_495,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509}),
            .WDATA({dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,N__21049,dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,N__21181,dangling_wire_521,dangling_wire_522,dangling_wire_523}),
            .RCLKE(),
            .RCLK(N__32030),
            .RE(N__29967),
            .WCLKE(N__14338),
            .WCLK(N__32031),
            .WE(N__30085));
    defparam \this_sprites_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_524,dangling_wire_525,dangling_wire_526,dangling_wire_527,\this_sprites_ram.mem_out_bus5_1 ,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,dangling_wire_533,dangling_wire_534,\this_sprites_ram.mem_out_bus5_0 ,dangling_wire_535,dangling_wire_536,dangling_wire_537}),
            .RADDR({N__11266,N__11713,N__11605,N__11491,N__11377,N__20395,N__15553,N__15703,N__23485,N__22117,N__22312}),
            .WADDR({N__22759,N__22906,N__23053,N__24280,N__23752,N__24913,N__26203,N__28306,N__22558,N__25558,N__26002}),
            .MASK({dangling_wire_538,dangling_wire_539,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553}),
            .WDATA({dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,N__21282,dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,N__21365,dangling_wire_565,dangling_wire_566,dangling_wire_567}),
            .RCLKE(),
            .RCLK(N__32042),
            .RE(N__30043),
            .WCLKE(N__14445),
            .WCLK(N__32043),
            .WE(N__30054));
    defparam \this_sprites_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_568,dangling_wire_569,dangling_wire_570,dangling_wire_571,\this_sprites_ram.mem_out_bus5_3 ,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,dangling_wire_577,dangling_wire_578,\this_sprites_ram.mem_out_bus5_2 ,dangling_wire_579,dangling_wire_580,dangling_wire_581}),
            .RADDR({N__11260,N__11707,N__11599,N__11485,N__11371,N__20389,N__15547,N__15697,N__23479,N__22111,N__22306}),
            .WADDR({N__22753,N__22900,N__23047,N__24274,N__23746,N__24907,N__26197,N__28300,N__22552,N__25552,N__25996}),
            .MASK({dangling_wire_582,dangling_wire_583,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597}),
            .WDATA({dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,N__21070,dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,N__21197,dangling_wire_609,dangling_wire_610,dangling_wire_611}),
            .RCLKE(),
            .RCLK(N__32049),
            .RE(N__30044),
            .WCLKE(N__14446),
            .WCLK(N__32050),
            .WE(N__30089));
    defparam \this_sprites_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_612,dangling_wire_613,dangling_wire_614,dangling_wire_615,\this_sprites_ram.mem_out_bus6_1 ,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,dangling_wire_621,dangling_wire_622,\this_sprites_ram.mem_out_bus6_0 ,dangling_wire_623,dangling_wire_624,dangling_wire_625}),
            .RADDR({N__11254,N__11701,N__11593,N__11479,N__11365,N__20383,N__15541,N__15691,N__23473,N__22105,N__22300}),
            .WADDR({N__22747,N__22894,N__23041,N__24268,N__23740,N__24901,N__26191,N__28294,N__22546,N__25546,N__25990}),
            .MASK({dangling_wire_626,dangling_wire_627,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641}),
            .WDATA({dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,N__21293,dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,N__21379,dangling_wire_653,dangling_wire_654,dangling_wire_655}),
            .RCLKE(),
            .RCLK(N__32051),
            .RE(N__30090),
            .WCLKE(N__15792),
            .WCLK(N__32052),
            .WE(N__30092));
    defparam \this_sprites_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_656,dangling_wire_657,dangling_wire_658,dangling_wire_659,\this_sprites_ram.mem_out_bus6_3 ,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,dangling_wire_665,dangling_wire_666,\this_sprites_ram.mem_out_bus6_2 ,dangling_wire_667,dangling_wire_668,dangling_wire_669}),
            .RADDR({N__11248,N__11695,N__11587,N__11473,N__11359,N__20377,N__15535,N__15685,N__23467,N__22099,N__22294}),
            .WADDR({N__22741,N__22888,N__23035,N__24262,N__23734,N__24895,N__26185,N__28288,N__22540,N__25540,N__25984}),
            .MASK({dangling_wire_670,dangling_wire_671,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685}),
            .WDATA({dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,N__21085,dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,N__21198,dangling_wire_697,dangling_wire_698,dangling_wire_699}),
            .RCLKE(),
            .RCLK(N__32053),
            .RE(N__30091),
            .WCLKE(N__15793),
            .WCLK(N__32054),
            .WE(N__30093));
    defparam \this_sprites_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_700,dangling_wire_701,dangling_wire_702,dangling_wire_703,\this_sprites_ram.mem_out_bus7_1 ,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,dangling_wire_709,dangling_wire_710,\this_sprites_ram.mem_out_bus7_0 ,dangling_wire_711,dangling_wire_712,dangling_wire_713}),
            .RADDR({N__11242,N__11689,N__11581,N__11467,N__11353,N__20371,N__15529,N__15678,N__23461,N__22093,N__22288}),
            .WADDR({N__22735,N__22882,N__23029,N__24256,N__23728,N__24889,N__26179,N__28282,N__22534,N__25534,N__25978}),
            .MASK({dangling_wire_714,dangling_wire_715,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,dangling_wire_723,dangling_wire_724,dangling_wire_725,dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729}),
            .WDATA({dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,N__21298,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,N__21387,dangling_wire_741,dangling_wire_742,dangling_wire_743}),
            .RCLKE(),
            .RCLK(N__32055),
            .RE(N__30115),
            .WCLKE(N__20556),
            .WCLK(N__32056),
            .WE(N__30117));
    defparam \this_sprites_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,\this_sprites_ram.mem_out_bus7_3 ,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,dangling_wire_753,dangling_wire_754,\this_sprites_ram.mem_out_bus7_2 ,dangling_wire_755,dangling_wire_756,dangling_wire_757}),
            .RADDR({N__11236,N__11683,N__11575,N__11461,N__11347,N__20365,N__15523,N__15666,N__23455,N__22087,N__22281}),
            .WADDR({N__22729,N__22876,N__23023,N__24250,N__23722,N__24883,N__26173,N__28276,N__22528,N__25528,N__25972}),
            .MASK({dangling_wire_758,dangling_wire_759,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,dangling_wire_767,dangling_wire_768,dangling_wire_769,dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773}),
            .WDATA({dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,N__21091,dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,N__21202,dangling_wire_785,dangling_wire_786,dangling_wire_787}),
            .RCLKE(),
            .RCLK(N__32059),
            .RE(N__30116),
            .WCLKE(N__20563),
            .WCLK(N__32060),
            .WE(N__30118));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_788,dangling_wire_789,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,dangling_wire_797,dangling_wire_798,dangling_wire_799,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_800,dangling_wire_801,dangling_wire_802,N__18607,N__14278,N__20893,N__13963,N__14353,N__13900,N__12184,N__12625}),
            .WADDR({dangling_wire_803,dangling_wire_804,dangling_wire_805,N__15681,N__33139,N__25116,N__23596,N__23958,N__23454,N__22086,N__22284}),
            .MASK({dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,dangling_wire_811,dangling_wire_812,dangling_wire_813,dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821}),
            .WDATA({dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829,dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,N__13720,N__20635,N__19912,N__16894}),
            .RCLKE(),
            .RCLK(N__32023),
            .RE(N__30078),
            .WCLKE(N__22225),
            .WCLK(N__32024),
            .WE(N__30106));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__34841),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__34843),
            .DIN(N__34842),
            .DOUT(N__34841),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__34843),
            .PADOUT(N__34842),
            .PADIN(N__34841),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__34832),
            .DIN(N__34831),
            .DOUT(N__34830),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__34832),
            .PADOUT(N__34831),
            .PADIN(N__34830),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__34823),
            .DIN(N__34822),
            .DOUT(N__34821),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__34823),
            .PADOUT(N__34822),
            .PADIN(N__34821),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__34814),
            .DIN(N__34813),
            .DOUT(N__34812),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__34814),
            .PADOUT(N__34813),
            .PADIN(N__34812),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12025),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__34805),
            .DIN(N__34804),
            .DOUT(N__34803),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__34805),
            .PADOUT(N__34804),
            .PADIN(N__34803),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11881),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__34796),
            .DIN(N__34795),
            .DOUT(N__34794),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__34796),
            .PADOUT(N__34795),
            .PADIN(N__34794),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29934),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__34787),
            .DIN(N__34786),
            .DOUT(N__34785),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__34787),
            .PADOUT(N__34786),
            .PADIN(N__34785),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__28585),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__34778),
            .DIN(N__34777),
            .DOUT(N__34776),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__34778),
            .PADOUT(N__34777),
            .PADIN(N__34776),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__34769),
            .DIN(N__34768),
            .DOUT(N__34767),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__34769),
            .PADOUT(N__34768),
            .PADIN(N__34767),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__34760),
            .DIN(N__34759),
            .DOUT(N__34758),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__34760),
            .PADOUT(N__34759),
            .PADIN(N__34758),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__34751),
            .DIN(N__34750),
            .DOUT(N__34749),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__34751),
            .PADOUT(N__34750),
            .PADIN(N__34749),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__34742),
            .DIN(N__34741),
            .DOUT(N__34740),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__34742),
            .PADOUT(N__34741),
            .PADIN(N__34740),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__34733),
            .DIN(N__34732),
            .DOUT(N__34731),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__34733),
            .PADOUT(N__34732),
            .PADIN(N__34731),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__34724),
            .DIN(N__34723),
            .DOUT(N__34722),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__34724),
            .PADOUT(N__34723),
            .PADIN(N__34722),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__28984),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21734));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__34715),
            .DIN(N__34714),
            .DOUT(N__34713),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__34715),
            .PADOUT(N__34714),
            .PADIN(N__34713),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__30376),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21867));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__34706),
            .DIN(N__34705),
            .DOUT(N__34704),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__34706),
            .PADOUT(N__34705),
            .PADIN(N__34704),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__30316),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21839));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__34697),
            .DIN(N__34696),
            .DOUT(N__34695),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__34697),
            .PADOUT(N__34696),
            .PADIN(N__34695),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__29251),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21866));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__34688),
            .DIN(N__34687),
            .DOUT(N__34686),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__34688),
            .PADOUT(N__34687),
            .PADIN(N__34686),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__30247),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21853));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__34679),
            .DIN(N__34678),
            .DOUT(N__34677),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__34679),
            .PADOUT(N__34678),
            .PADIN(N__34677),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__28753),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21826));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__34670),
            .DIN(N__34669),
            .DOUT(N__34668),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__34670),
            .PADOUT(N__34669),
            .PADIN(N__34668),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__28708),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21743));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__34661),
            .DIN(N__34660),
            .DOUT(N__34659),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__34661),
            .PADOUT(N__34660),
            .PADIN(N__34659),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__30994),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21775));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__34652),
            .DIN(N__34651),
            .DOUT(N__34650),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__34652),
            .PADOUT(N__34651),
            .PADIN(N__34650),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__30940),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21810));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__34643),
            .DIN(N__34642),
            .DOUT(N__34641),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__34643),
            .PADOUT(N__34642),
            .PADIN(N__34641),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29305),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21871));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__34634),
            .DIN(N__34633),
            .DOUT(N__34632),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__34634),
            .PADOUT(N__34633),
            .PADIN(N__34632),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__30436),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21854));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__34625),
            .DIN(N__34624),
            .DOUT(N__34623),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__34625),
            .PADOUT(N__34624),
            .PADIN(N__34623),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__28894),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21852));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__34616),
            .DIN(N__34615),
            .DOUT(N__34614),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__34616),
            .PADOUT(N__34615),
            .PADIN(N__34614),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__28849),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21822));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__34607),
            .DIN(N__34606),
            .DOUT(N__34605),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__34607),
            .PADOUT(N__34606),
            .PADIN(N__34605),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__30205),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21865));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__34598),
            .DIN(N__34597),
            .DOUT(N__34596),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__34598),
            .PADOUT(N__34597),
            .PADIN(N__34596),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29038),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21809));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__34589),
            .DIN(N__34588),
            .DOUT(N__34587),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__34589),
            .PADOUT(N__34588),
            .PADIN(N__34587),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__30901),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21858));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__34580),
            .DIN(N__34579),
            .DOUT(N__34578),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__34580),
            .PADOUT(N__34579),
            .PADIN(N__34578),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__34571),
            .DIN(N__34570),
            .DOUT(N__34569),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__34571),
            .PADOUT(N__34570),
            .PADIN(N__34569),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__34562),
            .DIN(N__34561),
            .DOUT(N__34560),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__34562),
            .PADOUT(N__34561),
            .PADIN(N__34560),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__34553),
            .DIN(N__34552),
            .DOUT(N__34551),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__34553),
            .PADOUT(N__34552),
            .PADIN(N__34551),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__34544),
            .DIN(N__34543),
            .DOUT(N__34542),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__34544),
            .PADOUT(N__34543),
            .PADIN(N__34542),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__34535),
            .DIN(N__34534),
            .DOUT(N__34533),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__34535),
            .PADOUT(N__34534),
            .PADIN(N__34533),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__34526),
            .DIN(N__34525),
            .DOUT(N__34524),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__34526),
            .PADOUT(N__34525),
            .PADIN(N__34524),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__34517),
            .DIN(N__34516),
            .DOUT(N__34515),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__34517),
            .PADOUT(N__34516),
            .PADIN(N__34515),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__34508),
            .DIN(N__34507),
            .DOUT(N__34506),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__34508),
            .PADOUT(N__34507),
            .PADIN(N__34506),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__34499),
            .DIN(N__34498),
            .DOUT(N__34497),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__34499),
            .PADOUT(N__34498),
            .PADIN(N__34497),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11812),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__34490),
            .DIN(N__34489),
            .DOUT(N__34488),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__34490),
            .PADOUT(N__34489),
            .PADIN(N__34488),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21898),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__34481),
            .DIN(N__34480),
            .DOUT(N__34479),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__34481),
            .PADOUT(N__34480),
            .PADIN(N__34479),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__34472),
            .DIN(N__34471),
            .DOUT(N__34470),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__34472),
            .PADOUT(N__34471),
            .PADIN(N__34470),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11863),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__34463),
            .DIN(N__34462),
            .DOUT(N__34461),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__34463),
            .PADOUT(N__34462),
            .PADIN(N__34461),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__30144),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21848));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__34454),
            .DIN(N__34453),
            .DOUT(N__34452),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__34454),
            .PADOUT(N__34453),
            .PADIN(N__34452),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11797),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__34445),
            .DIN(N__34444),
            .DOUT(N__34443),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__34445),
            .PADOUT(N__34444),
            .PADIN(N__34443),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11782),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__34436),
            .DIN(N__34435),
            .DOUT(N__34434),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__34436),
            .PADOUT(N__34435),
            .PADIN(N__34434),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11917),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__34427),
            .DIN(N__34426),
            .DOUT(N__34425),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__34427),
            .PADOUT(N__34426),
            .PADIN(N__34425),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11965),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__34418),
            .DIN(N__34417),
            .DOUT(N__34416),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__34418),
            .PADOUT(N__34417),
            .PADIN(N__34416),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11950),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__34409),
            .DIN(N__34408),
            .DOUT(N__34407),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__34409),
            .PADOUT(N__34408),
            .PADIN(N__34407),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11830),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__34400),
            .DIN(N__34399),
            .DOUT(N__34398),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__34400),
            .PADOUT(N__34399),
            .PADIN(N__34398),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__34391),
            .DIN(N__34390),
            .DOUT(N__34389),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__34391),
            .PADOUT(N__34390),
            .PADIN(N__34389),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12223),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__34382),
            .DIN(N__34381),
            .DOUT(N__34380),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__34382),
            .PADOUT(N__34381),
            .PADIN(N__34380),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12469),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__8553 (
            .O(N__34363),
            .I(N__34359));
    CascadeMux I__8552 (
            .O(N__34362),
            .I(N__34354));
    InMux I__8551 (
            .O(N__34359),
            .I(N__34351));
    InMux I__8550 (
            .O(N__34358),
            .I(N__34348));
    InMux I__8549 (
            .O(N__34357),
            .I(N__34344));
    InMux I__8548 (
            .O(N__34354),
            .I(N__34340));
    LocalMux I__8547 (
            .O(N__34351),
            .I(N__34337));
    LocalMux I__8546 (
            .O(N__34348),
            .I(N__34334));
    InMux I__8545 (
            .O(N__34347),
            .I(N__34328));
    LocalMux I__8544 (
            .O(N__34344),
            .I(N__34325));
    InMux I__8543 (
            .O(N__34343),
            .I(N__34322));
    LocalMux I__8542 (
            .O(N__34340),
            .I(N__34319));
    Span4Mux_v I__8541 (
            .O(N__34337),
            .I(N__34313));
    Span4Mux_v I__8540 (
            .O(N__34334),
            .I(N__34313));
    InMux I__8539 (
            .O(N__34333),
            .I(N__34310));
    CascadeMux I__8538 (
            .O(N__34332),
            .I(N__34307));
    CascadeMux I__8537 (
            .O(N__34331),
            .I(N__34303));
    LocalMux I__8536 (
            .O(N__34328),
            .I(N__34300));
    Span4Mux_v I__8535 (
            .O(N__34325),
            .I(N__34297));
    LocalMux I__8534 (
            .O(N__34322),
            .I(N__34294));
    Span4Mux_v I__8533 (
            .O(N__34319),
            .I(N__34291));
    InMux I__8532 (
            .O(N__34318),
            .I(N__34288));
    Sp12to4 I__8531 (
            .O(N__34313),
            .I(N__34285));
    LocalMux I__8530 (
            .O(N__34310),
            .I(N__34282));
    InMux I__8529 (
            .O(N__34307),
            .I(N__34279));
    InMux I__8528 (
            .O(N__34306),
            .I(N__34274));
    InMux I__8527 (
            .O(N__34303),
            .I(N__34274));
    Sp12to4 I__8526 (
            .O(N__34300),
            .I(N__34271));
    Span4Mux_h I__8525 (
            .O(N__34297),
            .I(N__34266));
    Span4Mux_h I__8524 (
            .O(N__34294),
            .I(N__34266));
    Span4Mux_v I__8523 (
            .O(N__34291),
            .I(N__34261));
    LocalMux I__8522 (
            .O(N__34288),
            .I(N__34261));
    Span12Mux_h I__8521 (
            .O(N__34285),
            .I(N__34258));
    Span12Mux_v I__8520 (
            .O(N__34282),
            .I(N__34251));
    LocalMux I__8519 (
            .O(N__34279),
            .I(N__34251));
    LocalMux I__8518 (
            .O(N__34274),
            .I(N__34251));
    Span12Mux_h I__8517 (
            .O(N__34271),
            .I(N__34246));
    Sp12to4 I__8516 (
            .O(N__34266),
            .I(N__34246));
    Span4Mux_h I__8515 (
            .O(N__34261),
            .I(N__34243));
    Span12Mux_v I__8514 (
            .O(N__34258),
            .I(N__34240));
    Span12Mux_h I__8513 (
            .O(N__34251),
            .I(N__34237));
    Span12Mux_v I__8512 (
            .O(N__34246),
            .I(N__34234));
    Span4Mux_h I__8511 (
            .O(N__34243),
            .I(N__34231));
    Odrv12 I__8510 (
            .O(N__34240),
            .I(port_data_c_3));
    Odrv12 I__8509 (
            .O(N__34237),
            .I(port_data_c_3));
    Odrv12 I__8508 (
            .O(N__34234),
            .I(port_data_c_3));
    Odrv4 I__8507 (
            .O(N__34231),
            .I(port_data_c_3));
    CascadeMux I__8506 (
            .O(N__34222),
            .I(N__34217));
    CascadeMux I__8505 (
            .O(N__34221),
            .I(N__34214));
    CascadeMux I__8504 (
            .O(N__34220),
            .I(N__34209));
    InMux I__8503 (
            .O(N__34217),
            .I(N__34206));
    InMux I__8502 (
            .O(N__34214),
            .I(N__34203));
    CascadeMux I__8501 (
            .O(N__34213),
            .I(N__34199));
    InMux I__8500 (
            .O(N__34212),
            .I(N__34196));
    InMux I__8499 (
            .O(N__34209),
            .I(N__34193));
    LocalMux I__8498 (
            .O(N__34206),
            .I(N__34189));
    LocalMux I__8497 (
            .O(N__34203),
            .I(N__34186));
    CascadeMux I__8496 (
            .O(N__34202),
            .I(N__34183));
    InMux I__8495 (
            .O(N__34199),
            .I(N__34180));
    LocalMux I__8494 (
            .O(N__34196),
            .I(N__34177));
    LocalMux I__8493 (
            .O(N__34193),
            .I(N__34174));
    InMux I__8492 (
            .O(N__34192),
            .I(N__34171));
    Span4Mux_v I__8491 (
            .O(N__34189),
            .I(N__34166));
    Span4Mux_v I__8490 (
            .O(N__34186),
            .I(N__34166));
    InMux I__8489 (
            .O(N__34183),
            .I(N__34163));
    LocalMux I__8488 (
            .O(N__34180),
            .I(N__34160));
    Span4Mux_h I__8487 (
            .O(N__34177),
            .I(N__34155));
    Span4Mux_v I__8486 (
            .O(N__34174),
            .I(N__34155));
    LocalMux I__8485 (
            .O(N__34171),
            .I(N__34152));
    Span4Mux_h I__8484 (
            .O(N__34166),
            .I(N__34145));
    LocalMux I__8483 (
            .O(N__34163),
            .I(N__34145));
    Span4Mux_v I__8482 (
            .O(N__34160),
            .I(N__34141));
    Span4Mux_h I__8481 (
            .O(N__34155),
            .I(N__34136));
    Span4Mux_v I__8480 (
            .O(N__34152),
            .I(N__34136));
    InMux I__8479 (
            .O(N__34151),
            .I(N__34133));
    CascadeMux I__8478 (
            .O(N__34150),
            .I(N__34130));
    Span4Mux_h I__8477 (
            .O(N__34145),
            .I(N__34126));
    InMux I__8476 (
            .O(N__34144),
            .I(N__34123));
    Sp12to4 I__8475 (
            .O(N__34141),
            .I(N__34120));
    Span4Mux_h I__8474 (
            .O(N__34136),
            .I(N__34115));
    LocalMux I__8473 (
            .O(N__34133),
            .I(N__34115));
    InMux I__8472 (
            .O(N__34130),
            .I(N__34112));
    InMux I__8471 (
            .O(N__34129),
            .I(N__34109));
    Span4Mux_v I__8470 (
            .O(N__34126),
            .I(N__34106));
    LocalMux I__8469 (
            .O(N__34123),
            .I(N__34103));
    Span12Mux_h I__8468 (
            .O(N__34120),
            .I(N__34100));
    Sp12to4 I__8467 (
            .O(N__34115),
            .I(N__34097));
    LocalMux I__8466 (
            .O(N__34112),
            .I(N__34092));
    LocalMux I__8465 (
            .O(N__34109),
            .I(N__34092));
    Span4Mux_v I__8464 (
            .O(N__34106),
            .I(N__34087));
    Span4Mux_h I__8463 (
            .O(N__34103),
            .I(N__34087));
    Span12Mux_v I__8462 (
            .O(N__34100),
            .I(N__34084));
    Span12Mux_v I__8461 (
            .O(N__34097),
            .I(N__34081));
    Span12Mux_h I__8460 (
            .O(N__34092),
            .I(N__34078));
    Span4Mux_v I__8459 (
            .O(N__34087),
            .I(N__34075));
    Odrv12 I__8458 (
            .O(N__34084),
            .I(port_data_c_2));
    Odrv12 I__8457 (
            .O(N__34081),
            .I(port_data_c_2));
    Odrv12 I__8456 (
            .O(N__34078),
            .I(port_data_c_2));
    Odrv4 I__8455 (
            .O(N__34075),
            .I(port_data_c_2));
    CascadeMux I__8454 (
            .O(N__34066),
            .I(\this_vga_signals.M_this_external_address_d21Z0Z_2_cascade_ ));
    CascadeMux I__8453 (
            .O(N__34063),
            .I(N__34060));
    InMux I__8452 (
            .O(N__34060),
            .I(N__34054));
    CascadeMux I__8451 (
            .O(N__34059),
            .I(N__34051));
    InMux I__8450 (
            .O(N__34058),
            .I(N__34047));
    InMux I__8449 (
            .O(N__34057),
            .I(N__34044));
    LocalMux I__8448 (
            .O(N__34054),
            .I(N__34041));
    InMux I__8447 (
            .O(N__34051),
            .I(N__34038));
    CascadeMux I__8446 (
            .O(N__34050),
            .I(N__34035));
    LocalMux I__8445 (
            .O(N__34047),
            .I(N__34032));
    LocalMux I__8444 (
            .O(N__34044),
            .I(N__34029));
    Span4Mux_h I__8443 (
            .O(N__34041),
            .I(N__34024));
    LocalMux I__8442 (
            .O(N__34038),
            .I(N__34024));
    InMux I__8441 (
            .O(N__34035),
            .I(N__34021));
    Span12Mux_h I__8440 (
            .O(N__34032),
            .I(N__34018));
    Span12Mux_h I__8439 (
            .O(N__34029),
            .I(N__34015));
    Span4Mux_h I__8438 (
            .O(N__34024),
            .I(N__34012));
    LocalMux I__8437 (
            .O(N__34021),
            .I(N__34009));
    Odrv12 I__8436 (
            .O(N__34018),
            .I(\this_vga_signals.M_this_external_address_dZ0Z21 ));
    Odrv12 I__8435 (
            .O(N__34015),
            .I(\this_vga_signals.M_this_external_address_dZ0Z21 ));
    Odrv4 I__8434 (
            .O(N__34012),
            .I(\this_vga_signals.M_this_external_address_dZ0Z21 ));
    Odrv12 I__8433 (
            .O(N__34009),
            .I(\this_vga_signals.M_this_external_address_dZ0Z21 ));
    InMux I__8432 (
            .O(N__34000),
            .I(N__33996));
    InMux I__8431 (
            .O(N__33999),
            .I(N__33993));
    LocalMux I__8430 (
            .O(N__33996),
            .I(N__33986));
    LocalMux I__8429 (
            .O(N__33993),
            .I(N__33983));
    CascadeMux I__8428 (
            .O(N__33992),
            .I(N__33978));
    CascadeMux I__8427 (
            .O(N__33991),
            .I(N__33975));
    CascadeMux I__8426 (
            .O(N__33990),
            .I(N__33972));
    InMux I__8425 (
            .O(N__33989),
            .I(N__33967));
    Span4Mux_h I__8424 (
            .O(N__33986),
            .I(N__33961));
    Span4Mux_v I__8423 (
            .O(N__33983),
            .I(N__33961));
    InMux I__8422 (
            .O(N__33982),
            .I(N__33958));
    CascadeMux I__8421 (
            .O(N__33981),
            .I(N__33955));
    InMux I__8420 (
            .O(N__33978),
            .I(N__33952));
    InMux I__8419 (
            .O(N__33975),
            .I(N__33949));
    InMux I__8418 (
            .O(N__33972),
            .I(N__33946));
    InMux I__8417 (
            .O(N__33971),
            .I(N__33940));
    InMux I__8416 (
            .O(N__33970),
            .I(N__33940));
    LocalMux I__8415 (
            .O(N__33967),
            .I(N__33937));
    CascadeMux I__8414 (
            .O(N__33966),
            .I(N__33934));
    Span4Mux_h I__8413 (
            .O(N__33961),
            .I(N__33929));
    LocalMux I__8412 (
            .O(N__33958),
            .I(N__33929));
    InMux I__8411 (
            .O(N__33955),
            .I(N__33926));
    LocalMux I__8410 (
            .O(N__33952),
            .I(N__33923));
    LocalMux I__8409 (
            .O(N__33949),
            .I(N__33918));
    LocalMux I__8408 (
            .O(N__33946),
            .I(N__33918));
    InMux I__8407 (
            .O(N__33945),
            .I(N__33915));
    LocalMux I__8406 (
            .O(N__33940),
            .I(N__33912));
    Span4Mux_v I__8405 (
            .O(N__33937),
            .I(N__33909));
    InMux I__8404 (
            .O(N__33934),
            .I(N__33906));
    Span4Mux_h I__8403 (
            .O(N__33929),
            .I(N__33901));
    LocalMux I__8402 (
            .O(N__33926),
            .I(N__33901));
    Span4Mux_v I__8401 (
            .O(N__33923),
            .I(N__33898));
    Span4Mux_v I__8400 (
            .O(N__33918),
            .I(N__33895));
    LocalMux I__8399 (
            .O(N__33915),
            .I(N__33892));
    Span12Mux_s7_h I__8398 (
            .O(N__33912),
            .I(N__33885));
    Sp12to4 I__8397 (
            .O(N__33909),
            .I(N__33885));
    LocalMux I__8396 (
            .O(N__33906),
            .I(N__33885));
    Span4Mux_v I__8395 (
            .O(N__33901),
            .I(N__33882));
    Span4Mux_v I__8394 (
            .O(N__33898),
            .I(N__33875));
    Span4Mux_v I__8393 (
            .O(N__33895),
            .I(N__33875));
    Span4Mux_v I__8392 (
            .O(N__33892),
            .I(N__33875));
    Span12Mux_h I__8391 (
            .O(N__33885),
            .I(N__33872));
    Span4Mux_h I__8390 (
            .O(N__33882),
            .I(N__33869));
    Sp12to4 I__8389 (
            .O(N__33875),
            .I(N__33866));
    Span12Mux_v I__8388 (
            .O(N__33872),
            .I(N__33863));
    Sp12to4 I__8387 (
            .O(N__33869),
            .I(N__33860));
    Span12Mux_h I__8386 (
            .O(N__33866),
            .I(N__33857));
    Odrv12 I__8385 (
            .O(N__33863),
            .I(port_data_c_1));
    Odrv12 I__8384 (
            .O(N__33860),
            .I(port_data_c_1));
    Odrv12 I__8383 (
            .O(N__33857),
            .I(port_data_c_1));
    CascadeMux I__8382 (
            .O(N__33850),
            .I(N__33847));
    InMux I__8381 (
            .O(N__33847),
            .I(N__33844));
    LocalMux I__8380 (
            .O(N__33844),
            .I(\this_vga_signals.M_this_external_address_d21Z0Z_2 ));
    CascadeMux I__8379 (
            .O(N__33841),
            .I(N__33838));
    InMux I__8378 (
            .O(N__33838),
            .I(N__33832));
    CascadeMux I__8377 (
            .O(N__33837),
            .I(N__33829));
    CascadeMux I__8376 (
            .O(N__33836),
            .I(N__33824));
    InMux I__8375 (
            .O(N__33835),
            .I(N__33819));
    LocalMux I__8374 (
            .O(N__33832),
            .I(N__33815));
    InMux I__8373 (
            .O(N__33829),
            .I(N__33808));
    InMux I__8372 (
            .O(N__33828),
            .I(N__33808));
    InMux I__8371 (
            .O(N__33827),
            .I(N__33803));
    InMux I__8370 (
            .O(N__33824),
            .I(N__33803));
    InMux I__8369 (
            .O(N__33823),
            .I(N__33798));
    InMux I__8368 (
            .O(N__33822),
            .I(N__33798));
    LocalMux I__8367 (
            .O(N__33819),
            .I(N__33795));
    InMux I__8366 (
            .O(N__33818),
            .I(N__33791));
    Span4Mux_v I__8365 (
            .O(N__33815),
            .I(N__33788));
    InMux I__8364 (
            .O(N__33814),
            .I(N__33785));
    InMux I__8363 (
            .O(N__33813),
            .I(N__33782));
    LocalMux I__8362 (
            .O(N__33808),
            .I(N__33779));
    LocalMux I__8361 (
            .O(N__33803),
            .I(N__33776));
    LocalMux I__8360 (
            .O(N__33798),
            .I(N__33773));
    Span4Mux_v I__8359 (
            .O(N__33795),
            .I(N__33770));
    InMux I__8358 (
            .O(N__33794),
            .I(N__33767));
    LocalMux I__8357 (
            .O(N__33791),
            .I(N__33764));
    Span4Mux_v I__8356 (
            .O(N__33788),
            .I(N__33761));
    LocalMux I__8355 (
            .O(N__33785),
            .I(N__33758));
    LocalMux I__8354 (
            .O(N__33782),
            .I(N__33755));
    Span4Mux_v I__8353 (
            .O(N__33779),
            .I(N__33752));
    Span4Mux_v I__8352 (
            .O(N__33776),
            .I(N__33749));
    Sp12to4 I__8351 (
            .O(N__33773),
            .I(N__33742));
    Sp12to4 I__8350 (
            .O(N__33770),
            .I(N__33742));
    LocalMux I__8349 (
            .O(N__33767),
            .I(N__33742));
    Span4Mux_h I__8348 (
            .O(N__33764),
            .I(N__33739));
    Span4Mux_v I__8347 (
            .O(N__33761),
            .I(N__33736));
    Span4Mux_v I__8346 (
            .O(N__33758),
            .I(N__33733));
    Span12Mux_h I__8345 (
            .O(N__33755),
            .I(N__33730));
    Sp12to4 I__8344 (
            .O(N__33752),
            .I(N__33725));
    Sp12to4 I__8343 (
            .O(N__33749),
            .I(N__33725));
    Span12Mux_h I__8342 (
            .O(N__33742),
            .I(N__33720));
    Sp12to4 I__8341 (
            .O(N__33739),
            .I(N__33720));
    Sp12to4 I__8340 (
            .O(N__33736),
            .I(N__33715));
    Sp12to4 I__8339 (
            .O(N__33733),
            .I(N__33715));
    Span12Mux_v I__8338 (
            .O(N__33730),
            .I(N__33712));
    Span12Mux_h I__8337 (
            .O(N__33725),
            .I(N__33709));
    Span12Mux_v I__8336 (
            .O(N__33720),
            .I(N__33704));
    Span12Mux_h I__8335 (
            .O(N__33715),
            .I(N__33704));
    Odrv12 I__8334 (
            .O(N__33712),
            .I(port_data_c_0));
    Odrv12 I__8333 (
            .O(N__33709),
            .I(port_data_c_0));
    Odrv12 I__8332 (
            .O(N__33704),
            .I(port_data_c_0));
    CascadeMux I__8331 (
            .O(N__33697),
            .I(N__33694));
    InMux I__8330 (
            .O(N__33694),
            .I(N__33689));
    InMux I__8329 (
            .O(N__33693),
            .I(N__33686));
    InMux I__8328 (
            .O(N__33692),
            .I(N__33683));
    LocalMux I__8327 (
            .O(N__33689),
            .I(N__33679));
    LocalMux I__8326 (
            .O(N__33686),
            .I(N__33676));
    LocalMux I__8325 (
            .O(N__33683),
            .I(N__33673));
    InMux I__8324 (
            .O(N__33682),
            .I(N__33670));
    Span4Mux_v I__8323 (
            .O(N__33679),
            .I(N__33665));
    Span4Mux_v I__8322 (
            .O(N__33676),
            .I(N__33665));
    Span4Mux_v I__8321 (
            .O(N__33673),
            .I(N__33662));
    LocalMux I__8320 (
            .O(N__33670),
            .I(N__33659));
    Span4Mux_h I__8319 (
            .O(N__33665),
            .I(N__33656));
    Span4Mux_h I__8318 (
            .O(N__33662),
            .I(N__33651));
    Span4Mux_v I__8317 (
            .O(N__33659),
            .I(N__33651));
    Odrv4 I__8316 (
            .O(N__33656),
            .I(\this_vga_signals.M_this_external_address_dZ0Z22 ));
    Odrv4 I__8315 (
            .O(N__33651),
            .I(\this_vga_signals.M_this_external_address_dZ0Z22 ));
    CascadeMux I__8314 (
            .O(N__33646),
            .I(N__33643));
    InMux I__8313 (
            .O(N__33643),
            .I(N__33638));
    CascadeMux I__8312 (
            .O(N__33642),
            .I(N__33634));
    CascadeMux I__8311 (
            .O(N__33641),
            .I(N__33631));
    LocalMux I__8310 (
            .O(N__33638),
            .I(N__33627));
    InMux I__8309 (
            .O(N__33637),
            .I(N__33624));
    InMux I__8308 (
            .O(N__33634),
            .I(N__33621));
    InMux I__8307 (
            .O(N__33631),
            .I(N__33618));
    InMux I__8306 (
            .O(N__33630),
            .I(N__33615));
    Span4Mux_h I__8305 (
            .O(N__33627),
            .I(N__33608));
    LocalMux I__8304 (
            .O(N__33624),
            .I(N__33608));
    LocalMux I__8303 (
            .O(N__33621),
            .I(N__33605));
    LocalMux I__8302 (
            .O(N__33618),
            .I(N__33602));
    LocalMux I__8301 (
            .O(N__33615),
            .I(N__33599));
    InMux I__8300 (
            .O(N__33614),
            .I(N__33596));
    InMux I__8299 (
            .O(N__33613),
            .I(N__33592));
    Span4Mux_h I__8298 (
            .O(N__33608),
            .I(N__33589));
    Span4Mux_v I__8297 (
            .O(N__33605),
            .I(N__33582));
    Span4Mux_v I__8296 (
            .O(N__33602),
            .I(N__33582));
    Span4Mux_v I__8295 (
            .O(N__33599),
            .I(N__33582));
    LocalMux I__8294 (
            .O(N__33596),
            .I(N__33579));
    InMux I__8293 (
            .O(N__33595),
            .I(N__33575));
    LocalMux I__8292 (
            .O(N__33592),
            .I(N__33572));
    Span4Mux_v I__8291 (
            .O(N__33589),
            .I(N__33565));
    Span4Mux_h I__8290 (
            .O(N__33582),
            .I(N__33565));
    Span4Mux_v I__8289 (
            .O(N__33579),
            .I(N__33565));
    InMux I__8288 (
            .O(N__33578),
            .I(N__33562));
    LocalMux I__8287 (
            .O(N__33575),
            .I(N__33559));
    Span12Mux_h I__8286 (
            .O(N__33572),
            .I(N__33556));
    Sp12to4 I__8285 (
            .O(N__33565),
            .I(N__33551));
    LocalMux I__8284 (
            .O(N__33562),
            .I(N__33551));
    Span12Mux_v I__8283 (
            .O(N__33559),
            .I(N__33548));
    Span12Mux_v I__8282 (
            .O(N__33556),
            .I(N__33543));
    Span12Mux_h I__8281 (
            .O(N__33551),
            .I(N__33543));
    Odrv12 I__8280 (
            .O(N__33548),
            .I(port_data_c_5));
    Odrv12 I__8279 (
            .O(N__33543),
            .I(port_data_c_5));
    CascadeMux I__8278 (
            .O(N__33538),
            .I(N__33533));
    InMux I__8277 (
            .O(N__33537),
            .I(N__33529));
    CascadeMux I__8276 (
            .O(N__33536),
            .I(N__33526));
    InMux I__8275 (
            .O(N__33533),
            .I(N__33523));
    CascadeMux I__8274 (
            .O(N__33532),
            .I(N__33520));
    LocalMux I__8273 (
            .O(N__33529),
            .I(N__33516));
    InMux I__8272 (
            .O(N__33526),
            .I(N__33513));
    LocalMux I__8271 (
            .O(N__33523),
            .I(N__33509));
    InMux I__8270 (
            .O(N__33520),
            .I(N__33505));
    InMux I__8269 (
            .O(N__33519),
            .I(N__33502));
    Span4Mux_v I__8268 (
            .O(N__33516),
            .I(N__33497));
    LocalMux I__8267 (
            .O(N__33513),
            .I(N__33497));
    InMux I__8266 (
            .O(N__33512),
            .I(N__33493));
    Span4Mux_v I__8265 (
            .O(N__33509),
            .I(N__33490));
    InMux I__8264 (
            .O(N__33508),
            .I(N__33487));
    LocalMux I__8263 (
            .O(N__33505),
            .I(N__33484));
    LocalMux I__8262 (
            .O(N__33502),
            .I(N__33481));
    Span4Mux_v I__8261 (
            .O(N__33497),
            .I(N__33477));
    InMux I__8260 (
            .O(N__33496),
            .I(N__33474));
    LocalMux I__8259 (
            .O(N__33493),
            .I(N__33471));
    Span4Mux_v I__8258 (
            .O(N__33490),
            .I(N__33468));
    LocalMux I__8257 (
            .O(N__33487),
            .I(N__33465));
    Span4Mux_h I__8256 (
            .O(N__33484),
            .I(N__33460));
    Span4Mux_h I__8255 (
            .O(N__33481),
            .I(N__33460));
    InMux I__8254 (
            .O(N__33480),
            .I(N__33457));
    Span4Mux_h I__8253 (
            .O(N__33477),
            .I(N__33452));
    LocalMux I__8252 (
            .O(N__33474),
            .I(N__33452));
    Span12Mux_v I__8251 (
            .O(N__33471),
            .I(N__33447));
    Sp12to4 I__8250 (
            .O(N__33468),
            .I(N__33447));
    Span12Mux_s9_v I__8249 (
            .O(N__33465),
            .I(N__33438));
    Sp12to4 I__8248 (
            .O(N__33460),
            .I(N__33438));
    LocalMux I__8247 (
            .O(N__33457),
            .I(N__33438));
    Sp12to4 I__8246 (
            .O(N__33452),
            .I(N__33438));
    Span12Mux_h I__8245 (
            .O(N__33447),
            .I(N__33435));
    Span12Mux_v I__8244 (
            .O(N__33438),
            .I(N__33432));
    Odrv12 I__8243 (
            .O(N__33435),
            .I(port_data_c_6));
    Odrv12 I__8242 (
            .O(N__33432),
            .I(port_data_c_6));
    CascadeMux I__8241 (
            .O(N__33427),
            .I(N__33423));
    CascadeMux I__8240 (
            .O(N__33426),
            .I(N__33418));
    InMux I__8239 (
            .O(N__33423),
            .I(N__33415));
    InMux I__8238 (
            .O(N__33422),
            .I(N__33412));
    InMux I__8237 (
            .O(N__33421),
            .I(N__33407));
    InMux I__8236 (
            .O(N__33418),
            .I(N__33407));
    LocalMux I__8235 (
            .O(N__33415),
            .I(N__33403));
    LocalMux I__8234 (
            .O(N__33412),
            .I(N__33400));
    LocalMux I__8233 (
            .O(N__33407),
            .I(N__33397));
    InMux I__8232 (
            .O(N__33406),
            .I(N__33394));
    Span4Mux_v I__8231 (
            .O(N__33403),
            .I(N__33391));
    Span4Mux_v I__8230 (
            .O(N__33400),
            .I(N__33382));
    Span4Mux_h I__8229 (
            .O(N__33397),
            .I(N__33382));
    LocalMux I__8228 (
            .O(N__33394),
            .I(N__33382));
    Span4Mux_h I__8227 (
            .O(N__33391),
            .I(N__33379));
    InMux I__8226 (
            .O(N__33390),
            .I(N__33376));
    CascadeMux I__8225 (
            .O(N__33389),
            .I(N__33373));
    Span4Mux_v I__8224 (
            .O(N__33382),
            .I(N__33370));
    Span4Mux_h I__8223 (
            .O(N__33379),
            .I(N__33365));
    LocalMux I__8222 (
            .O(N__33376),
            .I(N__33365));
    InMux I__8221 (
            .O(N__33373),
            .I(N__33362));
    Span4Mux_v I__8220 (
            .O(N__33370),
            .I(N__33357));
    Span4Mux_v I__8219 (
            .O(N__33365),
            .I(N__33357));
    LocalMux I__8218 (
            .O(N__33362),
            .I(N__33354));
    Span4Mux_h I__8217 (
            .O(N__33357),
            .I(N__33351));
    Span12Mux_v I__8216 (
            .O(N__33354),
            .I(N__33348));
    IoSpan4Mux I__8215 (
            .O(N__33351),
            .I(N__33345));
    Odrv12 I__8214 (
            .O(N__33348),
            .I(port_data_c_7));
    Odrv4 I__8213 (
            .O(N__33345),
            .I(port_data_c_7));
    CascadeMux I__8212 (
            .O(N__33340),
            .I(N__33337));
    InMux I__8211 (
            .O(N__33337),
            .I(N__33333));
    CascadeMux I__8210 (
            .O(N__33336),
            .I(N__33330));
    LocalMux I__8209 (
            .O(N__33333),
            .I(N__33323));
    InMux I__8208 (
            .O(N__33330),
            .I(N__33320));
    CascadeMux I__8207 (
            .O(N__33329),
            .I(N__33316));
    CascadeMux I__8206 (
            .O(N__33328),
            .I(N__33313));
    InMux I__8205 (
            .O(N__33327),
            .I(N__33308));
    CascadeMux I__8204 (
            .O(N__33326),
            .I(N__33305));
    Span4Mux_v I__8203 (
            .O(N__33323),
            .I(N__33300));
    LocalMux I__8202 (
            .O(N__33320),
            .I(N__33300));
    InMux I__8201 (
            .O(N__33319),
            .I(N__33297));
    InMux I__8200 (
            .O(N__33316),
            .I(N__33294));
    InMux I__8199 (
            .O(N__33313),
            .I(N__33291));
    InMux I__8198 (
            .O(N__33312),
            .I(N__33288));
    CascadeMux I__8197 (
            .O(N__33311),
            .I(N__33285));
    LocalMux I__8196 (
            .O(N__33308),
            .I(N__33282));
    InMux I__8195 (
            .O(N__33305),
            .I(N__33279));
    Span4Mux_h I__8194 (
            .O(N__33300),
            .I(N__33270));
    LocalMux I__8193 (
            .O(N__33297),
            .I(N__33270));
    LocalMux I__8192 (
            .O(N__33294),
            .I(N__33270));
    LocalMux I__8191 (
            .O(N__33291),
            .I(N__33270));
    LocalMux I__8190 (
            .O(N__33288),
            .I(N__33267));
    InMux I__8189 (
            .O(N__33285),
            .I(N__33263));
    Span4Mux_v I__8188 (
            .O(N__33282),
            .I(N__33258));
    LocalMux I__8187 (
            .O(N__33279),
            .I(N__33258));
    Span4Mux_v I__8186 (
            .O(N__33270),
            .I(N__33255));
    Span4Mux_v I__8185 (
            .O(N__33267),
            .I(N__33252));
    InMux I__8184 (
            .O(N__33266),
            .I(N__33249));
    LocalMux I__8183 (
            .O(N__33263),
            .I(N__33245));
    Span4Mux_v I__8182 (
            .O(N__33258),
            .I(N__33242));
    Span4Mux_h I__8181 (
            .O(N__33255),
            .I(N__33237));
    Span4Mux_v I__8180 (
            .O(N__33252),
            .I(N__33237));
    LocalMux I__8179 (
            .O(N__33249),
            .I(N__33234));
    InMux I__8178 (
            .O(N__33248),
            .I(N__33231));
    Span12Mux_v I__8177 (
            .O(N__33245),
            .I(N__33228));
    Span4Mux_v I__8176 (
            .O(N__33242),
            .I(N__33225));
    Span4Mux_v I__8175 (
            .O(N__33237),
            .I(N__33220));
    Span4Mux_v I__8174 (
            .O(N__33234),
            .I(N__33220));
    LocalMux I__8173 (
            .O(N__33231),
            .I(N__33217));
    Span12Mux_h I__8172 (
            .O(N__33228),
            .I(N__33214));
    Sp12to4 I__8171 (
            .O(N__33225),
            .I(N__33211));
    Sp12to4 I__8170 (
            .O(N__33220),
            .I(N__33206));
    Span12Mux_v I__8169 (
            .O(N__33217),
            .I(N__33206));
    Odrv12 I__8168 (
            .O(N__33214),
            .I(port_data_c_4));
    Odrv12 I__8167 (
            .O(N__33211),
            .I(port_data_c_4));
    Odrv12 I__8166 (
            .O(N__33206),
            .I(port_data_c_4));
    InMux I__8165 (
            .O(N__33199),
            .I(N__33193));
    InMux I__8164 (
            .O(N__33198),
            .I(N__33193));
    LocalMux I__8163 (
            .O(N__33193),
            .I(N__33190));
    Odrv4 I__8162 (
            .O(N__33190),
            .I(\this_vga_signals.M_this_external_address_d21Z0Z_6 ));
    InMux I__8161 (
            .O(N__33187),
            .I(N__33184));
    LocalMux I__8160 (
            .O(N__33184),
            .I(N__33181));
    Span4Mux_v I__8159 (
            .O(N__33181),
            .I(N__33178));
    Odrv4 I__8158 (
            .O(N__33178),
            .I(M_this_map_ram_write_data_7));
    InMux I__8157 (
            .O(N__33175),
            .I(N__33171));
    InMux I__8156 (
            .O(N__33174),
            .I(N__33168));
    LocalMux I__8155 (
            .O(N__33171),
            .I(N__33165));
    LocalMux I__8154 (
            .O(N__33168),
            .I(\this_ppu.M_haddress_qZ0Z_7 ));
    Odrv12 I__8153 (
            .O(N__33165),
            .I(\this_ppu.M_haddress_qZ0Z_7 ));
    CascadeMux I__8152 (
            .O(N__33160),
            .I(N__33157));
    CascadeBuf I__8151 (
            .O(N__33157),
            .I(N__33154));
    CascadeMux I__8150 (
            .O(N__33154),
            .I(N__33151));
    InMux I__8149 (
            .O(N__33151),
            .I(N__33148));
    LocalMux I__8148 (
            .O(N__33148),
            .I(N__33145));
    Span4Mux_v I__8147 (
            .O(N__33145),
            .I(N__33142));
    Odrv4 I__8146 (
            .O(N__33142),
            .I(M_this_ppu_map_addr_4));
    CascadeMux I__8145 (
            .O(N__33139),
            .I(N__33136));
    InMux I__8144 (
            .O(N__33136),
            .I(N__33133));
    LocalMux I__8143 (
            .O(N__33133),
            .I(N__33130));
    Span4Mux_h I__8142 (
            .O(N__33130),
            .I(N__33127));
    Span4Mux_v I__8141 (
            .O(N__33127),
            .I(N__33122));
    InMux I__8140 (
            .O(N__33126),
            .I(N__33117));
    InMux I__8139 (
            .O(N__33125),
            .I(N__33117));
    Span4Mux_v I__8138 (
            .O(N__33122),
            .I(N__33110));
    LocalMux I__8137 (
            .O(N__33117),
            .I(N__33110));
    InMux I__8136 (
            .O(N__33116),
            .I(N__33107));
    InMux I__8135 (
            .O(N__33115),
            .I(N__33104));
    Span4Mux_h I__8134 (
            .O(N__33110),
            .I(N__33101));
    LocalMux I__8133 (
            .O(N__33107),
            .I(M_this_ppu_vram_addr_6));
    LocalMux I__8132 (
            .O(N__33104),
            .I(M_this_ppu_vram_addr_6));
    Odrv4 I__8131 (
            .O(N__33101),
            .I(M_this_ppu_vram_addr_6));
    CascadeMux I__8130 (
            .O(N__33094),
            .I(N__33091));
    CascadeBuf I__8129 (
            .O(N__33091),
            .I(N__33088));
    CascadeMux I__8128 (
            .O(N__33088),
            .I(N__33085));
    InMux I__8127 (
            .O(N__33085),
            .I(N__33082));
    LocalMux I__8126 (
            .O(N__33082),
            .I(N__33079));
    Span4Mux_s3_v I__8125 (
            .O(N__33079),
            .I(N__33076));
    Odrv4 I__8124 (
            .O(N__33076),
            .I(M_this_ppu_vram_addr_i_6));
    InMux I__8123 (
            .O(N__33073),
            .I(N__33070));
    LocalMux I__8122 (
            .O(N__33070),
            .I(M_this_map_ram_write_data_2));
    InMux I__8121 (
            .O(N__33067),
            .I(N__33064));
    LocalMux I__8120 (
            .O(N__33064),
            .I(N__33061));
    Odrv4 I__8119 (
            .O(N__33061),
            .I(M_this_map_ram_write_data_1));
    InMux I__8118 (
            .O(N__33058),
            .I(N__33055));
    LocalMux I__8117 (
            .O(N__33055),
            .I(M_this_map_ram_write_data_0));
    InMux I__8116 (
            .O(N__33052),
            .I(N__33049));
    LocalMux I__8115 (
            .O(N__33049),
            .I(M_this_map_ram_write_data_5));
    CascadeMux I__8114 (
            .O(N__33046),
            .I(N__33040));
    CEMux I__8113 (
            .O(N__33045),
            .I(N__33036));
    CEMux I__8112 (
            .O(N__33044),
            .I(N__33033));
    InMux I__8111 (
            .O(N__33043),
            .I(N__33030));
    InMux I__8110 (
            .O(N__33040),
            .I(N__33025));
    InMux I__8109 (
            .O(N__33039),
            .I(N__33025));
    LocalMux I__8108 (
            .O(N__33036),
            .I(N__33019));
    LocalMux I__8107 (
            .O(N__33033),
            .I(N__33012));
    LocalMux I__8106 (
            .O(N__33030),
            .I(N__33012));
    LocalMux I__8105 (
            .O(N__33025),
            .I(N__33012));
    InMux I__8104 (
            .O(N__33024),
            .I(N__33007));
    InMux I__8103 (
            .O(N__33023),
            .I(N__33007));
    InMux I__8102 (
            .O(N__33022),
            .I(N__33002));
    Span4Mux_v I__8101 (
            .O(N__33019),
            .I(N__32994));
    Span4Mux_v I__8100 (
            .O(N__33012),
            .I(N__32994));
    LocalMux I__8099 (
            .O(N__33007),
            .I(N__32994));
    InMux I__8098 (
            .O(N__33006),
            .I(N__32989));
    InMux I__8097 (
            .O(N__33005),
            .I(N__32989));
    LocalMux I__8096 (
            .O(N__33002),
            .I(N__32986));
    InMux I__8095 (
            .O(N__33001),
            .I(N__32981));
    Span4Mux_h I__8094 (
            .O(N__32994),
            .I(N__32978));
    LocalMux I__8093 (
            .O(N__32989),
            .I(N__32975));
    Span12Mux_h I__8092 (
            .O(N__32986),
            .I(N__32972));
    InMux I__8091 (
            .O(N__32985),
            .I(N__32967));
    InMux I__8090 (
            .O(N__32984),
            .I(N__32967));
    LocalMux I__8089 (
            .O(N__32981),
            .I(N__32960));
    Span4Mux_v I__8088 (
            .O(N__32978),
            .I(N__32960));
    Span4Mux_h I__8087 (
            .O(N__32975),
            .I(N__32960));
    Span12Mux_v I__8086 (
            .O(N__32972),
            .I(N__32957));
    LocalMux I__8085 (
            .O(N__32967),
            .I(N__32952));
    Span4Mux_v I__8084 (
            .O(N__32960),
            .I(N__32952));
    Odrv12 I__8083 (
            .O(N__32957),
            .I(M_this_map_ram_write_en_0));
    Odrv4 I__8082 (
            .O(N__32952),
            .I(M_this_map_ram_write_en_0));
    InMux I__8081 (
            .O(N__32947),
            .I(N__32944));
    LocalMux I__8080 (
            .O(N__32944),
            .I(M_this_map_ram_write_data_4));
    InMux I__8079 (
            .O(N__32941),
            .I(N__32938));
    LocalMux I__8078 (
            .O(N__32938),
            .I(M_this_data_count_q_cry_9_THRU_CO));
    CascadeMux I__8077 (
            .O(N__32935),
            .I(M_this_data_count_q_3_10_cascade_));
    CascadeMux I__8076 (
            .O(N__32932),
            .I(N__32926));
    InMux I__8075 (
            .O(N__32931),
            .I(N__32920));
    InMux I__8074 (
            .O(N__32930),
            .I(N__32917));
    InMux I__8073 (
            .O(N__32929),
            .I(N__32913));
    InMux I__8072 (
            .O(N__32926),
            .I(N__32910));
    InMux I__8071 (
            .O(N__32925),
            .I(N__32907));
    InMux I__8070 (
            .O(N__32924),
            .I(N__32904));
    InMux I__8069 (
            .O(N__32923),
            .I(N__32901));
    LocalMux I__8068 (
            .O(N__32920),
            .I(N__32898));
    LocalMux I__8067 (
            .O(N__32917),
            .I(N__32895));
    InMux I__8066 (
            .O(N__32916),
            .I(N__32892));
    LocalMux I__8065 (
            .O(N__32913),
            .I(N__32889));
    LocalMux I__8064 (
            .O(N__32910),
            .I(N__32886));
    LocalMux I__8063 (
            .O(N__32907),
            .I(N__32883));
    LocalMux I__8062 (
            .O(N__32904),
            .I(N__32880));
    LocalMux I__8061 (
            .O(N__32901),
            .I(N__32877));
    Span4Mux_h I__8060 (
            .O(N__32898),
            .I(N__32872));
    Span4Mux_h I__8059 (
            .O(N__32895),
            .I(N__32872));
    LocalMux I__8058 (
            .O(N__32892),
            .I(N__32861));
    Span4Mux_v I__8057 (
            .O(N__32889),
            .I(N__32861));
    Span4Mux_v I__8056 (
            .O(N__32886),
            .I(N__32861));
    Span4Mux_v I__8055 (
            .O(N__32883),
            .I(N__32861));
    Span4Mux_h I__8054 (
            .O(N__32880),
            .I(N__32861));
    Odrv12 I__8053 (
            .O(N__32877),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__8052 (
            .O(N__32872),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__8051 (
            .O(N__32861),
            .I(M_this_state_qZ0Z_8));
    InMux I__8050 (
            .O(N__32854),
            .I(N__32840));
    InMux I__8049 (
            .O(N__32853),
            .I(N__32835));
    InMux I__8048 (
            .O(N__32852),
            .I(N__32835));
    CascadeMux I__8047 (
            .O(N__32851),
            .I(N__32831));
    InMux I__8046 (
            .O(N__32850),
            .I(N__32818));
    InMux I__8045 (
            .O(N__32849),
            .I(N__32815));
    InMux I__8044 (
            .O(N__32848),
            .I(N__32812));
    InMux I__8043 (
            .O(N__32847),
            .I(N__32805));
    InMux I__8042 (
            .O(N__32846),
            .I(N__32805));
    InMux I__8041 (
            .O(N__32845),
            .I(N__32805));
    InMux I__8040 (
            .O(N__32844),
            .I(N__32800));
    InMux I__8039 (
            .O(N__32843),
            .I(N__32800));
    LocalMux I__8038 (
            .O(N__32840),
            .I(N__32795));
    LocalMux I__8037 (
            .O(N__32835),
            .I(N__32795));
    InMux I__8036 (
            .O(N__32834),
            .I(N__32792));
    InMux I__8035 (
            .O(N__32831),
            .I(N__32781));
    InMux I__8034 (
            .O(N__32830),
            .I(N__32778));
    InMux I__8033 (
            .O(N__32829),
            .I(N__32765));
    InMux I__8032 (
            .O(N__32828),
            .I(N__32765));
    InMux I__8031 (
            .O(N__32827),
            .I(N__32762));
    InMux I__8030 (
            .O(N__32826),
            .I(N__32747));
    InMux I__8029 (
            .O(N__32825),
            .I(N__32743));
    InMux I__8028 (
            .O(N__32824),
            .I(N__32740));
    InMux I__8027 (
            .O(N__32823),
            .I(N__32735));
    InMux I__8026 (
            .O(N__32822),
            .I(N__32735));
    InMux I__8025 (
            .O(N__32821),
            .I(N__32732));
    LocalMux I__8024 (
            .O(N__32818),
            .I(N__32727));
    LocalMux I__8023 (
            .O(N__32815),
            .I(N__32727));
    LocalMux I__8022 (
            .O(N__32812),
            .I(N__32724));
    LocalMux I__8021 (
            .O(N__32805),
            .I(N__32716));
    LocalMux I__8020 (
            .O(N__32800),
            .I(N__32716));
    Span4Mux_h I__8019 (
            .O(N__32795),
            .I(N__32716));
    LocalMux I__8018 (
            .O(N__32792),
            .I(N__32713));
    InMux I__8017 (
            .O(N__32791),
            .I(N__32710));
    InMux I__8016 (
            .O(N__32790),
            .I(N__32707));
    InMux I__8015 (
            .O(N__32789),
            .I(N__32704));
    InMux I__8014 (
            .O(N__32788),
            .I(N__32699));
    InMux I__8013 (
            .O(N__32787),
            .I(N__32699));
    InMux I__8012 (
            .O(N__32786),
            .I(N__32696));
    InMux I__8011 (
            .O(N__32785),
            .I(N__32691));
    InMux I__8010 (
            .O(N__32784),
            .I(N__32691));
    LocalMux I__8009 (
            .O(N__32781),
            .I(N__32688));
    LocalMux I__8008 (
            .O(N__32778),
            .I(N__32685));
    InMux I__8007 (
            .O(N__32777),
            .I(N__32682));
    InMux I__8006 (
            .O(N__32776),
            .I(N__32675));
    InMux I__8005 (
            .O(N__32775),
            .I(N__32675));
    InMux I__8004 (
            .O(N__32774),
            .I(N__32675));
    InMux I__8003 (
            .O(N__32773),
            .I(N__32672));
    InMux I__8002 (
            .O(N__32772),
            .I(N__32669));
    InMux I__8001 (
            .O(N__32771),
            .I(N__32664));
    InMux I__8000 (
            .O(N__32770),
            .I(N__32664));
    LocalMux I__7999 (
            .O(N__32765),
            .I(N__32659));
    LocalMux I__7998 (
            .O(N__32762),
            .I(N__32659));
    InMux I__7997 (
            .O(N__32761),
            .I(N__32650));
    InMux I__7996 (
            .O(N__32760),
            .I(N__32650));
    InMux I__7995 (
            .O(N__32759),
            .I(N__32650));
    InMux I__7994 (
            .O(N__32758),
            .I(N__32650));
    InMux I__7993 (
            .O(N__32757),
            .I(N__32645));
    InMux I__7992 (
            .O(N__32756),
            .I(N__32645));
    InMux I__7991 (
            .O(N__32755),
            .I(N__32640));
    InMux I__7990 (
            .O(N__32754),
            .I(N__32640));
    InMux I__7989 (
            .O(N__32753),
            .I(N__32634));
    InMux I__7988 (
            .O(N__32752),
            .I(N__32629));
    InMux I__7987 (
            .O(N__32751),
            .I(N__32629));
    InMux I__7986 (
            .O(N__32750),
            .I(N__32626));
    LocalMux I__7985 (
            .O(N__32747),
            .I(N__32617));
    InMux I__7984 (
            .O(N__32746),
            .I(N__32613));
    LocalMux I__7983 (
            .O(N__32743),
            .I(N__32600));
    LocalMux I__7982 (
            .O(N__32740),
            .I(N__32600));
    LocalMux I__7981 (
            .O(N__32735),
            .I(N__32600));
    LocalMux I__7980 (
            .O(N__32732),
            .I(N__32600));
    Sp12to4 I__7979 (
            .O(N__32727),
            .I(N__32600));
    Sp12to4 I__7978 (
            .O(N__32724),
            .I(N__32600));
    InMux I__7977 (
            .O(N__32723),
            .I(N__32597));
    Span4Mux_v I__7976 (
            .O(N__32716),
            .I(N__32590));
    Span4Mux_h I__7975 (
            .O(N__32713),
            .I(N__32590));
    LocalMux I__7974 (
            .O(N__32710),
            .I(N__32590));
    LocalMux I__7973 (
            .O(N__32707),
            .I(N__32585));
    LocalMux I__7972 (
            .O(N__32704),
            .I(N__32582));
    LocalMux I__7971 (
            .O(N__32699),
            .I(N__32577));
    LocalMux I__7970 (
            .O(N__32696),
            .I(N__32577));
    LocalMux I__7969 (
            .O(N__32691),
            .I(N__32574));
    Span4Mux_v I__7968 (
            .O(N__32688),
            .I(N__32567));
    Span4Mux_v I__7967 (
            .O(N__32685),
            .I(N__32567));
    LocalMux I__7966 (
            .O(N__32682),
            .I(N__32567));
    LocalMux I__7965 (
            .O(N__32675),
            .I(N__32564));
    LocalMux I__7964 (
            .O(N__32672),
            .I(N__32561));
    LocalMux I__7963 (
            .O(N__32669),
            .I(N__32548));
    LocalMux I__7962 (
            .O(N__32664),
            .I(N__32548));
    Span4Mux_h I__7961 (
            .O(N__32659),
            .I(N__32548));
    LocalMux I__7960 (
            .O(N__32650),
            .I(N__32548));
    LocalMux I__7959 (
            .O(N__32645),
            .I(N__32548));
    LocalMux I__7958 (
            .O(N__32640),
            .I(N__32548));
    InMux I__7957 (
            .O(N__32639),
            .I(N__32545));
    InMux I__7956 (
            .O(N__32638),
            .I(N__32542));
    InMux I__7955 (
            .O(N__32637),
            .I(N__32539));
    LocalMux I__7954 (
            .O(N__32634),
            .I(N__32532));
    LocalMux I__7953 (
            .O(N__32629),
            .I(N__32532));
    LocalMux I__7952 (
            .O(N__32626),
            .I(N__32532));
    InMux I__7951 (
            .O(N__32625),
            .I(N__32529));
    InMux I__7950 (
            .O(N__32624),
            .I(N__32526));
    InMux I__7949 (
            .O(N__32623),
            .I(N__32523));
    InMux I__7948 (
            .O(N__32622),
            .I(N__32518));
    InMux I__7947 (
            .O(N__32621),
            .I(N__32518));
    InMux I__7946 (
            .O(N__32620),
            .I(N__32515));
    Span12Mux_h I__7945 (
            .O(N__32617),
            .I(N__32512));
    InMux I__7944 (
            .O(N__32616),
            .I(N__32509));
    LocalMux I__7943 (
            .O(N__32613),
            .I(N__32502));
    Span12Mux_v I__7942 (
            .O(N__32600),
            .I(N__32502));
    LocalMux I__7941 (
            .O(N__32597),
            .I(N__32502));
    Span4Mux_v I__7940 (
            .O(N__32590),
            .I(N__32499));
    InMux I__7939 (
            .O(N__32589),
            .I(N__32494));
    InMux I__7938 (
            .O(N__32588),
            .I(N__32494));
    Span4Mux_h I__7937 (
            .O(N__32585),
            .I(N__32487));
    Span4Mux_h I__7936 (
            .O(N__32582),
            .I(N__32487));
    Span4Mux_h I__7935 (
            .O(N__32577),
            .I(N__32487));
    Span4Mux_h I__7934 (
            .O(N__32574),
            .I(N__32476));
    Span4Mux_h I__7933 (
            .O(N__32567),
            .I(N__32476));
    Span4Mux_h I__7932 (
            .O(N__32564),
            .I(N__32476));
    Span4Mux_h I__7931 (
            .O(N__32561),
            .I(N__32476));
    Span4Mux_v I__7930 (
            .O(N__32548),
            .I(N__32476));
    LocalMux I__7929 (
            .O(N__32545),
            .I(N__32471));
    LocalMux I__7928 (
            .O(N__32542),
            .I(N__32471));
    LocalMux I__7927 (
            .O(N__32539),
            .I(N__32464));
    Span4Mux_v I__7926 (
            .O(N__32532),
            .I(N__32464));
    LocalMux I__7925 (
            .O(N__32529),
            .I(N__32464));
    LocalMux I__7924 (
            .O(N__32526),
            .I(N_389_0));
    LocalMux I__7923 (
            .O(N__32523),
            .I(N_389_0));
    LocalMux I__7922 (
            .O(N__32518),
            .I(N_389_0));
    LocalMux I__7921 (
            .O(N__32515),
            .I(N_389_0));
    Odrv12 I__7920 (
            .O(N__32512),
            .I(N_389_0));
    LocalMux I__7919 (
            .O(N__32509),
            .I(N_389_0));
    Odrv12 I__7918 (
            .O(N__32502),
            .I(N_389_0));
    Odrv4 I__7917 (
            .O(N__32499),
            .I(N_389_0));
    LocalMux I__7916 (
            .O(N__32494),
            .I(N_389_0));
    Odrv4 I__7915 (
            .O(N__32487),
            .I(N_389_0));
    Odrv4 I__7914 (
            .O(N__32476),
            .I(N_389_0));
    Odrv12 I__7913 (
            .O(N__32471),
            .I(N_389_0));
    Odrv4 I__7912 (
            .O(N__32464),
            .I(N_389_0));
    InMux I__7911 (
            .O(N__32437),
            .I(N__32424));
    InMux I__7910 (
            .O(N__32436),
            .I(N__32421));
    InMux I__7909 (
            .O(N__32435),
            .I(N__32418));
    InMux I__7908 (
            .O(N__32434),
            .I(N__32415));
    InMux I__7907 (
            .O(N__32433),
            .I(N__32412));
    InMux I__7906 (
            .O(N__32432),
            .I(N__32409));
    InMux I__7905 (
            .O(N__32431),
            .I(N__32406));
    InMux I__7904 (
            .O(N__32430),
            .I(N__32403));
    InMux I__7903 (
            .O(N__32429),
            .I(N__32400));
    InMux I__7902 (
            .O(N__32428),
            .I(N__32397));
    InMux I__7901 (
            .O(N__32427),
            .I(N__32394));
    LocalMux I__7900 (
            .O(N__32424),
            .I(N__32370));
    LocalMux I__7899 (
            .O(N__32421),
            .I(N__32367));
    LocalMux I__7898 (
            .O(N__32418),
            .I(N__32364));
    LocalMux I__7897 (
            .O(N__32415),
            .I(N__32361));
    LocalMux I__7896 (
            .O(N__32412),
            .I(N__32358));
    LocalMux I__7895 (
            .O(N__32409),
            .I(N__32355));
    LocalMux I__7894 (
            .O(N__32406),
            .I(N__32352));
    LocalMux I__7893 (
            .O(N__32403),
            .I(N__32349));
    LocalMux I__7892 (
            .O(N__32400),
            .I(N__32346));
    LocalMux I__7891 (
            .O(N__32397),
            .I(N__32343));
    LocalMux I__7890 (
            .O(N__32394),
            .I(N__32340));
    SRMux I__7889 (
            .O(N__32393),
            .I(N__32275));
    SRMux I__7888 (
            .O(N__32392),
            .I(N__32275));
    SRMux I__7887 (
            .O(N__32391),
            .I(N__32275));
    SRMux I__7886 (
            .O(N__32390),
            .I(N__32275));
    SRMux I__7885 (
            .O(N__32389),
            .I(N__32275));
    SRMux I__7884 (
            .O(N__32388),
            .I(N__32275));
    SRMux I__7883 (
            .O(N__32387),
            .I(N__32275));
    SRMux I__7882 (
            .O(N__32386),
            .I(N__32275));
    SRMux I__7881 (
            .O(N__32385),
            .I(N__32275));
    SRMux I__7880 (
            .O(N__32384),
            .I(N__32275));
    SRMux I__7879 (
            .O(N__32383),
            .I(N__32275));
    SRMux I__7878 (
            .O(N__32382),
            .I(N__32275));
    SRMux I__7877 (
            .O(N__32381),
            .I(N__32275));
    SRMux I__7876 (
            .O(N__32380),
            .I(N__32275));
    SRMux I__7875 (
            .O(N__32379),
            .I(N__32275));
    SRMux I__7874 (
            .O(N__32378),
            .I(N__32275));
    SRMux I__7873 (
            .O(N__32377),
            .I(N__32275));
    SRMux I__7872 (
            .O(N__32376),
            .I(N__32275));
    SRMux I__7871 (
            .O(N__32375),
            .I(N__32275));
    SRMux I__7870 (
            .O(N__32374),
            .I(N__32275));
    SRMux I__7869 (
            .O(N__32373),
            .I(N__32275));
    Glb2LocalMux I__7868 (
            .O(N__32370),
            .I(N__32275));
    Glb2LocalMux I__7867 (
            .O(N__32367),
            .I(N__32275));
    Glb2LocalMux I__7866 (
            .O(N__32364),
            .I(N__32275));
    Glb2LocalMux I__7865 (
            .O(N__32361),
            .I(N__32275));
    Glb2LocalMux I__7864 (
            .O(N__32358),
            .I(N__32275));
    Glb2LocalMux I__7863 (
            .O(N__32355),
            .I(N__32275));
    Glb2LocalMux I__7862 (
            .O(N__32352),
            .I(N__32275));
    Glb2LocalMux I__7861 (
            .O(N__32349),
            .I(N__32275));
    Glb2LocalMux I__7860 (
            .O(N__32346),
            .I(N__32275));
    Glb2LocalMux I__7859 (
            .O(N__32343),
            .I(N__32275));
    Glb2LocalMux I__7858 (
            .O(N__32340),
            .I(N__32275));
    GlobalMux I__7857 (
            .O(N__32275),
            .I(N__32272));
    gio2CtrlBuf I__7856 (
            .O(N__32272),
            .I(M_this_reset_cond_out_g_0));
    CascadeMux I__7855 (
            .O(N__32269),
            .I(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8_cascade_ ));
    InMux I__7854 (
            .O(N__32266),
            .I(N__32263));
    LocalMux I__7853 (
            .O(N__32263),
            .I(N__32260));
    Odrv4 I__7852 (
            .O(N__32260),
            .I(\this_vga_signals.M_this_data_count_q_3_bmZ0Z_13 ));
    CascadeMux I__7851 (
            .O(N__32257),
            .I(\this_vga_signals.M_this_data_count_q_3_amZ0Z_13_cascade_ ));
    InMux I__7850 (
            .O(N__32254),
            .I(N__32242));
    InMux I__7849 (
            .O(N__32253),
            .I(N__32242));
    InMux I__7848 (
            .O(N__32252),
            .I(N__32242));
    InMux I__7847 (
            .O(N__32251),
            .I(N__32227));
    InMux I__7846 (
            .O(N__32250),
            .I(N__32227));
    InMux I__7845 (
            .O(N__32249),
            .I(N__32227));
    LocalMux I__7844 (
            .O(N__32242),
            .I(N__32224));
    InMux I__7843 (
            .O(N__32241),
            .I(N__32219));
    InMux I__7842 (
            .O(N__32240),
            .I(N__32219));
    InMux I__7841 (
            .O(N__32239),
            .I(N__32214));
    InMux I__7840 (
            .O(N__32238),
            .I(N__32214));
    InMux I__7839 (
            .O(N__32237),
            .I(N__32205));
    InMux I__7838 (
            .O(N__32236),
            .I(N__32205));
    InMux I__7837 (
            .O(N__32235),
            .I(N__32205));
    InMux I__7836 (
            .O(N__32234),
            .I(N__32205));
    LocalMux I__7835 (
            .O(N__32227),
            .I(N__32200));
    Sp12to4 I__7834 (
            .O(N__32224),
            .I(N__32193));
    LocalMux I__7833 (
            .O(N__32219),
            .I(N__32193));
    LocalMux I__7832 (
            .O(N__32214),
            .I(N__32193));
    LocalMux I__7831 (
            .O(N__32205),
            .I(N__32190));
    InMux I__7830 (
            .O(N__32204),
            .I(N__32185));
    InMux I__7829 (
            .O(N__32203),
            .I(N__32185));
    Odrv4 I__7828 (
            .O(N__32200),
            .I(M_this_data_count_q_3_sn_N_2));
    Odrv12 I__7827 (
            .O(N__32193),
            .I(M_this_data_count_q_3_sn_N_2));
    Odrv4 I__7826 (
            .O(N__32190),
            .I(M_this_data_count_q_3_sn_N_2));
    LocalMux I__7825 (
            .O(N__32185),
            .I(M_this_data_count_q_3_sn_N_2));
    InMux I__7824 (
            .O(N__32176),
            .I(N__32173));
    LocalMux I__7823 (
            .O(N__32173),
            .I(M_this_data_count_q_cry_12_THRU_CO));
    CascadeMux I__7822 (
            .O(N__32170),
            .I(M_this_data_count_q_3_13_cascade_));
    InMux I__7821 (
            .O(N__32167),
            .I(N__32147));
    InMux I__7820 (
            .O(N__32166),
            .I(N__32147));
    InMux I__7819 (
            .O(N__32165),
            .I(N__32147));
    InMux I__7818 (
            .O(N__32164),
            .I(N__32138));
    InMux I__7817 (
            .O(N__32163),
            .I(N__32138));
    InMux I__7816 (
            .O(N__32162),
            .I(N__32138));
    InMux I__7815 (
            .O(N__32161),
            .I(N__32138));
    InMux I__7814 (
            .O(N__32160),
            .I(N__32127));
    InMux I__7813 (
            .O(N__32159),
            .I(N__32127));
    InMux I__7812 (
            .O(N__32158),
            .I(N__32127));
    InMux I__7811 (
            .O(N__32157),
            .I(N__32127));
    InMux I__7810 (
            .O(N__32156),
            .I(N__32120));
    InMux I__7809 (
            .O(N__32155),
            .I(N__32120));
    InMux I__7808 (
            .O(N__32154),
            .I(N__32120));
    LocalMux I__7807 (
            .O(N__32147),
            .I(N__32115));
    LocalMux I__7806 (
            .O(N__32138),
            .I(N__32115));
    InMux I__7805 (
            .O(N__32137),
            .I(N__32110));
    InMux I__7804 (
            .O(N__32136),
            .I(N__32110));
    LocalMux I__7803 (
            .O(N__32127),
            .I(N__32107));
    LocalMux I__7802 (
            .O(N__32120),
            .I(N__32104));
    Span4Mux_v I__7801 (
            .O(N__32115),
            .I(N__32099));
    LocalMux I__7800 (
            .O(N__32110),
            .I(N__32099));
    Odrv4 I__7799 (
            .O(N__32107),
            .I(N_570_0_i));
    Odrv4 I__7798 (
            .O(N__32104),
            .I(N_570_0_i));
    Odrv4 I__7797 (
            .O(N__32099),
            .I(N_570_0_i));
    InMux I__7796 (
            .O(N__32092),
            .I(N__32089));
    LocalMux I__7795 (
            .O(N__32089),
            .I(N__32083));
    InMux I__7794 (
            .O(N__32088),
            .I(N__32080));
    InMux I__7793 (
            .O(N__32087),
            .I(N__32077));
    InMux I__7792 (
            .O(N__32086),
            .I(N__32074));
    Span4Mux_h I__7791 (
            .O(N__32083),
            .I(N__32071));
    LocalMux I__7790 (
            .O(N__32080),
            .I(M_this_data_count_qZ0Z_13));
    LocalMux I__7789 (
            .O(N__32077),
            .I(M_this_data_count_qZ0Z_13));
    LocalMux I__7788 (
            .O(N__32074),
            .I(M_this_data_count_qZ0Z_13));
    Odrv4 I__7787 (
            .O(N__32071),
            .I(M_this_data_count_qZ0Z_13));
    ClkMux I__7786 (
            .O(N__32062),
            .I(N__31684));
    ClkMux I__7785 (
            .O(N__32061),
            .I(N__31684));
    ClkMux I__7784 (
            .O(N__32060),
            .I(N__31684));
    ClkMux I__7783 (
            .O(N__32059),
            .I(N__31684));
    ClkMux I__7782 (
            .O(N__32058),
            .I(N__31684));
    ClkMux I__7781 (
            .O(N__32057),
            .I(N__31684));
    ClkMux I__7780 (
            .O(N__32056),
            .I(N__31684));
    ClkMux I__7779 (
            .O(N__32055),
            .I(N__31684));
    ClkMux I__7778 (
            .O(N__32054),
            .I(N__31684));
    ClkMux I__7777 (
            .O(N__32053),
            .I(N__31684));
    ClkMux I__7776 (
            .O(N__32052),
            .I(N__31684));
    ClkMux I__7775 (
            .O(N__32051),
            .I(N__31684));
    ClkMux I__7774 (
            .O(N__32050),
            .I(N__31684));
    ClkMux I__7773 (
            .O(N__32049),
            .I(N__31684));
    ClkMux I__7772 (
            .O(N__32048),
            .I(N__31684));
    ClkMux I__7771 (
            .O(N__32047),
            .I(N__31684));
    ClkMux I__7770 (
            .O(N__32046),
            .I(N__31684));
    ClkMux I__7769 (
            .O(N__32045),
            .I(N__31684));
    ClkMux I__7768 (
            .O(N__32044),
            .I(N__31684));
    ClkMux I__7767 (
            .O(N__32043),
            .I(N__31684));
    ClkMux I__7766 (
            .O(N__32042),
            .I(N__31684));
    ClkMux I__7765 (
            .O(N__32041),
            .I(N__31684));
    ClkMux I__7764 (
            .O(N__32040),
            .I(N__31684));
    ClkMux I__7763 (
            .O(N__32039),
            .I(N__31684));
    ClkMux I__7762 (
            .O(N__32038),
            .I(N__31684));
    ClkMux I__7761 (
            .O(N__32037),
            .I(N__31684));
    ClkMux I__7760 (
            .O(N__32036),
            .I(N__31684));
    ClkMux I__7759 (
            .O(N__32035),
            .I(N__31684));
    ClkMux I__7758 (
            .O(N__32034),
            .I(N__31684));
    ClkMux I__7757 (
            .O(N__32033),
            .I(N__31684));
    ClkMux I__7756 (
            .O(N__32032),
            .I(N__31684));
    ClkMux I__7755 (
            .O(N__32031),
            .I(N__31684));
    ClkMux I__7754 (
            .O(N__32030),
            .I(N__31684));
    ClkMux I__7753 (
            .O(N__32029),
            .I(N__31684));
    ClkMux I__7752 (
            .O(N__32028),
            .I(N__31684));
    ClkMux I__7751 (
            .O(N__32027),
            .I(N__31684));
    ClkMux I__7750 (
            .O(N__32026),
            .I(N__31684));
    ClkMux I__7749 (
            .O(N__32025),
            .I(N__31684));
    ClkMux I__7748 (
            .O(N__32024),
            .I(N__31684));
    ClkMux I__7747 (
            .O(N__32023),
            .I(N__31684));
    ClkMux I__7746 (
            .O(N__32022),
            .I(N__31684));
    ClkMux I__7745 (
            .O(N__32021),
            .I(N__31684));
    ClkMux I__7744 (
            .O(N__32020),
            .I(N__31684));
    ClkMux I__7743 (
            .O(N__32019),
            .I(N__31684));
    ClkMux I__7742 (
            .O(N__32018),
            .I(N__31684));
    ClkMux I__7741 (
            .O(N__32017),
            .I(N__31684));
    ClkMux I__7740 (
            .O(N__32016),
            .I(N__31684));
    ClkMux I__7739 (
            .O(N__32015),
            .I(N__31684));
    ClkMux I__7738 (
            .O(N__32014),
            .I(N__31684));
    ClkMux I__7737 (
            .O(N__32013),
            .I(N__31684));
    ClkMux I__7736 (
            .O(N__32012),
            .I(N__31684));
    ClkMux I__7735 (
            .O(N__32011),
            .I(N__31684));
    ClkMux I__7734 (
            .O(N__32010),
            .I(N__31684));
    ClkMux I__7733 (
            .O(N__32009),
            .I(N__31684));
    ClkMux I__7732 (
            .O(N__32008),
            .I(N__31684));
    ClkMux I__7731 (
            .O(N__32007),
            .I(N__31684));
    ClkMux I__7730 (
            .O(N__32006),
            .I(N__31684));
    ClkMux I__7729 (
            .O(N__32005),
            .I(N__31684));
    ClkMux I__7728 (
            .O(N__32004),
            .I(N__31684));
    ClkMux I__7727 (
            .O(N__32003),
            .I(N__31684));
    ClkMux I__7726 (
            .O(N__32002),
            .I(N__31684));
    ClkMux I__7725 (
            .O(N__32001),
            .I(N__31684));
    ClkMux I__7724 (
            .O(N__32000),
            .I(N__31684));
    ClkMux I__7723 (
            .O(N__31999),
            .I(N__31684));
    ClkMux I__7722 (
            .O(N__31998),
            .I(N__31684));
    ClkMux I__7721 (
            .O(N__31997),
            .I(N__31684));
    ClkMux I__7720 (
            .O(N__31996),
            .I(N__31684));
    ClkMux I__7719 (
            .O(N__31995),
            .I(N__31684));
    ClkMux I__7718 (
            .O(N__31994),
            .I(N__31684));
    ClkMux I__7717 (
            .O(N__31993),
            .I(N__31684));
    ClkMux I__7716 (
            .O(N__31992),
            .I(N__31684));
    ClkMux I__7715 (
            .O(N__31991),
            .I(N__31684));
    ClkMux I__7714 (
            .O(N__31990),
            .I(N__31684));
    ClkMux I__7713 (
            .O(N__31989),
            .I(N__31684));
    ClkMux I__7712 (
            .O(N__31988),
            .I(N__31684));
    ClkMux I__7711 (
            .O(N__31987),
            .I(N__31684));
    ClkMux I__7710 (
            .O(N__31986),
            .I(N__31684));
    ClkMux I__7709 (
            .O(N__31985),
            .I(N__31684));
    ClkMux I__7708 (
            .O(N__31984),
            .I(N__31684));
    ClkMux I__7707 (
            .O(N__31983),
            .I(N__31684));
    ClkMux I__7706 (
            .O(N__31982),
            .I(N__31684));
    ClkMux I__7705 (
            .O(N__31981),
            .I(N__31684));
    ClkMux I__7704 (
            .O(N__31980),
            .I(N__31684));
    ClkMux I__7703 (
            .O(N__31979),
            .I(N__31684));
    ClkMux I__7702 (
            .O(N__31978),
            .I(N__31684));
    ClkMux I__7701 (
            .O(N__31977),
            .I(N__31684));
    ClkMux I__7700 (
            .O(N__31976),
            .I(N__31684));
    ClkMux I__7699 (
            .O(N__31975),
            .I(N__31684));
    ClkMux I__7698 (
            .O(N__31974),
            .I(N__31684));
    ClkMux I__7697 (
            .O(N__31973),
            .I(N__31684));
    ClkMux I__7696 (
            .O(N__31972),
            .I(N__31684));
    ClkMux I__7695 (
            .O(N__31971),
            .I(N__31684));
    ClkMux I__7694 (
            .O(N__31970),
            .I(N__31684));
    ClkMux I__7693 (
            .O(N__31969),
            .I(N__31684));
    ClkMux I__7692 (
            .O(N__31968),
            .I(N__31684));
    ClkMux I__7691 (
            .O(N__31967),
            .I(N__31684));
    ClkMux I__7690 (
            .O(N__31966),
            .I(N__31684));
    ClkMux I__7689 (
            .O(N__31965),
            .I(N__31684));
    ClkMux I__7688 (
            .O(N__31964),
            .I(N__31684));
    ClkMux I__7687 (
            .O(N__31963),
            .I(N__31684));
    ClkMux I__7686 (
            .O(N__31962),
            .I(N__31684));
    ClkMux I__7685 (
            .O(N__31961),
            .I(N__31684));
    ClkMux I__7684 (
            .O(N__31960),
            .I(N__31684));
    ClkMux I__7683 (
            .O(N__31959),
            .I(N__31684));
    ClkMux I__7682 (
            .O(N__31958),
            .I(N__31684));
    ClkMux I__7681 (
            .O(N__31957),
            .I(N__31684));
    ClkMux I__7680 (
            .O(N__31956),
            .I(N__31684));
    ClkMux I__7679 (
            .O(N__31955),
            .I(N__31684));
    ClkMux I__7678 (
            .O(N__31954),
            .I(N__31684));
    ClkMux I__7677 (
            .O(N__31953),
            .I(N__31684));
    ClkMux I__7676 (
            .O(N__31952),
            .I(N__31684));
    ClkMux I__7675 (
            .O(N__31951),
            .I(N__31684));
    ClkMux I__7674 (
            .O(N__31950),
            .I(N__31684));
    ClkMux I__7673 (
            .O(N__31949),
            .I(N__31684));
    ClkMux I__7672 (
            .O(N__31948),
            .I(N__31684));
    ClkMux I__7671 (
            .O(N__31947),
            .I(N__31684));
    ClkMux I__7670 (
            .O(N__31946),
            .I(N__31684));
    ClkMux I__7669 (
            .O(N__31945),
            .I(N__31684));
    ClkMux I__7668 (
            .O(N__31944),
            .I(N__31684));
    ClkMux I__7667 (
            .O(N__31943),
            .I(N__31684));
    ClkMux I__7666 (
            .O(N__31942),
            .I(N__31684));
    ClkMux I__7665 (
            .O(N__31941),
            .I(N__31684));
    ClkMux I__7664 (
            .O(N__31940),
            .I(N__31684));
    ClkMux I__7663 (
            .O(N__31939),
            .I(N__31684));
    ClkMux I__7662 (
            .O(N__31938),
            .I(N__31684));
    ClkMux I__7661 (
            .O(N__31937),
            .I(N__31684));
    GlobalMux I__7660 (
            .O(N__31684),
            .I(N__31681));
    gio2CtrlBuf I__7659 (
            .O(N__31681),
            .I(clk_0_c_g));
    CEMux I__7658 (
            .O(N__31678),
            .I(N__31673));
    CEMux I__7657 (
            .O(N__31677),
            .I(N__31670));
    CEMux I__7656 (
            .O(N__31676),
            .I(N__31665));
    LocalMux I__7655 (
            .O(N__31673),
            .I(N__31660));
    LocalMux I__7654 (
            .O(N__31670),
            .I(N__31660));
    CEMux I__7653 (
            .O(N__31669),
            .I(N__31657));
    CEMux I__7652 (
            .O(N__31668),
            .I(N__31654));
    LocalMux I__7651 (
            .O(N__31665),
            .I(N__31651));
    Span4Mux_v I__7650 (
            .O(N__31660),
            .I(N__31648));
    LocalMux I__7649 (
            .O(N__31657),
            .I(N__31643));
    LocalMux I__7648 (
            .O(N__31654),
            .I(N__31643));
    Odrv4 I__7647 (
            .O(N__31651),
            .I(M_this_data_count_qe_0_i));
    Odrv4 I__7646 (
            .O(N__31648),
            .I(M_this_data_count_qe_0_i));
    Odrv4 I__7645 (
            .O(N__31643),
            .I(M_this_data_count_qe_0_i));
    InMux I__7644 (
            .O(N__31636),
            .I(N__31631));
    InMux I__7643 (
            .O(N__31635),
            .I(N__31628));
    InMux I__7642 (
            .O(N__31634),
            .I(N__31625));
    LocalMux I__7641 (
            .O(N__31631),
            .I(N__31622));
    LocalMux I__7640 (
            .O(N__31628),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__7639 (
            .O(N__31625),
            .I(M_this_data_count_qZ0Z_9));
    Odrv4 I__7638 (
            .O(N__31622),
            .I(M_this_data_count_qZ0Z_9));
    CascadeMux I__7637 (
            .O(N__31615),
            .I(N__31612));
    InMux I__7636 (
            .O(N__31612),
            .I(N__31607));
    InMux I__7635 (
            .O(N__31611),
            .I(N__31604));
    InMux I__7634 (
            .O(N__31610),
            .I(N__31601));
    LocalMux I__7633 (
            .O(N__31607),
            .I(N__31598));
    LocalMux I__7632 (
            .O(N__31604),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__7631 (
            .O(N__31601),
            .I(M_this_data_count_qZ0Z_11));
    Odrv4 I__7630 (
            .O(N__31598),
            .I(M_this_data_count_qZ0Z_11));
    CascadeMux I__7629 (
            .O(N__31591),
            .I(N__31586));
    InMux I__7628 (
            .O(N__31590),
            .I(N__31583));
    InMux I__7627 (
            .O(N__31589),
            .I(N__31580));
    InMux I__7626 (
            .O(N__31586),
            .I(N__31577));
    LocalMux I__7625 (
            .O(N__31583),
            .I(N__31574));
    LocalMux I__7624 (
            .O(N__31580),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__7623 (
            .O(N__31577),
            .I(M_this_data_count_qZ0Z_8));
    Odrv4 I__7622 (
            .O(N__31574),
            .I(M_this_data_count_qZ0Z_8));
    InMux I__7621 (
            .O(N__31567),
            .I(N__31563));
    InMux I__7620 (
            .O(N__31566),
            .I(N__31560));
    LocalMux I__7619 (
            .O(N__31563),
            .I(N__31557));
    LocalMux I__7618 (
            .O(N__31560),
            .I(N__31552));
    Span4Mux_v I__7617 (
            .O(N__31557),
            .I(N__31552));
    Span4Mux_v I__7616 (
            .O(N__31552),
            .I(N__31549));
    Odrv4 I__7615 (
            .O(N__31549),
            .I(M_this_state_d88_10));
    CascadeMux I__7614 (
            .O(N__31546),
            .I(N__31541));
    InMux I__7613 (
            .O(N__31545),
            .I(N__31538));
    InMux I__7612 (
            .O(N__31544),
            .I(N__31534));
    InMux I__7611 (
            .O(N__31541),
            .I(N__31531));
    LocalMux I__7610 (
            .O(N__31538),
            .I(N__31528));
    InMux I__7609 (
            .O(N__31537),
            .I(N__31525));
    LocalMux I__7608 (
            .O(N__31534),
            .I(M_this_data_count_qZ0Z_10));
    LocalMux I__7607 (
            .O(N__31531),
            .I(M_this_data_count_qZ0Z_10));
    Odrv4 I__7606 (
            .O(N__31528),
            .I(M_this_data_count_qZ0Z_10));
    LocalMux I__7605 (
            .O(N__31525),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__7604 (
            .O(N__31516),
            .I(N__31509));
    InMux I__7603 (
            .O(N__31515),
            .I(N__31509));
    InMux I__7602 (
            .O(N__31514),
            .I(N__31502));
    LocalMux I__7601 (
            .O(N__31509),
            .I(N__31499));
    InMux I__7600 (
            .O(N__31508),
            .I(N__31490));
    InMux I__7599 (
            .O(N__31507),
            .I(N__31490));
    InMux I__7598 (
            .O(N__31506),
            .I(N__31490));
    InMux I__7597 (
            .O(N__31505),
            .I(N__31490));
    LocalMux I__7596 (
            .O(N__31502),
            .I(N__31487));
    Odrv4 I__7595 (
            .O(N__31499),
            .I(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8 ));
    LocalMux I__7594 (
            .O(N__31490),
            .I(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8 ));
    Odrv4 I__7593 (
            .O(N__31487),
            .I(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8 ));
    InMux I__7592 (
            .O(N__31480),
            .I(N__31477));
    LocalMux I__7591 (
            .O(N__31477),
            .I(N__31474));
    Odrv4 I__7590 (
            .O(N__31474),
            .I(\this_vga_signals.M_this_data_count_q_3_amZ0Z_10 ));
    InMux I__7589 (
            .O(N__31471),
            .I(N__31468));
    LocalMux I__7588 (
            .O(N__31468),
            .I(N__31465));
    Span4Mux_s2_v I__7587 (
            .O(N__31465),
            .I(N__31462));
    Span4Mux_v I__7586 (
            .O(N__31462),
            .I(N__31459));
    Odrv4 I__7585 (
            .O(N__31459),
            .I(M_this_map_ram_write_data_6));
    CascadeMux I__7584 (
            .O(N__31456),
            .I(N__31453));
    InMux I__7583 (
            .O(N__31453),
            .I(N__31450));
    LocalMux I__7582 (
            .O(N__31450),
            .I(M_this_data_count_q_s_11));
    InMux I__7581 (
            .O(N__31447),
            .I(N__31444));
    LocalMux I__7580 (
            .O(N__31444),
            .I(M_this_data_count_q_s_12));
    CascadeMux I__7579 (
            .O(N__31441),
            .I(N_518_cascade_));
    CascadeMux I__7578 (
            .O(N__31438),
            .I(N__31433));
    InMux I__7577 (
            .O(N__31437),
            .I(N__31430));
    InMux I__7576 (
            .O(N__31436),
            .I(N__31427));
    InMux I__7575 (
            .O(N__31433),
            .I(N__31424));
    LocalMux I__7574 (
            .O(N__31430),
            .I(N__31421));
    LocalMux I__7573 (
            .O(N__31427),
            .I(M_this_data_count_qZ0Z_12));
    LocalMux I__7572 (
            .O(N__31424),
            .I(M_this_data_count_qZ0Z_12));
    Odrv4 I__7571 (
            .O(N__31421),
            .I(M_this_data_count_qZ0Z_12));
    InMux I__7570 (
            .O(N__31414),
            .I(N__31411));
    LocalMux I__7569 (
            .O(N__31411),
            .I(M_this_data_count_q_s_14));
    CascadeMux I__7568 (
            .O(N__31408),
            .I(N_520_cascade_));
    CascadeMux I__7567 (
            .O(N__31405),
            .I(N__31400));
    InMux I__7566 (
            .O(N__31404),
            .I(N__31397));
    InMux I__7565 (
            .O(N__31403),
            .I(N__31394));
    InMux I__7564 (
            .O(N__31400),
            .I(N__31391));
    LocalMux I__7563 (
            .O(N__31397),
            .I(N__31388));
    LocalMux I__7562 (
            .O(N__31394),
            .I(M_this_data_count_qZ0Z_14));
    LocalMux I__7561 (
            .O(N__31391),
            .I(M_this_data_count_qZ0Z_14));
    Odrv4 I__7560 (
            .O(N__31388),
            .I(M_this_data_count_qZ0Z_14));
    InMux I__7559 (
            .O(N__31381),
            .I(N__31378));
    LocalMux I__7558 (
            .O(N__31378),
            .I(M_this_data_count_q_s_15));
    CascadeMux I__7557 (
            .O(N__31375),
            .I(N_521_cascade_));
    CascadeMux I__7556 (
            .O(N__31372),
            .I(N__31369));
    InMux I__7555 (
            .O(N__31369),
            .I(N__31364));
    InMux I__7554 (
            .O(N__31368),
            .I(N__31361));
    InMux I__7553 (
            .O(N__31367),
            .I(N__31358));
    LocalMux I__7552 (
            .O(N__31364),
            .I(N__31355));
    LocalMux I__7551 (
            .O(N__31361),
            .I(M_this_data_count_qZ0Z_15));
    LocalMux I__7550 (
            .O(N__31358),
            .I(M_this_data_count_qZ0Z_15));
    Odrv4 I__7549 (
            .O(N__31355),
            .I(M_this_data_count_qZ0Z_15));
    InMux I__7548 (
            .O(N__31348),
            .I(N__31345));
    LocalMux I__7547 (
            .O(N__31345),
            .I(N_517));
    InMux I__7546 (
            .O(N__31342),
            .I(N__31339));
    LocalMux I__7545 (
            .O(N__31339),
            .I(N__31336));
    Span4Mux_v I__7544 (
            .O(N__31336),
            .I(N__31333));
    Span4Mux_h I__7543 (
            .O(N__31333),
            .I(N__31330));
    Odrv4 I__7542 (
            .O(N__31330),
            .I(\this_vga_signals.M_this_data_count_q_3_bmZ0Z_10 ));
    CascadeMux I__7541 (
            .O(N__31327),
            .I(N__31324));
    InMux I__7540 (
            .O(N__31324),
            .I(N__31320));
    CascadeMux I__7539 (
            .O(N__31323),
            .I(N__31313));
    LocalMux I__7538 (
            .O(N__31320),
            .I(N__31310));
    InMux I__7537 (
            .O(N__31319),
            .I(N__31307));
    InMux I__7536 (
            .O(N__31318),
            .I(N__31304));
    InMux I__7535 (
            .O(N__31317),
            .I(N__31301));
    InMux I__7534 (
            .O(N__31316),
            .I(N__31296));
    InMux I__7533 (
            .O(N__31313),
            .I(N__31296));
    Span4Mux_v I__7532 (
            .O(N__31310),
            .I(N__31290));
    LocalMux I__7531 (
            .O(N__31307),
            .I(N__31290));
    LocalMux I__7530 (
            .O(N__31304),
            .I(N__31287));
    LocalMux I__7529 (
            .O(N__31301),
            .I(N__31284));
    LocalMux I__7528 (
            .O(N__31296),
            .I(N__31281));
    InMux I__7527 (
            .O(N__31295),
            .I(N__31278));
    Span4Mux_h I__7526 (
            .O(N__31290),
            .I(N__31275));
    Span4Mux_h I__7525 (
            .O(N__31287),
            .I(N__31272));
    Span4Mux_h I__7524 (
            .O(N__31284),
            .I(N__31267));
    Span4Mux_h I__7523 (
            .O(N__31281),
            .I(N__31267));
    LocalMux I__7522 (
            .O(N__31278),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__7521 (
            .O(N__31275),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__7520 (
            .O(N__31272),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__7519 (
            .O(N__31267),
            .I(M_this_state_qZ0Z_13));
    CascadeMux I__7518 (
            .O(N__31258),
            .I(N__31255));
    InMux I__7517 (
            .O(N__31255),
            .I(N__31249));
    InMux I__7516 (
            .O(N__31254),
            .I(N__31246));
    InMux I__7515 (
            .O(N__31253),
            .I(N__31243));
    InMux I__7514 (
            .O(N__31252),
            .I(N__31240));
    LocalMux I__7513 (
            .O(N__31249),
            .I(N__31237));
    LocalMux I__7512 (
            .O(N__31246),
            .I(N__31232));
    LocalMux I__7511 (
            .O(N__31243),
            .I(N__31232));
    LocalMux I__7510 (
            .O(N__31240),
            .I(N__31228));
    Span4Mux_h I__7509 (
            .O(N__31237),
            .I(N__31223));
    Span4Mux_v I__7508 (
            .O(N__31232),
            .I(N__31223));
    InMux I__7507 (
            .O(N__31231),
            .I(N__31220));
    Span12Mux_h I__7506 (
            .O(N__31228),
            .I(N__31217));
    Odrv4 I__7505 (
            .O(N__31223),
            .I(N_391_0));
    LocalMux I__7504 (
            .O(N__31220),
            .I(N_391_0));
    Odrv12 I__7503 (
            .O(N__31217),
            .I(N_391_0));
    InMux I__7502 (
            .O(N__31210),
            .I(N__31207));
    LocalMux I__7501 (
            .O(N__31207),
            .I(\this_vga_signals.un1_M_this_state_q_18Z0Z_1 ));
    InMux I__7500 (
            .O(N__31204),
            .I(N__31194));
    InMux I__7499 (
            .O(N__31203),
            .I(N__31194));
    InMux I__7498 (
            .O(N__31202),
            .I(N__31191));
    InMux I__7497 (
            .O(N__31201),
            .I(N__31188));
    InMux I__7496 (
            .O(N__31200),
            .I(N__31185));
    CascadeMux I__7495 (
            .O(N__31199),
            .I(N__31182));
    LocalMux I__7494 (
            .O(N__31194),
            .I(N__31179));
    LocalMux I__7493 (
            .O(N__31191),
            .I(N__31176));
    LocalMux I__7492 (
            .O(N__31188),
            .I(N__31171));
    LocalMux I__7491 (
            .O(N__31185),
            .I(N__31171));
    InMux I__7490 (
            .O(N__31182),
            .I(N__31168));
    Span4Mux_v I__7489 (
            .O(N__31179),
            .I(N__31165));
    Span4Mux_v I__7488 (
            .O(N__31176),
            .I(N__31162));
    Span4Mux_v I__7487 (
            .O(N__31171),
            .I(N__31159));
    LocalMux I__7486 (
            .O(N__31168),
            .I(M_this_state_qZ0Z_11));
    Odrv4 I__7485 (
            .O(N__31165),
            .I(M_this_state_qZ0Z_11));
    Odrv4 I__7484 (
            .O(N__31162),
            .I(M_this_state_qZ0Z_11));
    Odrv4 I__7483 (
            .O(N__31159),
            .I(M_this_state_qZ0Z_11));
    InMux I__7482 (
            .O(N__31150),
            .I(N__31143));
    InMux I__7481 (
            .O(N__31149),
            .I(N__31143));
    CascadeMux I__7480 (
            .O(N__31148),
            .I(N__31140));
    LocalMux I__7479 (
            .O(N__31143),
            .I(N__31137));
    InMux I__7478 (
            .O(N__31140),
            .I(N__31134));
    Span4Mux_v I__7477 (
            .O(N__31137),
            .I(N__31129));
    LocalMux I__7476 (
            .O(N__31134),
            .I(N__31129));
    Span4Mux_h I__7475 (
            .O(N__31129),
            .I(N__31125));
    InMux I__7474 (
            .O(N__31128),
            .I(N__31122));
    Odrv4 I__7473 (
            .O(N__31125),
            .I(\this_vga_signals.N_387_0 ));
    LocalMux I__7472 (
            .O(N__31122),
            .I(\this_vga_signals.N_387_0 ));
    InMux I__7471 (
            .O(N__31117),
            .I(N__31108));
    InMux I__7470 (
            .O(N__31116),
            .I(N__31108));
    InMux I__7469 (
            .O(N__31115),
            .I(N__31108));
    LocalMux I__7468 (
            .O(N__31108),
            .I(N__31104));
    InMux I__7467 (
            .O(N__31107),
            .I(N__31097));
    Span4Mux_h I__7466 (
            .O(N__31104),
            .I(N__31094));
    InMux I__7465 (
            .O(N__31103),
            .I(N__31091));
    InMux I__7464 (
            .O(N__31102),
            .I(N__31088));
    InMux I__7463 (
            .O(N__31101),
            .I(N__31083));
    InMux I__7462 (
            .O(N__31100),
            .I(N__31083));
    LocalMux I__7461 (
            .O(N__31097),
            .I(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0 ));
    Odrv4 I__7460 (
            .O(N__31094),
            .I(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0 ));
    LocalMux I__7459 (
            .O(N__31091),
            .I(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0 ));
    LocalMux I__7458 (
            .O(N__31088),
            .I(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0 ));
    LocalMux I__7457 (
            .O(N__31083),
            .I(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0 ));
    InMux I__7456 (
            .O(N__31072),
            .I(N__31069));
    LocalMux I__7455 (
            .O(N__31069),
            .I(N_513));
    CascadeMux I__7454 (
            .O(N__31066),
            .I(N__31063));
    InMux I__7453 (
            .O(N__31063),
            .I(N__31060));
    LocalMux I__7452 (
            .O(N__31060),
            .I(M_this_data_count_q_s_7));
    CascadeMux I__7451 (
            .O(N__31057),
            .I(N__31054));
    InMux I__7450 (
            .O(N__31054),
            .I(N__31049));
    InMux I__7449 (
            .O(N__31053),
            .I(N__31046));
    InMux I__7448 (
            .O(N__31052),
            .I(N__31043));
    LocalMux I__7447 (
            .O(N__31049),
            .I(N__31040));
    LocalMux I__7446 (
            .O(N__31046),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__7445 (
            .O(N__31043),
            .I(M_this_data_count_qZ0Z_7));
    Odrv4 I__7444 (
            .O(N__31040),
            .I(M_this_data_count_qZ0Z_7));
    InMux I__7443 (
            .O(N__31033),
            .I(N__31030));
    LocalMux I__7442 (
            .O(N__31030),
            .I(M_this_data_count_q_s_8));
    CascadeMux I__7441 (
            .O(N__31027),
            .I(N_514_cascade_));
    InMux I__7440 (
            .O(N__31024),
            .I(N__31021));
    LocalMux I__7439 (
            .O(N__31021),
            .I(M_this_data_count_q_s_9));
    CascadeMux I__7438 (
            .O(N__31018),
            .I(N_515_cascade_));
    InMux I__7437 (
            .O(N__31015),
            .I(N__31012));
    LocalMux I__7436 (
            .O(N__31012),
            .I(N__31009));
    Span4Mux_v I__7435 (
            .O(N__31009),
            .I(N__31006));
    Odrv4 I__7434 (
            .O(N__31006),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_7 ));
    CascadeMux I__7433 (
            .O(N__31003),
            .I(\this_vga_signals.M_this_external_address_d_8_mZ0Z_7_cascade_ ));
    InMux I__7432 (
            .O(N__31000),
            .I(N__30997));
    LocalMux I__7431 (
            .O(N__30997),
            .I(un1_M_this_external_address_q_cry_6_c_RNIS2NBZ0));
    IoInMux I__7430 (
            .O(N__30994),
            .I(N__30991));
    LocalMux I__7429 (
            .O(N__30991),
            .I(N__30988));
    Span4Mux_s1_h I__7428 (
            .O(N__30988),
            .I(N__30985));
    Span4Mux_v I__7427 (
            .O(N__30985),
            .I(N__30982));
    Span4Mux_v I__7426 (
            .O(N__30982),
            .I(N__30979));
    Span4Mux_h I__7425 (
            .O(N__30979),
            .I(N__30975));
    InMux I__7424 (
            .O(N__30978),
            .I(N__30972));
    Span4Mux_h I__7423 (
            .O(N__30975),
            .I(N__30966));
    LocalMux I__7422 (
            .O(N__30972),
            .I(N__30966));
    InMux I__7421 (
            .O(N__30971),
            .I(N__30962));
    Span4Mux_v I__7420 (
            .O(N__30966),
            .I(N__30959));
    InMux I__7419 (
            .O(N__30965),
            .I(N__30956));
    LocalMux I__7418 (
            .O(N__30962),
            .I(M_this_external_address_qZ0Z_7));
    Odrv4 I__7417 (
            .O(N__30959),
            .I(M_this_external_address_qZ0Z_7));
    LocalMux I__7416 (
            .O(N__30956),
            .I(M_this_external_address_qZ0Z_7));
    CascadeMux I__7415 (
            .O(N__30949),
            .I(\this_vga_signals.M_this_external_address_d_5_mZ0Z_10_cascade_ ));
    InMux I__7414 (
            .O(N__30946),
            .I(N__30943));
    LocalMux I__7413 (
            .O(N__30943),
            .I(un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0));
    IoInMux I__7412 (
            .O(N__30940),
            .I(N__30937));
    LocalMux I__7411 (
            .O(N__30937),
            .I(N__30933));
    InMux I__7410 (
            .O(N__30936),
            .I(N__30929));
    Span12Mux_s11_v I__7409 (
            .O(N__30933),
            .I(N__30925));
    InMux I__7408 (
            .O(N__30932),
            .I(N__30922));
    LocalMux I__7407 (
            .O(N__30929),
            .I(N__30919));
    InMux I__7406 (
            .O(N__30928),
            .I(N__30916));
    Odrv12 I__7405 (
            .O(N__30925),
            .I(M_this_external_address_qZ0Z_10));
    LocalMux I__7404 (
            .O(N__30922),
            .I(M_this_external_address_qZ0Z_10));
    Odrv4 I__7403 (
            .O(N__30919),
            .I(M_this_external_address_qZ0Z_10));
    LocalMux I__7402 (
            .O(N__30916),
            .I(M_this_external_address_qZ0Z_10));
    InMux I__7401 (
            .O(N__30907),
            .I(N__30904));
    LocalMux I__7400 (
            .O(N__30904),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_10 ));
    IoInMux I__7399 (
            .O(N__30901),
            .I(N__30898));
    LocalMux I__7398 (
            .O(N__30898),
            .I(N__30895));
    Span4Mux_s2_v I__7397 (
            .O(N__30895),
            .I(N__30892));
    Span4Mux_v I__7396 (
            .O(N__30892),
            .I(N__30888));
    InMux I__7395 (
            .O(N__30891),
            .I(N__30884));
    Span4Mux_v I__7394 (
            .O(N__30888),
            .I(N__30880));
    InMux I__7393 (
            .O(N__30887),
            .I(N__30877));
    LocalMux I__7392 (
            .O(N__30884),
            .I(N__30874));
    InMux I__7391 (
            .O(N__30883),
            .I(N__30871));
    Odrv4 I__7390 (
            .O(N__30880),
            .I(M_this_external_address_qZ0Z_9));
    LocalMux I__7389 (
            .O(N__30877),
            .I(M_this_external_address_qZ0Z_9));
    Odrv12 I__7388 (
            .O(N__30874),
            .I(M_this_external_address_qZ0Z_9));
    LocalMux I__7387 (
            .O(N__30871),
            .I(M_this_external_address_qZ0Z_9));
    CascadeMux I__7386 (
            .O(N__30862),
            .I(N__30853));
    CascadeMux I__7385 (
            .O(N__30861),
            .I(N__30849));
    InMux I__7384 (
            .O(N__30860),
            .I(N__30844));
    InMux I__7383 (
            .O(N__30859),
            .I(N__30835));
    InMux I__7382 (
            .O(N__30858),
            .I(N__30828));
    InMux I__7381 (
            .O(N__30857),
            .I(N__30828));
    InMux I__7380 (
            .O(N__30856),
            .I(N__30828));
    InMux I__7379 (
            .O(N__30853),
            .I(N__30823));
    InMux I__7378 (
            .O(N__30852),
            .I(N__30823));
    InMux I__7377 (
            .O(N__30849),
            .I(N__30818));
    InMux I__7376 (
            .O(N__30848),
            .I(N__30818));
    InMux I__7375 (
            .O(N__30847),
            .I(N__30815));
    LocalMux I__7374 (
            .O(N__30844),
            .I(N__30812));
    InMux I__7373 (
            .O(N__30843),
            .I(N__30809));
    InMux I__7372 (
            .O(N__30842),
            .I(N__30806));
    InMux I__7371 (
            .O(N__30841),
            .I(N__30801));
    InMux I__7370 (
            .O(N__30840),
            .I(N__30801));
    InMux I__7369 (
            .O(N__30839),
            .I(N__30797));
    InMux I__7368 (
            .O(N__30838),
            .I(N__30794));
    LocalMux I__7367 (
            .O(N__30835),
            .I(N__30785));
    LocalMux I__7366 (
            .O(N__30828),
            .I(N__30785));
    LocalMux I__7365 (
            .O(N__30823),
            .I(N__30785));
    LocalMux I__7364 (
            .O(N__30818),
            .I(N__30785));
    LocalMux I__7363 (
            .O(N__30815),
            .I(N__30781));
    Span4Mux_h I__7362 (
            .O(N__30812),
            .I(N__30778));
    LocalMux I__7361 (
            .O(N__30809),
            .I(N__30771));
    LocalMux I__7360 (
            .O(N__30806),
            .I(N__30771));
    LocalMux I__7359 (
            .O(N__30801),
            .I(N__30771));
    InMux I__7358 (
            .O(N__30800),
            .I(N__30768));
    LocalMux I__7357 (
            .O(N__30797),
            .I(N__30765));
    LocalMux I__7356 (
            .O(N__30794),
            .I(N__30760));
    Span4Mux_v I__7355 (
            .O(N__30785),
            .I(N__30760));
    InMux I__7354 (
            .O(N__30784),
            .I(N__30757));
    Span4Mux_h I__7353 (
            .O(N__30781),
            .I(N__30745));
    Span4Mux_v I__7352 (
            .O(N__30778),
            .I(N__30745));
    Span4Mux_v I__7351 (
            .O(N__30771),
            .I(N__30745));
    LocalMux I__7350 (
            .O(N__30768),
            .I(N__30745));
    Span4Mux_v I__7349 (
            .O(N__30765),
            .I(N__30740));
    Span4Mux_v I__7348 (
            .O(N__30760),
            .I(N__30740));
    LocalMux I__7347 (
            .O(N__30757),
            .I(N__30737));
    InMux I__7346 (
            .O(N__30756),
            .I(N__30734));
    InMux I__7345 (
            .O(N__30755),
            .I(N__30731));
    InMux I__7344 (
            .O(N__30754),
            .I(N__30728));
    Span4Mux_v I__7343 (
            .O(N__30745),
            .I(N__30725));
    Span4Mux_h I__7342 (
            .O(N__30740),
            .I(N__30720));
    Span4Mux_h I__7341 (
            .O(N__30737),
            .I(N__30720));
    LocalMux I__7340 (
            .O(N__30734),
            .I(N__30715));
    LocalMux I__7339 (
            .O(N__30731),
            .I(N__30715));
    LocalMux I__7338 (
            .O(N__30728),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__7337 (
            .O(N__30725),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__7336 (
            .O(N__30720),
            .I(M_this_state_qZ0Z_6));
    Odrv12 I__7335 (
            .O(N__30715),
            .I(M_this_state_qZ0Z_6));
    InMux I__7334 (
            .O(N__30706),
            .I(N__30703));
    LocalMux I__7333 (
            .O(N__30703),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_9 ));
    InMux I__7332 (
            .O(N__30700),
            .I(N__30692));
    InMux I__7331 (
            .O(N__30699),
            .I(N__30689));
    CascadeMux I__7330 (
            .O(N__30698),
            .I(N__30686));
    InMux I__7329 (
            .O(N__30697),
            .I(N__30677));
    InMux I__7328 (
            .O(N__30696),
            .I(N__30677));
    InMux I__7327 (
            .O(N__30695),
            .I(N__30672));
    LocalMux I__7326 (
            .O(N__30692),
            .I(N__30664));
    LocalMux I__7325 (
            .O(N__30689),
            .I(N__30664));
    InMux I__7324 (
            .O(N__30686),
            .I(N__30661));
    InMux I__7323 (
            .O(N__30685),
            .I(N__30658));
    InMux I__7322 (
            .O(N__30684),
            .I(N__30655));
    InMux I__7321 (
            .O(N__30683),
            .I(N__30652));
    InMux I__7320 (
            .O(N__30682),
            .I(N__30649));
    LocalMux I__7319 (
            .O(N__30677),
            .I(N__30645));
    InMux I__7318 (
            .O(N__30676),
            .I(N__30640));
    InMux I__7317 (
            .O(N__30675),
            .I(N__30640));
    LocalMux I__7316 (
            .O(N__30672),
            .I(N__30637));
    InMux I__7315 (
            .O(N__30671),
            .I(N__30633));
    InMux I__7314 (
            .O(N__30670),
            .I(N__30630));
    InMux I__7313 (
            .O(N__30669),
            .I(N__30627));
    Span4Mux_v I__7312 (
            .O(N__30664),
            .I(N__30618));
    LocalMux I__7311 (
            .O(N__30661),
            .I(N__30618));
    LocalMux I__7310 (
            .O(N__30658),
            .I(N__30618));
    LocalMux I__7309 (
            .O(N__30655),
            .I(N__30618));
    LocalMux I__7308 (
            .O(N__30652),
            .I(N__30613));
    LocalMux I__7307 (
            .O(N__30649),
            .I(N__30613));
    CascadeMux I__7306 (
            .O(N__30648),
            .I(N__30610));
    Span4Mux_v I__7305 (
            .O(N__30645),
            .I(N__30602));
    LocalMux I__7304 (
            .O(N__30640),
            .I(N__30602));
    Span4Mux_v I__7303 (
            .O(N__30637),
            .I(N__30602));
    InMux I__7302 (
            .O(N__30636),
            .I(N__30599));
    LocalMux I__7301 (
            .O(N__30633),
            .I(N__30592));
    LocalMux I__7300 (
            .O(N__30630),
            .I(N__30592));
    LocalMux I__7299 (
            .O(N__30627),
            .I(N__30585));
    Span4Mux_v I__7298 (
            .O(N__30618),
            .I(N__30585));
    Span4Mux_v I__7297 (
            .O(N__30613),
            .I(N__30585));
    InMux I__7296 (
            .O(N__30610),
            .I(N__30582));
    InMux I__7295 (
            .O(N__30609),
            .I(N__30579));
    Span4Mux_h I__7294 (
            .O(N__30602),
            .I(N__30573));
    LocalMux I__7293 (
            .O(N__30599),
            .I(N__30573));
    InMux I__7292 (
            .O(N__30598),
            .I(N__30570));
    InMux I__7291 (
            .O(N__30597),
            .I(N__30567));
    Span12Mux_h I__7290 (
            .O(N__30592),
            .I(N__30564));
    Span4Mux_h I__7289 (
            .O(N__30585),
            .I(N__30561));
    LocalMux I__7288 (
            .O(N__30582),
            .I(N__30556));
    LocalMux I__7287 (
            .O(N__30579),
            .I(N__30556));
    InMux I__7286 (
            .O(N__30578),
            .I(N__30553));
    Span4Mux_h I__7285 (
            .O(N__30573),
            .I(N__30550));
    LocalMux I__7284 (
            .O(N__30570),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__7283 (
            .O(N__30567),
            .I(M_this_state_qZ0Z_5));
    Odrv12 I__7282 (
            .O(N__30564),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__7281 (
            .O(N__30561),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__7280 (
            .O(N__30556),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__7279 (
            .O(N__30553),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__7278 (
            .O(N__30550),
            .I(M_this_state_qZ0Z_5));
    InMux I__7277 (
            .O(N__30535),
            .I(N__30532));
    LocalMux I__7276 (
            .O(N__30532),
            .I(\this_vga_signals.M_this_external_address_d_5_mZ0Z_12 ));
    InMux I__7275 (
            .O(N__30529),
            .I(N__30515));
    InMux I__7274 (
            .O(N__30528),
            .I(N__30510));
    InMux I__7273 (
            .O(N__30527),
            .I(N__30510));
    InMux I__7272 (
            .O(N__30526),
            .I(N__30503));
    InMux I__7271 (
            .O(N__30525),
            .I(N__30503));
    InMux I__7270 (
            .O(N__30524),
            .I(N__30503));
    InMux I__7269 (
            .O(N__30523),
            .I(N__30496));
    InMux I__7268 (
            .O(N__30522),
            .I(N__30496));
    InMux I__7267 (
            .O(N__30521),
            .I(N__30496));
    InMux I__7266 (
            .O(N__30520),
            .I(N__30489));
    InMux I__7265 (
            .O(N__30519),
            .I(N__30489));
    InMux I__7264 (
            .O(N__30518),
            .I(N__30489));
    LocalMux I__7263 (
            .O(N__30515),
            .I(N__30476));
    LocalMux I__7262 (
            .O(N__30510),
            .I(N__30476));
    LocalMux I__7261 (
            .O(N__30503),
            .I(N__30476));
    LocalMux I__7260 (
            .O(N__30496),
            .I(N__30476));
    LocalMux I__7259 (
            .O(N__30489),
            .I(N__30476));
    InMux I__7258 (
            .O(N__30488),
            .I(N__30471));
    InMux I__7257 (
            .O(N__30487),
            .I(N__30471));
    Span4Mux_v I__7256 (
            .O(N__30476),
            .I(N__30467));
    LocalMux I__7255 (
            .O(N__30471),
            .I(N__30464));
    InMux I__7254 (
            .O(N__30470),
            .I(N__30461));
    Odrv4 I__7253 (
            .O(N__30467),
            .I(\this_vga_signals.un1_M_this_state_q_21_0 ));
    Odrv4 I__7252 (
            .O(N__30464),
            .I(\this_vga_signals.un1_M_this_state_q_21_0 ));
    LocalMux I__7251 (
            .O(N__30461),
            .I(\this_vga_signals.un1_M_this_state_q_21_0 ));
    CascadeMux I__7250 (
            .O(N__30454),
            .I(N__30451));
    InMux I__7249 (
            .O(N__30451),
            .I(N__30448));
    LocalMux I__7248 (
            .O(N__30448),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_12 ));
    InMux I__7247 (
            .O(N__30445),
            .I(N__30442));
    LocalMux I__7246 (
            .O(N__30442),
            .I(N__30439));
    Odrv4 I__7245 (
            .O(N__30439),
            .I(un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0));
    IoInMux I__7244 (
            .O(N__30436),
            .I(N__30433));
    LocalMux I__7243 (
            .O(N__30433),
            .I(N__30430));
    IoSpan4Mux I__7242 (
            .O(N__30430),
            .I(N__30427));
    Span4Mux_s2_h I__7241 (
            .O(N__30427),
            .I(N__30423));
    InMux I__7240 (
            .O(N__30426),
            .I(N__30418));
    Span4Mux_h I__7239 (
            .O(N__30423),
            .I(N__30415));
    InMux I__7238 (
            .O(N__30422),
            .I(N__30410));
    InMux I__7237 (
            .O(N__30421),
            .I(N__30410));
    LocalMux I__7236 (
            .O(N__30418),
            .I(N__30407));
    Odrv4 I__7235 (
            .O(N__30415),
            .I(M_this_external_address_qZ0Z_12));
    LocalMux I__7234 (
            .O(N__30410),
            .I(M_this_external_address_qZ0Z_12));
    Odrv4 I__7233 (
            .O(N__30407),
            .I(M_this_external_address_qZ0Z_12));
    InMux I__7232 (
            .O(N__30400),
            .I(N__30397));
    LocalMux I__7231 (
            .O(N__30397),
            .I(N__30394));
    Odrv4 I__7230 (
            .O(N__30394),
            .I(M_this_map_ram_write_data_3));
    InMux I__7229 (
            .O(N__30391),
            .I(N__30388));
    LocalMux I__7228 (
            .O(N__30388),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_1 ));
    CascadeMux I__7227 (
            .O(N__30385),
            .I(\this_vga_signals.M_this_external_address_d_8_mZ0Z_1_cascade_ ));
    InMux I__7226 (
            .O(N__30382),
            .I(N__30379));
    LocalMux I__7225 (
            .O(N__30379),
            .I(un1_M_this_external_address_q_cry_0_c_RNIGGGBZ0));
    IoInMux I__7224 (
            .O(N__30376),
            .I(N__30373));
    LocalMux I__7223 (
            .O(N__30373),
            .I(N__30370));
    IoSpan4Mux I__7222 (
            .O(N__30370),
            .I(N__30367));
    Sp12to4 I__7221 (
            .O(N__30367),
            .I(N__30364));
    Span12Mux_v I__7220 (
            .O(N__30364),
            .I(N__30358));
    InMux I__7219 (
            .O(N__30363),
            .I(N__30355));
    InMux I__7218 (
            .O(N__30362),
            .I(N__30352));
    InMux I__7217 (
            .O(N__30361),
            .I(N__30349));
    Odrv12 I__7216 (
            .O(N__30358),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__7215 (
            .O(N__30355),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__7214 (
            .O(N__30352),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__7213 (
            .O(N__30349),
            .I(M_this_external_address_qZ0Z_1));
    InMux I__7212 (
            .O(N__30340),
            .I(N__30337));
    LocalMux I__7211 (
            .O(N__30337),
            .I(N__30334));
    Span4Mux_v I__7210 (
            .O(N__30334),
            .I(N__30331));
    Span4Mux_h I__7209 (
            .O(N__30331),
            .I(N__30328));
    Odrv4 I__7208 (
            .O(N__30328),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_2 ));
    CascadeMux I__7207 (
            .O(N__30325),
            .I(\this_vga_signals.M_this_external_address_d_8_mZ0Z_2_cascade_ ));
    InMux I__7206 (
            .O(N__30322),
            .I(N__30319));
    LocalMux I__7205 (
            .O(N__30319),
            .I(un1_M_this_external_address_q_cry_1_c_RNIIJHBZ0));
    IoInMux I__7204 (
            .O(N__30316),
            .I(N__30313));
    LocalMux I__7203 (
            .O(N__30313),
            .I(N__30310));
    Span4Mux_s0_v I__7202 (
            .O(N__30310),
            .I(N__30307));
    Sp12to4 I__7201 (
            .O(N__30307),
            .I(N__30303));
    InMux I__7200 (
            .O(N__30306),
            .I(N__30300));
    Span12Mux_h I__7199 (
            .O(N__30303),
            .I(N__30296));
    LocalMux I__7198 (
            .O(N__30300),
            .I(N__30293));
    InMux I__7197 (
            .O(N__30299),
            .I(N__30289));
    Span12Mux_v I__7196 (
            .O(N__30296),
            .I(N__30284));
    Span12Mux_v I__7195 (
            .O(N__30293),
            .I(N__30284));
    InMux I__7194 (
            .O(N__30292),
            .I(N__30281));
    LocalMux I__7193 (
            .O(N__30289),
            .I(M_this_external_address_qZ0Z_2));
    Odrv12 I__7192 (
            .O(N__30284),
            .I(M_this_external_address_qZ0Z_2));
    LocalMux I__7191 (
            .O(N__30281),
            .I(M_this_external_address_qZ0Z_2));
    InMux I__7190 (
            .O(N__30274),
            .I(N__30271));
    LocalMux I__7189 (
            .O(N__30271),
            .I(N__30268));
    Odrv4 I__7188 (
            .O(N__30268),
            .I(\this_vga_signals.M_this_external_address_d_8_mZ0Z_4 ));
    CascadeMux I__7187 (
            .O(N__30265),
            .I(N__30262));
    InMux I__7186 (
            .O(N__30262),
            .I(N__30259));
    LocalMux I__7185 (
            .O(N__30259),
            .I(N__30256));
    Odrv4 I__7184 (
            .O(N__30256),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_4 ));
    InMux I__7183 (
            .O(N__30253),
            .I(N__30250));
    LocalMux I__7182 (
            .O(N__30250),
            .I(un1_M_this_external_address_q_cry_3_c_RNIMPJBZ0));
    IoInMux I__7181 (
            .O(N__30247),
            .I(N__30244));
    LocalMux I__7180 (
            .O(N__30244),
            .I(N__30241));
    IoSpan4Mux I__7179 (
            .O(N__30241),
            .I(N__30238));
    Span4Mux_s3_h I__7178 (
            .O(N__30238),
            .I(N__30233));
    InMux I__7177 (
            .O(N__30237),
            .I(N__30228));
    InMux I__7176 (
            .O(N__30236),
            .I(N__30228));
    Span4Mux_h I__7175 (
            .O(N__30233),
            .I(N__30222));
    LocalMux I__7174 (
            .O(N__30228),
            .I(N__30222));
    InMux I__7173 (
            .O(N__30227),
            .I(N__30219));
    Odrv4 I__7172 (
            .O(N__30222),
            .I(M_this_external_address_qZ0Z_4));
    LocalMux I__7171 (
            .O(N__30219),
            .I(M_this_external_address_qZ0Z_4));
    CascadeMux I__7170 (
            .O(N__30214),
            .I(\this_vga_signals.M_this_external_address_d_5_i_mZ0Z_15_cascade_ ));
    InMux I__7169 (
            .O(N__30211),
            .I(N__30208));
    LocalMux I__7168 (
            .O(N__30208),
            .I(un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0));
    IoInMux I__7167 (
            .O(N__30205),
            .I(N__30202));
    LocalMux I__7166 (
            .O(N__30202),
            .I(N__30199));
    Span12Mux_s9_h I__7165 (
            .O(N__30199),
            .I(N__30196));
    Span12Mux_v I__7164 (
            .O(N__30196),
            .I(N__30190));
    InMux I__7163 (
            .O(N__30195),
            .I(N__30187));
    InMux I__7162 (
            .O(N__30194),
            .I(N__30182));
    InMux I__7161 (
            .O(N__30193),
            .I(N__30182));
    Odrv12 I__7160 (
            .O(N__30190),
            .I(M_this_external_address_qZ0Z_15));
    LocalMux I__7159 (
            .O(N__30187),
            .I(M_this_external_address_qZ0Z_15));
    LocalMux I__7158 (
            .O(N__30182),
            .I(M_this_external_address_qZ0Z_15));
    InMux I__7157 (
            .O(N__30175),
            .I(N__30172));
    LocalMux I__7156 (
            .O(N__30172),
            .I(\this_vga_signals.M_this_external_address_q_i_mZ0Z_15 ));
    InMux I__7155 (
            .O(N__30169),
            .I(M_this_data_count_q_cry_10));
    InMux I__7154 (
            .O(N__30166),
            .I(M_this_data_count_q_cry_11));
    InMux I__7153 (
            .O(N__30163),
            .I(M_this_data_count_q_cry_12));
    SRMux I__7152 (
            .O(N__30160),
            .I(N__30157));
    LocalMux I__7151 (
            .O(N__30157),
            .I(N__30152));
    SRMux I__7150 (
            .O(N__30156),
            .I(N__30149));
    SRMux I__7149 (
            .O(N__30155),
            .I(N__30146));
    Span4Mux_s2_v I__7148 (
            .O(N__30152),
            .I(N__30141));
    LocalMux I__7147 (
            .O(N__30149),
            .I(N__30138));
    LocalMux I__7146 (
            .O(N__30146),
            .I(N__30135));
    SRMux I__7145 (
            .O(N__30145),
            .I(N__30132));
    IoInMux I__7144 (
            .O(N__30144),
            .I(N__30129));
    Span4Mux_h I__7143 (
            .O(N__30141),
            .I(N__30124));
    Span4Mux_h I__7142 (
            .O(N__30138),
            .I(N__30124));
    Span4Mux_s2_v I__7141 (
            .O(N__30135),
            .I(N__30119));
    LocalMux I__7140 (
            .O(N__30132),
            .I(N__30119));
    LocalMux I__7139 (
            .O(N__30129),
            .I(N__30112));
    Span4Mux_v I__7138 (
            .O(N__30124),
            .I(N__30107));
    Span4Mux_v I__7137 (
            .O(N__30119),
            .I(N__30107));
    SRMux I__7136 (
            .O(N__30118),
            .I(N__30103));
    SRMux I__7135 (
            .O(N__30117),
            .I(N__30100));
    SRMux I__7134 (
            .O(N__30116),
            .I(N__30097));
    SRMux I__7133 (
            .O(N__30115),
            .I(N__30094));
    IoSpan4Mux I__7132 (
            .O(N__30112),
            .I(N__30086));
    Span4Mux_v I__7131 (
            .O(N__30107),
            .I(N__30082));
    SRMux I__7130 (
            .O(N__30106),
            .I(N__30079));
    LocalMux I__7129 (
            .O(N__30103),
            .I(N__30066));
    LocalMux I__7128 (
            .O(N__30100),
            .I(N__30066));
    LocalMux I__7127 (
            .O(N__30097),
            .I(N__30061));
    LocalMux I__7126 (
            .O(N__30094),
            .I(N__30061));
    SRMux I__7125 (
            .O(N__30093),
            .I(N__30058));
    SRMux I__7124 (
            .O(N__30092),
            .I(N__30055));
    SRMux I__7123 (
            .O(N__30091),
            .I(N__30051));
    SRMux I__7122 (
            .O(N__30090),
            .I(N__30048));
    SRMux I__7121 (
            .O(N__30089),
            .I(N__30045));
    Span4Mux_s0_h I__7120 (
            .O(N__30086),
            .I(N__30035));
    SRMux I__7119 (
            .O(N__30085),
            .I(N__30032));
    Span4Mux_v I__7118 (
            .O(N__30082),
            .I(N__30025));
    LocalMux I__7117 (
            .O(N__30079),
            .I(N__30025));
    SRMux I__7116 (
            .O(N__30078),
            .I(N__30022));
    CascadeMux I__7115 (
            .O(N__30077),
            .I(N__30018));
    CascadeMux I__7114 (
            .O(N__30076),
            .I(N__30015));
    CascadeMux I__7113 (
            .O(N__30075),
            .I(N__30009));
    CascadeMux I__7112 (
            .O(N__30074),
            .I(N__30006));
    CascadeMux I__7111 (
            .O(N__30073),
            .I(N__30002));
    CascadeMux I__7110 (
            .O(N__30072),
            .I(N__29998));
    CascadeMux I__7109 (
            .O(N__30071),
            .I(N__29994));
    Span4Mux_v I__7108 (
            .O(N__30066),
            .I(N__29985));
    Span4Mux_v I__7107 (
            .O(N__30061),
            .I(N__29985));
    LocalMux I__7106 (
            .O(N__30058),
            .I(N__29985));
    LocalMux I__7105 (
            .O(N__30055),
            .I(N__29985));
    SRMux I__7104 (
            .O(N__30054),
            .I(N__29982));
    LocalMux I__7103 (
            .O(N__30051),
            .I(N__29977));
    LocalMux I__7102 (
            .O(N__30048),
            .I(N__29977));
    LocalMux I__7101 (
            .O(N__30045),
            .I(N__29974));
    SRMux I__7100 (
            .O(N__30044),
            .I(N__29971));
    SRMux I__7099 (
            .O(N__30043),
            .I(N__29968));
    SRMux I__7098 (
            .O(N__30042),
            .I(N__29963));
    SRMux I__7097 (
            .O(N__30041),
            .I(N__29958));
    SRMux I__7096 (
            .O(N__30040),
            .I(N__29955));
    SRMux I__7095 (
            .O(N__30039),
            .I(N__29952));
    SRMux I__7094 (
            .O(N__30038),
            .I(N__29949));
    Span4Mux_h I__7093 (
            .O(N__30035),
            .I(N__29942));
    LocalMux I__7092 (
            .O(N__30032),
            .I(N__29942));
    SRMux I__7091 (
            .O(N__30031),
            .I(N__29939));
    SRMux I__7090 (
            .O(N__30030),
            .I(N__29936));
    Span4Mux_v I__7089 (
            .O(N__30025),
            .I(N__29931));
    LocalMux I__7088 (
            .O(N__30022),
            .I(N__29928));
    InMux I__7087 (
            .O(N__30021),
            .I(N__29913));
    InMux I__7086 (
            .O(N__30018),
            .I(N__29913));
    InMux I__7085 (
            .O(N__30015),
            .I(N__29913));
    InMux I__7084 (
            .O(N__30014),
            .I(N__29913));
    InMux I__7083 (
            .O(N__30013),
            .I(N__29913));
    InMux I__7082 (
            .O(N__30012),
            .I(N__29913));
    InMux I__7081 (
            .O(N__30009),
            .I(N__29913));
    InMux I__7080 (
            .O(N__30006),
            .I(N__29898));
    InMux I__7079 (
            .O(N__30005),
            .I(N__29898));
    InMux I__7078 (
            .O(N__30002),
            .I(N__29898));
    InMux I__7077 (
            .O(N__30001),
            .I(N__29898));
    InMux I__7076 (
            .O(N__29998),
            .I(N__29898));
    InMux I__7075 (
            .O(N__29997),
            .I(N__29898));
    InMux I__7074 (
            .O(N__29994),
            .I(N__29898));
    Span4Mux_v I__7073 (
            .O(N__29985),
            .I(N__29895));
    LocalMux I__7072 (
            .O(N__29982),
            .I(N__29892));
    Span4Mux_v I__7071 (
            .O(N__29977),
            .I(N__29883));
    Span4Mux_h I__7070 (
            .O(N__29974),
            .I(N__29883));
    LocalMux I__7069 (
            .O(N__29971),
            .I(N__29883));
    LocalMux I__7068 (
            .O(N__29968),
            .I(N__29883));
    SRMux I__7067 (
            .O(N__29967),
            .I(N__29880));
    SRMux I__7066 (
            .O(N__29966),
            .I(N__29877));
    LocalMux I__7065 (
            .O(N__29963),
            .I(N__29873));
    SRMux I__7064 (
            .O(N__29962),
            .I(N__29870));
    SRMux I__7063 (
            .O(N__29961),
            .I(N__29866));
    LocalMux I__7062 (
            .O(N__29958),
            .I(N__29863));
    LocalMux I__7061 (
            .O(N__29955),
            .I(N__29860));
    LocalMux I__7060 (
            .O(N__29952),
            .I(N__29855));
    LocalMux I__7059 (
            .O(N__29949),
            .I(N__29855));
    SRMux I__7058 (
            .O(N__29948),
            .I(N__29852));
    SRMux I__7057 (
            .O(N__29947),
            .I(N__29849));
    Span4Mux_h I__7056 (
            .O(N__29942),
            .I(N__29843));
    LocalMux I__7055 (
            .O(N__29939),
            .I(N__29843));
    LocalMux I__7054 (
            .O(N__29936),
            .I(N__29840));
    SRMux I__7053 (
            .O(N__29935),
            .I(N__29837));
    IoInMux I__7052 (
            .O(N__29934),
            .I(N__29833));
    Span4Mux_v I__7051 (
            .O(N__29931),
            .I(N__29828));
    Span4Mux_v I__7050 (
            .O(N__29928),
            .I(N__29828));
    LocalMux I__7049 (
            .O(N__29913),
            .I(N__29822));
    LocalMux I__7048 (
            .O(N__29898),
            .I(N__29822));
    Span4Mux_v I__7047 (
            .O(N__29895),
            .I(N__29811));
    Span4Mux_v I__7046 (
            .O(N__29892),
            .I(N__29811));
    Span4Mux_v I__7045 (
            .O(N__29883),
            .I(N__29811));
    LocalMux I__7044 (
            .O(N__29880),
            .I(N__29811));
    LocalMux I__7043 (
            .O(N__29877),
            .I(N__29811));
    SRMux I__7042 (
            .O(N__29876),
            .I(N__29808));
    Span4Mux_v I__7041 (
            .O(N__29873),
            .I(N__29803));
    LocalMux I__7040 (
            .O(N__29870),
            .I(N__29803));
    SRMux I__7039 (
            .O(N__29869),
            .I(N__29800));
    LocalMux I__7038 (
            .O(N__29866),
            .I(N__29797));
    Span4Mux_s3_v I__7037 (
            .O(N__29863),
            .I(N__29786));
    Span4Mux_h I__7036 (
            .O(N__29860),
            .I(N__29786));
    Span4Mux_s3_v I__7035 (
            .O(N__29855),
            .I(N__29786));
    LocalMux I__7034 (
            .O(N__29852),
            .I(N__29786));
    LocalMux I__7033 (
            .O(N__29849),
            .I(N__29786));
    SRMux I__7032 (
            .O(N__29848),
            .I(N__29783));
    Span4Mux_v I__7031 (
            .O(N__29843),
            .I(N__29776));
    Span4Mux_h I__7030 (
            .O(N__29840),
            .I(N__29776));
    LocalMux I__7029 (
            .O(N__29837),
            .I(N__29776));
    SRMux I__7028 (
            .O(N__29836),
            .I(N__29773));
    LocalMux I__7027 (
            .O(N__29833),
            .I(N__29770));
    Span4Mux_h I__7026 (
            .O(N__29828),
            .I(N__29767));
    InMux I__7025 (
            .O(N__29827),
            .I(N__29763));
    Span4Mux_v I__7024 (
            .O(N__29822),
            .I(N__29760));
    Span4Mux_v I__7023 (
            .O(N__29811),
            .I(N__29751));
    LocalMux I__7022 (
            .O(N__29808),
            .I(N__29751));
    Span4Mux_v I__7021 (
            .O(N__29803),
            .I(N__29751));
    LocalMux I__7020 (
            .O(N__29800),
            .I(N__29751));
    Span4Mux_h I__7019 (
            .O(N__29797),
            .I(N__29740));
    Span4Mux_v I__7018 (
            .O(N__29786),
            .I(N__29740));
    LocalMux I__7017 (
            .O(N__29783),
            .I(N__29740));
    Span4Mux_v I__7016 (
            .O(N__29776),
            .I(N__29740));
    LocalMux I__7015 (
            .O(N__29773),
            .I(N__29740));
    Span12Mux_s8_h I__7014 (
            .O(N__29770),
            .I(N__29737));
    Span4Mux_h I__7013 (
            .O(N__29767),
            .I(N__29734));
    SRMux I__7012 (
            .O(N__29766),
            .I(N__29731));
    LocalMux I__7011 (
            .O(N__29763),
            .I(N__29728));
    Span4Mux_v I__7010 (
            .O(N__29760),
            .I(N__29725));
    Span4Mux_v I__7009 (
            .O(N__29751),
            .I(N__29720));
    Span4Mux_v I__7008 (
            .O(N__29740),
            .I(N__29720));
    Span12Mux_h I__7007 (
            .O(N__29737),
            .I(N__29717));
    Span4Mux_h I__7006 (
            .O(N__29734),
            .I(N__29714));
    LocalMux I__7005 (
            .O(N__29731),
            .I(N__29711));
    Span12Mux_v I__7004 (
            .O(N__29728),
            .I(N__29704));
    Sp12to4 I__7003 (
            .O(N__29725),
            .I(N__29704));
    Sp12to4 I__7002 (
            .O(N__29720),
            .I(N__29704));
    Odrv12 I__7001 (
            .O(N__29717),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7000 (
            .O(N__29714),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6999 (
            .O(N__29711),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6998 (
            .O(N__29704),
            .I(CONSTANT_ONE_NET));
    InMux I__6997 (
            .O(N__29695),
            .I(M_this_data_count_q_cry_13));
    InMux I__6996 (
            .O(N__29692),
            .I(M_this_data_count_q_cry_14));
    InMux I__6995 (
            .O(N__29689),
            .I(N__29686));
    LocalMux I__6994 (
            .O(N__29686),
            .I(N__29683));
    Span12Mux_v I__6993 (
            .O(N__29683),
            .I(N__29680));
    Span12Mux_v I__6992 (
            .O(N__29680),
            .I(N__29677));
    Odrv12 I__6991 (
            .O(N__29677),
            .I(M_this_map_ram_read_data_6));
    InMux I__6990 (
            .O(N__29674),
            .I(N__29669));
    CascadeMux I__6989 (
            .O(N__29673),
            .I(N__29666));
    CascadeMux I__6988 (
            .O(N__29672),
            .I(N__29663));
    LocalMux I__6987 (
            .O(N__29669),
            .I(N__29660));
    InMux I__6986 (
            .O(N__29666),
            .I(N__29657));
    InMux I__6985 (
            .O(N__29663),
            .I(N__29654));
    Span4Mux_h I__6984 (
            .O(N__29660),
            .I(N__29651));
    LocalMux I__6983 (
            .O(N__29657),
            .I(N__29646));
    LocalMux I__6982 (
            .O(N__29654),
            .I(N__29646));
    Span4Mux_h I__6981 (
            .O(N__29651),
            .I(N__29640));
    Span4Mux_v I__6980 (
            .O(N__29646),
            .I(N__29640));
    InMux I__6979 (
            .O(N__29645),
            .I(N__29637));
    Span4Mux_h I__6978 (
            .O(N__29640),
            .I(N__29634));
    LocalMux I__6977 (
            .O(N__29637),
            .I(N__29631));
    Span4Mux_h I__6976 (
            .O(N__29634),
            .I(N__29628));
    Span12Mux_h I__6975 (
            .O(N__29631),
            .I(N__29625));
    Odrv4 I__6974 (
            .O(N__29628),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv12 I__6973 (
            .O(N__29625),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    InMux I__6972 (
            .O(N__29620),
            .I(N__29613));
    InMux I__6971 (
            .O(N__29619),
            .I(N__29610));
    InMux I__6970 (
            .O(N__29618),
            .I(N__29607));
    InMux I__6969 (
            .O(N__29617),
            .I(N__29603));
    InMux I__6968 (
            .O(N__29616),
            .I(N__29600));
    LocalMux I__6967 (
            .O(N__29613),
            .I(N__29597));
    LocalMux I__6966 (
            .O(N__29610),
            .I(N__29592));
    LocalMux I__6965 (
            .O(N__29607),
            .I(N__29589));
    CascadeMux I__6964 (
            .O(N__29606),
            .I(N__29586));
    LocalMux I__6963 (
            .O(N__29603),
            .I(N__29581));
    LocalMux I__6962 (
            .O(N__29600),
            .I(N__29581));
    Span4Mux_v I__6961 (
            .O(N__29597),
            .I(N__29578));
    InMux I__6960 (
            .O(N__29596),
            .I(N__29575));
    InMux I__6959 (
            .O(N__29595),
            .I(N__29572));
    Span4Mux_h I__6958 (
            .O(N__29592),
            .I(N__29567));
    Span4Mux_h I__6957 (
            .O(N__29589),
            .I(N__29567));
    InMux I__6956 (
            .O(N__29586),
            .I(N__29564));
    Span4Mux_h I__6955 (
            .O(N__29581),
            .I(N__29561));
    Odrv4 I__6954 (
            .O(N__29578),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__6953 (
            .O(N__29575),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__6952 (
            .O(N__29572),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__6951 (
            .O(N__29567),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__6950 (
            .O(N__29564),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__6949 (
            .O(N__29561),
            .I(M_this_state_qZ0Z_7));
    InMux I__6948 (
            .O(N__29548),
            .I(N__29545));
    LocalMux I__6947 (
            .O(N__29545),
            .I(M_this_data_count_q_s_2));
    InMux I__6946 (
            .O(N__29542),
            .I(M_this_data_count_q_cry_1));
    InMux I__6945 (
            .O(N__29539),
            .I(N__29534));
    InMux I__6944 (
            .O(N__29538),
            .I(N__29531));
    InMux I__6943 (
            .O(N__29537),
            .I(N__29528));
    LocalMux I__6942 (
            .O(N__29534),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__6941 (
            .O(N__29531),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__6940 (
            .O(N__29528),
            .I(M_this_data_count_qZ0Z_3));
    CascadeMux I__6939 (
            .O(N__29521),
            .I(N__29518));
    InMux I__6938 (
            .O(N__29518),
            .I(N__29515));
    LocalMux I__6937 (
            .O(N__29515),
            .I(M_this_data_count_q_s_3));
    InMux I__6936 (
            .O(N__29512),
            .I(M_this_data_count_q_cry_2));
    CascadeMux I__6935 (
            .O(N__29509),
            .I(N__29505));
    InMux I__6934 (
            .O(N__29508),
            .I(N__29501));
    InMux I__6933 (
            .O(N__29505),
            .I(N__29498));
    InMux I__6932 (
            .O(N__29504),
            .I(N__29495));
    LocalMux I__6931 (
            .O(N__29501),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__6930 (
            .O(N__29498),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__6929 (
            .O(N__29495),
            .I(M_this_data_count_qZ0Z_4));
    InMux I__6928 (
            .O(N__29488),
            .I(N__29485));
    LocalMux I__6927 (
            .O(N__29485),
            .I(M_this_data_count_q_s_4));
    InMux I__6926 (
            .O(N__29482),
            .I(M_this_data_count_q_cry_3));
    InMux I__6925 (
            .O(N__29479),
            .I(N__29474));
    InMux I__6924 (
            .O(N__29478),
            .I(N__29469));
    InMux I__6923 (
            .O(N__29477),
            .I(N__29469));
    LocalMux I__6922 (
            .O(N__29474),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__6921 (
            .O(N__29469),
            .I(M_this_data_count_qZ0Z_5));
    CascadeMux I__6920 (
            .O(N__29464),
            .I(N__29461));
    InMux I__6919 (
            .O(N__29461),
            .I(N__29458));
    LocalMux I__6918 (
            .O(N__29458),
            .I(M_this_data_count_q_s_5));
    InMux I__6917 (
            .O(N__29455),
            .I(M_this_data_count_q_cry_4));
    CascadeMux I__6916 (
            .O(N__29452),
            .I(N__29449));
    InMux I__6915 (
            .O(N__29449),
            .I(N__29444));
    InMux I__6914 (
            .O(N__29448),
            .I(N__29439));
    InMux I__6913 (
            .O(N__29447),
            .I(N__29439));
    LocalMux I__6912 (
            .O(N__29444),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__6911 (
            .O(N__29439),
            .I(M_this_data_count_qZ0Z_6));
    CascadeMux I__6910 (
            .O(N__29434),
            .I(N__29431));
    InMux I__6909 (
            .O(N__29431),
            .I(N__29428));
    LocalMux I__6908 (
            .O(N__29428),
            .I(M_this_data_count_q_s_6));
    InMux I__6907 (
            .O(N__29425),
            .I(M_this_data_count_q_cry_5));
    InMux I__6906 (
            .O(N__29422),
            .I(M_this_data_count_q_cry_6));
    InMux I__6905 (
            .O(N__29419),
            .I(bfn_23_18_0_));
    InMux I__6904 (
            .O(N__29416),
            .I(M_this_data_count_q_cry_8));
    InMux I__6903 (
            .O(N__29413),
            .I(M_this_data_count_q_cry_9));
    InMux I__6902 (
            .O(N__29410),
            .I(N__29407));
    LocalMux I__6901 (
            .O(N__29407),
            .I(N_509));
    CascadeMux I__6900 (
            .O(N__29404),
            .I(N_510_cascade_));
    InMux I__6899 (
            .O(N__29401),
            .I(N__29398));
    LocalMux I__6898 (
            .O(N__29398),
            .I(N_511));
    InMux I__6897 (
            .O(N__29395),
            .I(N__29392));
    LocalMux I__6896 (
            .O(N__29392),
            .I(N_512));
    InMux I__6895 (
            .O(N__29389),
            .I(N__29386));
    LocalMux I__6894 (
            .O(N__29386),
            .I(N__29383));
    Span4Mux_v I__6893 (
            .O(N__29383),
            .I(N__29379));
    InMux I__6892 (
            .O(N__29382),
            .I(N__29374));
    Span4Mux_v I__6891 (
            .O(N__29379),
            .I(N__29371));
    InMux I__6890 (
            .O(N__29378),
            .I(N__29368));
    InMux I__6889 (
            .O(N__29377),
            .I(N__29365));
    LocalMux I__6888 (
            .O(N__29374),
            .I(M_this_data_count_qZ0Z_0));
    Odrv4 I__6887 (
            .O(N__29371),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__6886 (
            .O(N__29368),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__6885 (
            .O(N__29365),
            .I(M_this_data_count_qZ0Z_0));
    InMux I__6884 (
            .O(N__29356),
            .I(N__29351));
    InMux I__6883 (
            .O(N__29355),
            .I(N__29348));
    InMux I__6882 (
            .O(N__29354),
            .I(N__29345));
    LocalMux I__6881 (
            .O(N__29351),
            .I(N__29342));
    LocalMux I__6880 (
            .O(N__29348),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__6879 (
            .O(N__29345),
            .I(M_this_data_count_qZ0Z_1));
    Odrv4 I__6878 (
            .O(N__29342),
            .I(M_this_data_count_qZ0Z_1));
    InMux I__6877 (
            .O(N__29335),
            .I(N__29332));
    LocalMux I__6876 (
            .O(N__29332),
            .I(M_this_data_count_q_s_1));
    InMux I__6875 (
            .O(N__29329),
            .I(M_this_data_count_q_cry_0));
    CascadeMux I__6874 (
            .O(N__29326),
            .I(N__29322));
    InMux I__6873 (
            .O(N__29325),
            .I(N__29318));
    InMux I__6872 (
            .O(N__29322),
            .I(N__29315));
    InMux I__6871 (
            .O(N__29321),
            .I(N__29312));
    LocalMux I__6870 (
            .O(N__29318),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__6869 (
            .O(N__29315),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__6868 (
            .O(N__29312),
            .I(M_this_data_count_qZ0Z_2));
    IoInMux I__6867 (
            .O(N__29305),
            .I(N__29302));
    LocalMux I__6866 (
            .O(N__29302),
            .I(N__29299));
    Span4Mux_s0_v I__6865 (
            .O(N__29299),
            .I(N__29296));
    Sp12to4 I__6864 (
            .O(N__29296),
            .I(N__29292));
    InMux I__6863 (
            .O(N__29295),
            .I(N__29287));
    Span12Mux_s10_h I__6862 (
            .O(N__29292),
            .I(N__29284));
    InMux I__6861 (
            .O(N__29291),
            .I(N__29279));
    InMux I__6860 (
            .O(N__29290),
            .I(N__29279));
    LocalMux I__6859 (
            .O(N__29287),
            .I(N__29276));
    Odrv12 I__6858 (
            .O(N__29284),
            .I(M_this_external_address_qZ0Z_11));
    LocalMux I__6857 (
            .O(N__29279),
            .I(M_this_external_address_qZ0Z_11));
    Odrv4 I__6856 (
            .O(N__29276),
            .I(M_this_external_address_qZ0Z_11));
    InMux I__6855 (
            .O(N__29269),
            .I(N__29266));
    LocalMux I__6854 (
            .O(N__29266),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_11 ));
    CascadeMux I__6853 (
            .O(N__29263),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_3_cascade_ ));
    InMux I__6852 (
            .O(N__29260),
            .I(N__29257));
    LocalMux I__6851 (
            .O(N__29257),
            .I(N__29254));
    Odrv4 I__6850 (
            .O(N__29254),
            .I(un1_M_this_external_address_q_cry_2_c_RNIKMIBZ0));
    IoInMux I__6849 (
            .O(N__29251),
            .I(N__29248));
    LocalMux I__6848 (
            .O(N__29248),
            .I(N__29245));
    IoSpan4Mux I__6847 (
            .O(N__29245),
            .I(N__29242));
    Span4Mux_s1_h I__6846 (
            .O(N__29242),
            .I(N__29239));
    Span4Mux_v I__6845 (
            .O(N__29239),
            .I(N__29234));
    CascadeMux I__6844 (
            .O(N__29238),
            .I(N__29231));
    InMux I__6843 (
            .O(N__29237),
            .I(N__29227));
    Sp12to4 I__6842 (
            .O(N__29234),
            .I(N__29224));
    InMux I__6841 (
            .O(N__29231),
            .I(N__29219));
    InMux I__6840 (
            .O(N__29230),
            .I(N__29219));
    LocalMux I__6839 (
            .O(N__29227),
            .I(N__29216));
    Odrv12 I__6838 (
            .O(N__29224),
            .I(M_this_external_address_qZ0Z_3));
    LocalMux I__6837 (
            .O(N__29219),
            .I(M_this_external_address_qZ0Z_3));
    Odrv4 I__6836 (
            .O(N__29216),
            .I(M_this_external_address_qZ0Z_3));
    InMux I__6835 (
            .O(N__29209),
            .I(N__29206));
    LocalMux I__6834 (
            .O(N__29206),
            .I(\this_vga_signals.M_this_external_address_d_8_mZ0Z_3 ));
    InMux I__6833 (
            .O(N__29203),
            .I(N__29200));
    LocalMux I__6832 (
            .O(N__29200),
            .I(N__29197));
    Span12Mux_v I__6831 (
            .O(N__29197),
            .I(N__29194));
    Odrv12 I__6830 (
            .O(N__29194),
            .I(M_this_data_count_q_s_0));
    InMux I__6829 (
            .O(N__29191),
            .I(N__29182));
    InMux I__6828 (
            .O(N__29190),
            .I(N__29182));
    InMux I__6827 (
            .O(N__29189),
            .I(N__29177));
    InMux I__6826 (
            .O(N__29188),
            .I(N__29174));
    InMux I__6825 (
            .O(N__29187),
            .I(N__29171));
    LocalMux I__6824 (
            .O(N__29182),
            .I(N__29168));
    InMux I__6823 (
            .O(N__29181),
            .I(N__29165));
    InMux I__6822 (
            .O(N__29180),
            .I(N__29156));
    LocalMux I__6821 (
            .O(N__29177),
            .I(N__29153));
    LocalMux I__6820 (
            .O(N__29174),
            .I(N__29146));
    LocalMux I__6819 (
            .O(N__29171),
            .I(N__29146));
    Span4Mux_h I__6818 (
            .O(N__29168),
            .I(N__29146));
    LocalMux I__6817 (
            .O(N__29165),
            .I(N__29143));
    InMux I__6816 (
            .O(N__29164),
            .I(N__29140));
    InMux I__6815 (
            .O(N__29163),
            .I(N__29137));
    InMux I__6814 (
            .O(N__29162),
            .I(N__29134));
    InMux I__6813 (
            .O(N__29161),
            .I(N__29131));
    InMux I__6812 (
            .O(N__29160),
            .I(N__29128));
    InMux I__6811 (
            .O(N__29159),
            .I(N__29125));
    LocalMux I__6810 (
            .O(N__29156),
            .I(N__29122));
    Span4Mux_h I__6809 (
            .O(N__29153),
            .I(N__29119));
    Span4Mux_v I__6808 (
            .O(N__29146),
            .I(N__29114));
    Span4Mux_h I__6807 (
            .O(N__29143),
            .I(N__29114));
    LocalMux I__6806 (
            .O(N__29140),
            .I(N__29111));
    LocalMux I__6805 (
            .O(N__29137),
            .I(N__29102));
    LocalMux I__6804 (
            .O(N__29134),
            .I(N__29102));
    LocalMux I__6803 (
            .O(N__29131),
            .I(N__29102));
    LocalMux I__6802 (
            .O(N__29128),
            .I(N__29102));
    LocalMux I__6801 (
            .O(N__29125),
            .I(M_this_state_qZ0Z_10));
    Odrv4 I__6800 (
            .O(N__29122),
            .I(M_this_state_qZ0Z_10));
    Odrv4 I__6799 (
            .O(N__29119),
            .I(M_this_state_qZ0Z_10));
    Odrv4 I__6798 (
            .O(N__29114),
            .I(M_this_state_qZ0Z_10));
    Odrv12 I__6797 (
            .O(N__29111),
            .I(M_this_state_qZ0Z_10));
    Odrv4 I__6796 (
            .O(N__29102),
            .I(M_this_state_qZ0Z_10));
    CascadeMux I__6795 (
            .O(N__29089),
            .I(\this_vga_signals.N_292_cascade_ ));
    InMux I__6794 (
            .O(N__29086),
            .I(N__29083));
    LocalMux I__6793 (
            .O(N__29083),
            .I(N__29079));
    InMux I__6792 (
            .O(N__29082),
            .I(N__29076));
    Span4Mux_h I__6791 (
            .O(N__29079),
            .I(N__29073));
    LocalMux I__6790 (
            .O(N__29076),
            .I(N__29070));
    Odrv4 I__6789 (
            .O(N__29073),
            .I(\this_vga_signals.M_this_external_address_d_2_sqmuxaZ0 ));
    Odrv4 I__6788 (
            .O(N__29070),
            .I(\this_vga_signals.M_this_external_address_d_2_sqmuxaZ0 ));
    InMux I__6787 (
            .O(N__29065),
            .I(N__29062));
    LocalMux I__6786 (
            .O(N__29062),
            .I(M_this_state_d88_9));
    CascadeMux I__6785 (
            .O(N__29059),
            .I(N__29056));
    InMux I__6784 (
            .O(N__29056),
            .I(N__29053));
    LocalMux I__6783 (
            .O(N__29053),
            .I(N__29050));
    Odrv4 I__6782 (
            .O(N__29050),
            .I(N_506));
    InMux I__6781 (
            .O(N__29047),
            .I(N__29044));
    LocalMux I__6780 (
            .O(N__29044),
            .I(un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0));
    CascadeMux I__6779 (
            .O(N__29041),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_8_cascade_ ));
    IoInMux I__6778 (
            .O(N__29038),
            .I(N__29035));
    LocalMux I__6777 (
            .O(N__29035),
            .I(N__29032));
    Span4Mux_s1_v I__6776 (
            .O(N__29032),
            .I(N__29029));
    Sp12to4 I__6775 (
            .O(N__29029),
            .I(N__29025));
    CascadeMux I__6774 (
            .O(N__29028),
            .I(N__29022));
    Span12Mux_h I__6773 (
            .O(N__29025),
            .I(N__29017));
    InMux I__6772 (
            .O(N__29022),
            .I(N__29012));
    InMux I__6771 (
            .O(N__29021),
            .I(N__29012));
    InMux I__6770 (
            .O(N__29020),
            .I(N__29009));
    Odrv12 I__6769 (
            .O(N__29017),
            .I(M_this_external_address_qZ0Z_8));
    LocalMux I__6768 (
            .O(N__29012),
            .I(M_this_external_address_qZ0Z_8));
    LocalMux I__6767 (
            .O(N__29009),
            .I(M_this_external_address_qZ0Z_8));
    InMux I__6766 (
            .O(N__29002),
            .I(N__28999));
    LocalMux I__6765 (
            .O(N__28999),
            .I(\this_vga_signals.M_this_external_address_d_5_mZ0Z_8 ));
    CascadeMux I__6764 (
            .O(N__28996),
            .I(\this_vga_signals.M_this_external_address_d_8_mZ0Z_0_cascade_ ));
    InMux I__6763 (
            .O(N__28993),
            .I(N__28990));
    LocalMux I__6762 (
            .O(N__28990),
            .I(N__28987));
    Odrv12 I__6761 (
            .O(N__28987),
            .I(M_this_external_address_q_RNIE44V9Z0Z_0));
    IoInMux I__6760 (
            .O(N__28984),
            .I(N__28981));
    LocalMux I__6759 (
            .O(N__28981),
            .I(N__28978));
    IoSpan4Mux I__6758 (
            .O(N__28978),
            .I(N__28975));
    Span4Mux_s2_v I__6757 (
            .O(N__28975),
            .I(N__28972));
    Span4Mux_v I__6756 (
            .O(N__28972),
            .I(N__28968));
    InMux I__6755 (
            .O(N__28971),
            .I(N__28963));
    Span4Mux_v I__6754 (
            .O(N__28968),
            .I(N__28960));
    InMux I__6753 (
            .O(N__28967),
            .I(N__28955));
    InMux I__6752 (
            .O(N__28966),
            .I(N__28955));
    LocalMux I__6751 (
            .O(N__28963),
            .I(N__28952));
    Odrv4 I__6750 (
            .O(N__28960),
            .I(M_this_external_address_qZ0Z_0));
    LocalMux I__6749 (
            .O(N__28955),
            .I(M_this_external_address_qZ0Z_0));
    Odrv4 I__6748 (
            .O(N__28952),
            .I(M_this_external_address_qZ0Z_0));
    InMux I__6747 (
            .O(N__28945),
            .I(N__28942));
    LocalMux I__6746 (
            .O(N__28942),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_0 ));
    CascadeMux I__6745 (
            .O(N__28939),
            .I(N__28936));
    InMux I__6744 (
            .O(N__28936),
            .I(N__28933));
    LocalMux I__6743 (
            .O(N__28933),
            .I(N__28930));
    Odrv4 I__6742 (
            .O(N__28930),
            .I(\this_vga_signals.M_this_external_address_d_5_mZ0Z_9 ));
    InMux I__6741 (
            .O(N__28927),
            .I(N__28924));
    LocalMux I__6740 (
            .O(N__28924),
            .I(un1_M_this_external_address_q_cry_8_c_RNI09PBZ0));
    CascadeMux I__6739 (
            .O(N__28921),
            .I(\this_vga_signals.M_this_external_address_d_5_mZ0Z_11_cascade_ ));
    InMux I__6738 (
            .O(N__28918),
            .I(N__28915));
    LocalMux I__6737 (
            .O(N__28915),
            .I(N__28912));
    Odrv4 I__6736 (
            .O(N__28912),
            .I(un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0));
    InMux I__6735 (
            .O(N__28909),
            .I(bfn_22_21_0_));
    InMux I__6734 (
            .O(N__28906),
            .I(un1_M_this_external_address_q_cry_8));
    InMux I__6733 (
            .O(N__28903),
            .I(un1_M_this_external_address_q_cry_9));
    InMux I__6732 (
            .O(N__28900),
            .I(un1_M_this_external_address_q_cry_10));
    InMux I__6731 (
            .O(N__28897),
            .I(un1_M_this_external_address_q_cry_11));
    IoInMux I__6730 (
            .O(N__28894),
            .I(N__28891));
    LocalMux I__6729 (
            .O(N__28891),
            .I(N__28888));
    Span4Mux_s2_h I__6728 (
            .O(N__28888),
            .I(N__28885));
    Span4Mux_h I__6727 (
            .O(N__28885),
            .I(N__28881));
    InMux I__6726 (
            .O(N__28884),
            .I(N__28878));
    Span4Mux_h I__6725 (
            .O(N__28881),
            .I(N__28871));
    LocalMux I__6724 (
            .O(N__28878),
            .I(N__28871));
    InMux I__6723 (
            .O(N__28877),
            .I(N__28866));
    InMux I__6722 (
            .O(N__28876),
            .I(N__28866));
    Odrv4 I__6721 (
            .O(N__28871),
            .I(M_this_external_address_qZ0Z_13));
    LocalMux I__6720 (
            .O(N__28866),
            .I(M_this_external_address_qZ0Z_13));
    InMux I__6719 (
            .O(N__28861),
            .I(N__28858));
    LocalMux I__6718 (
            .O(N__28858),
            .I(N__28855));
    Odrv4 I__6717 (
            .O(N__28855),
            .I(un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0));
    InMux I__6716 (
            .O(N__28852),
            .I(un1_M_this_external_address_q_cry_12));
    IoInMux I__6715 (
            .O(N__28849),
            .I(N__28846));
    LocalMux I__6714 (
            .O(N__28846),
            .I(N__28843));
    Span4Mux_s3_h I__6713 (
            .O(N__28843),
            .I(N__28839));
    InMux I__6712 (
            .O(N__28842),
            .I(N__28835));
    Span4Mux_h I__6711 (
            .O(N__28839),
            .I(N__28832));
    CascadeMux I__6710 (
            .O(N__28838),
            .I(N__28829));
    LocalMux I__6709 (
            .O(N__28835),
            .I(N__28826));
    Span4Mux_h I__6708 (
            .O(N__28832),
            .I(N__28822));
    InMux I__6707 (
            .O(N__28829),
            .I(N__28819));
    Span4Mux_h I__6706 (
            .O(N__28826),
            .I(N__28816));
    InMux I__6705 (
            .O(N__28825),
            .I(N__28813));
    Odrv4 I__6704 (
            .O(N__28822),
            .I(M_this_external_address_qZ0Z_14));
    LocalMux I__6703 (
            .O(N__28819),
            .I(M_this_external_address_qZ0Z_14));
    Odrv4 I__6702 (
            .O(N__28816),
            .I(M_this_external_address_qZ0Z_14));
    LocalMux I__6701 (
            .O(N__28813),
            .I(M_this_external_address_qZ0Z_14));
    InMux I__6700 (
            .O(N__28804),
            .I(N__28801));
    LocalMux I__6699 (
            .O(N__28801),
            .I(N__28798));
    Span4Mux_h I__6698 (
            .O(N__28798),
            .I(N__28795));
    Odrv4 I__6697 (
            .O(N__28795),
            .I(un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0));
    InMux I__6696 (
            .O(N__28792),
            .I(un1_M_this_external_address_q_cry_13));
    InMux I__6695 (
            .O(N__28789),
            .I(un1_M_this_external_address_q_cry_14));
    CascadeMux I__6694 (
            .O(N__28786),
            .I(N__28781));
    InMux I__6693 (
            .O(N__28785),
            .I(N__28778));
    InMux I__6692 (
            .O(N__28784),
            .I(N__28775));
    InMux I__6691 (
            .O(N__28781),
            .I(N__28772));
    LocalMux I__6690 (
            .O(N__28778),
            .I(un1_M_this_state_q_16_0));
    LocalMux I__6689 (
            .O(N__28775),
            .I(un1_M_this_state_q_16_0));
    LocalMux I__6688 (
            .O(N__28772),
            .I(un1_M_this_state_q_16_0));
    InMux I__6687 (
            .O(N__28765),
            .I(un1_M_this_external_address_q_cry_0));
    InMux I__6686 (
            .O(N__28762),
            .I(un1_M_this_external_address_q_cry_1));
    InMux I__6685 (
            .O(N__28759),
            .I(un1_M_this_external_address_q_cry_2));
    InMux I__6684 (
            .O(N__28756),
            .I(un1_M_this_external_address_q_cry_3));
    IoInMux I__6683 (
            .O(N__28753),
            .I(N__28750));
    LocalMux I__6682 (
            .O(N__28750),
            .I(N__28745));
    CascadeMux I__6681 (
            .O(N__28749),
            .I(N__28741));
    CascadeMux I__6680 (
            .O(N__28748),
            .I(N__28738));
    Span12Mux_s4_h I__6679 (
            .O(N__28745),
            .I(N__28735));
    InMux I__6678 (
            .O(N__28744),
            .I(N__28732));
    InMux I__6677 (
            .O(N__28741),
            .I(N__28729));
    InMux I__6676 (
            .O(N__28738),
            .I(N__28726));
    Odrv12 I__6675 (
            .O(N__28735),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__6674 (
            .O(N__28732),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__6673 (
            .O(N__28729),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__6672 (
            .O(N__28726),
            .I(M_this_external_address_qZ0Z_5));
    InMux I__6671 (
            .O(N__28717),
            .I(N__28714));
    LocalMux I__6670 (
            .O(N__28714),
            .I(un1_M_this_external_address_q_cry_4_c_RNIOSKBZ0));
    InMux I__6669 (
            .O(N__28711),
            .I(un1_M_this_external_address_q_cry_4));
    IoInMux I__6668 (
            .O(N__28708),
            .I(N__28705));
    LocalMux I__6667 (
            .O(N__28705),
            .I(N__28702));
    Span4Mux_s2_h I__6666 (
            .O(N__28702),
            .I(N__28699));
    Span4Mux_v I__6665 (
            .O(N__28699),
            .I(N__28695));
    InMux I__6664 (
            .O(N__28698),
            .I(N__28691));
    Sp12to4 I__6663 (
            .O(N__28695),
            .I(N__28687));
    InMux I__6662 (
            .O(N__28694),
            .I(N__28684));
    LocalMux I__6661 (
            .O(N__28691),
            .I(N__28681));
    InMux I__6660 (
            .O(N__28690),
            .I(N__28678));
    Odrv12 I__6659 (
            .O(N__28687),
            .I(M_this_external_address_qZ0Z_6));
    LocalMux I__6658 (
            .O(N__28684),
            .I(M_this_external_address_qZ0Z_6));
    Odrv12 I__6657 (
            .O(N__28681),
            .I(M_this_external_address_qZ0Z_6));
    LocalMux I__6656 (
            .O(N__28678),
            .I(M_this_external_address_qZ0Z_6));
    InMux I__6655 (
            .O(N__28669),
            .I(N__28666));
    LocalMux I__6654 (
            .O(N__28666),
            .I(un1_M_this_external_address_q_cry_5_c_RNIQVLBZ0));
    InMux I__6653 (
            .O(N__28663),
            .I(un1_M_this_external_address_q_cry_5));
    InMux I__6652 (
            .O(N__28660),
            .I(un1_M_this_external_address_q_cry_6));
    CascadeMux I__6651 (
            .O(N__28657),
            .I(N_508_cascade_));
    InMux I__6650 (
            .O(N__28654),
            .I(N__28651));
    LocalMux I__6649 (
            .O(N__28651),
            .I(N__28648));
    Odrv4 I__6648 (
            .O(N__28648),
            .I(M_this_state_d88_11));
    CascadeMux I__6647 (
            .O(N__28645),
            .I(M_this_state_d88_11_cascade_));
    InMux I__6646 (
            .O(N__28642),
            .I(N__28639));
    LocalMux I__6645 (
            .O(N__28639),
            .I(N__28636));
    Odrv12 I__6644 (
            .O(N__28636),
            .I(M_this_state_d88_12));
    InMux I__6643 (
            .O(N__28633),
            .I(N__28630));
    LocalMux I__6642 (
            .O(N__28630),
            .I(N__28627));
    Odrv4 I__6641 (
            .O(N__28627),
            .I(N_436));
    InMux I__6640 (
            .O(N__28624),
            .I(N__28621));
    LocalMux I__6639 (
            .O(N__28621),
            .I(N__28618));
    Span4Mux_v I__6638 (
            .O(N__28618),
            .I(N__28615));
    Span4Mux_h I__6637 (
            .O(N__28615),
            .I(N__28612));
    Odrv4 I__6636 (
            .O(N__28612),
            .I(N_465));
    InMux I__6635 (
            .O(N__28609),
            .I(N__28606));
    LocalMux I__6634 (
            .O(N__28606),
            .I(N__28603));
    Span4Mux_h I__6633 (
            .O(N__28603),
            .I(N__28600));
    Odrv4 I__6632 (
            .O(N__28600),
            .I(N_435));
    CascadeMux I__6631 (
            .O(N__28597),
            .I(M_this_state_qsr_0_cascade_));
    InMux I__6630 (
            .O(N__28594),
            .I(N__28591));
    LocalMux I__6629 (
            .O(N__28591),
            .I(N__28588));
    Odrv4 I__6628 (
            .O(N__28588),
            .I(N_466));
    IoInMux I__6627 (
            .O(N__28585),
            .I(N__28582));
    LocalMux I__6626 (
            .O(N__28582),
            .I(N__28579));
    Span4Mux_s2_h I__6625 (
            .O(N__28579),
            .I(N__28575));
    CascadeMux I__6624 (
            .O(N__28578),
            .I(N__28571));
    Span4Mux_h I__6623 (
            .O(N__28575),
            .I(N__28568));
    InMux I__6622 (
            .O(N__28574),
            .I(N__28565));
    InMux I__6621 (
            .O(N__28571),
            .I(N__28562));
    Sp12to4 I__6620 (
            .O(N__28568),
            .I(N__28556));
    LocalMux I__6619 (
            .O(N__28565),
            .I(N__28551));
    LocalMux I__6618 (
            .O(N__28562),
            .I(N__28551));
    InMux I__6617 (
            .O(N__28561),
            .I(N__28544));
    InMux I__6616 (
            .O(N__28560),
            .I(N__28544));
    InMux I__6615 (
            .O(N__28559),
            .I(N__28544));
    Span12Mux_v I__6614 (
            .O(N__28556),
            .I(N__28541));
    Span4Mux_h I__6613 (
            .O(N__28551),
            .I(N__28538));
    LocalMux I__6612 (
            .O(N__28544),
            .I(N__28535));
    Odrv12 I__6611 (
            .O(N__28541),
            .I(led_c_1));
    Odrv4 I__6610 (
            .O(N__28538),
            .I(led_c_1));
    Odrv4 I__6609 (
            .O(N__28535),
            .I(led_c_1));
    InMux I__6608 (
            .O(N__28528),
            .I(N__28525));
    LocalMux I__6607 (
            .O(N__28525),
            .I(N__28520));
    InMux I__6606 (
            .O(N__28524),
            .I(N__28517));
    InMux I__6605 (
            .O(N__28523),
            .I(N__28514));
    Span4Mux_v I__6604 (
            .O(N__28520),
            .I(N__28509));
    LocalMux I__6603 (
            .O(N__28517),
            .I(N__28509));
    LocalMux I__6602 (
            .O(N__28514),
            .I(N__28506));
    Span4Mux_h I__6601 (
            .O(N__28509),
            .I(N__28501));
    Span4Mux_h I__6600 (
            .O(N__28506),
            .I(N__28498));
    InMux I__6599 (
            .O(N__28505),
            .I(N__28495));
    InMux I__6598 (
            .O(N__28504),
            .I(N__28492));
    Odrv4 I__6597 (
            .O(N__28501),
            .I(M_this_state_d88));
    Odrv4 I__6596 (
            .O(N__28498),
            .I(M_this_state_d88));
    LocalMux I__6595 (
            .O(N__28495),
            .I(M_this_state_d88));
    LocalMux I__6594 (
            .O(N__28492),
            .I(M_this_state_d88));
    InMux I__6593 (
            .O(N__28483),
            .I(N__28478));
    InMux I__6592 (
            .O(N__28482),
            .I(N__28475));
    InMux I__6591 (
            .O(N__28481),
            .I(N__28472));
    LocalMux I__6590 (
            .O(N__28478),
            .I(N__28462));
    LocalMux I__6589 (
            .O(N__28475),
            .I(N__28457));
    LocalMux I__6588 (
            .O(N__28472),
            .I(N__28457));
    InMux I__6587 (
            .O(N__28471),
            .I(N__28452));
    InMux I__6586 (
            .O(N__28470),
            .I(N__28452));
    InMux I__6585 (
            .O(N__28469),
            .I(N__28445));
    InMux I__6584 (
            .O(N__28468),
            .I(N__28445));
    InMux I__6583 (
            .O(N__28467),
            .I(N__28445));
    InMux I__6582 (
            .O(N__28466),
            .I(N__28440));
    InMux I__6581 (
            .O(N__28465),
            .I(N__28440));
    Span4Mux_h I__6580 (
            .O(N__28462),
            .I(N__28435));
    Span4Mux_h I__6579 (
            .O(N__28457),
            .I(N__28435));
    LocalMux I__6578 (
            .O(N__28452),
            .I(N__28432));
    LocalMux I__6577 (
            .O(N__28445),
            .I(N__28429));
    LocalMux I__6576 (
            .O(N__28440),
            .I(N__28426));
    Span4Mux_v I__6575 (
            .O(N__28435),
            .I(N__28423));
    Span4Mux_h I__6574 (
            .O(N__28432),
            .I(N__28420));
    Span4Mux_v I__6573 (
            .O(N__28429),
            .I(N__28417));
    Span12Mux_h I__6572 (
            .O(N__28426),
            .I(N__28414));
    Span4Mux_v I__6571 (
            .O(N__28423),
            .I(N__28411));
    Span4Mux_v I__6570 (
            .O(N__28420),
            .I(N__28408));
    Span4Mux_v I__6569 (
            .O(N__28417),
            .I(N__28405));
    Span12Mux_v I__6568 (
            .O(N__28414),
            .I(N__28402));
    Span4Mux_v I__6567 (
            .O(N__28411),
            .I(N__28399));
    Span4Mux_v I__6566 (
            .O(N__28408),
            .I(N__28396));
    IoSpan4Mux I__6565 (
            .O(N__28405),
            .I(N__28393));
    Odrv12 I__6564 (
            .O(N__28402),
            .I(rst_n_c));
    Odrv4 I__6563 (
            .O(N__28399),
            .I(rst_n_c));
    Odrv4 I__6562 (
            .O(N__28396),
            .I(rst_n_c));
    Odrv4 I__6561 (
            .O(N__28393),
            .I(rst_n_c));
    InMux I__6560 (
            .O(N__28384),
            .I(N__28381));
    LocalMux I__6559 (
            .O(N__28381),
            .I(N__28378));
    Span4Mux_h I__6558 (
            .O(N__28378),
            .I(N__28375));
    Odrv4 I__6557 (
            .O(N__28375),
            .I(\this_reset_cond.M_stage_qZ0Z_7 ));
    InMux I__6556 (
            .O(N__28372),
            .I(N__28369));
    LocalMux I__6555 (
            .O(N__28369),
            .I(\this_reset_cond.M_stage_qZ0Z_8 ));
    CascadeMux I__6554 (
            .O(N__28366),
            .I(N__28363));
    CascadeBuf I__6553 (
            .O(N__28363),
            .I(N__28360));
    CascadeMux I__6552 (
            .O(N__28360),
            .I(N__28357));
    CascadeBuf I__6551 (
            .O(N__28357),
            .I(N__28354));
    CascadeMux I__6550 (
            .O(N__28354),
            .I(N__28351));
    CascadeBuf I__6549 (
            .O(N__28351),
            .I(N__28348));
    CascadeMux I__6548 (
            .O(N__28348),
            .I(N__28345));
    CascadeBuf I__6547 (
            .O(N__28345),
            .I(N__28342));
    CascadeMux I__6546 (
            .O(N__28342),
            .I(N__28339));
    CascadeBuf I__6545 (
            .O(N__28339),
            .I(N__28336));
    CascadeMux I__6544 (
            .O(N__28336),
            .I(N__28333));
    CascadeBuf I__6543 (
            .O(N__28333),
            .I(N__28330));
    CascadeMux I__6542 (
            .O(N__28330),
            .I(N__28327));
    CascadeBuf I__6541 (
            .O(N__28327),
            .I(N__28324));
    CascadeMux I__6540 (
            .O(N__28324),
            .I(N__28321));
    CascadeBuf I__6539 (
            .O(N__28321),
            .I(N__28318));
    CascadeMux I__6538 (
            .O(N__28318),
            .I(N__28315));
    CascadeBuf I__6537 (
            .O(N__28315),
            .I(N__28312));
    CascadeMux I__6536 (
            .O(N__28312),
            .I(N__28309));
    CascadeBuf I__6535 (
            .O(N__28309),
            .I(N__28306));
    CascadeMux I__6534 (
            .O(N__28306),
            .I(N__28303));
    CascadeBuf I__6533 (
            .O(N__28303),
            .I(N__28300));
    CascadeMux I__6532 (
            .O(N__28300),
            .I(N__28297));
    CascadeBuf I__6531 (
            .O(N__28297),
            .I(N__28294));
    CascadeMux I__6530 (
            .O(N__28294),
            .I(N__28291));
    CascadeBuf I__6529 (
            .O(N__28291),
            .I(N__28288));
    CascadeMux I__6528 (
            .O(N__28288),
            .I(N__28285));
    CascadeBuf I__6527 (
            .O(N__28285),
            .I(N__28282));
    CascadeMux I__6526 (
            .O(N__28282),
            .I(N__28279));
    CascadeBuf I__6525 (
            .O(N__28279),
            .I(N__28276));
    CascadeMux I__6524 (
            .O(N__28276),
            .I(N__28273));
    InMux I__6523 (
            .O(N__28273),
            .I(N__28270));
    LocalMux I__6522 (
            .O(N__28270),
            .I(N__28267));
    Span4Mux_s1_v I__6521 (
            .O(N__28267),
            .I(N__28263));
    InMux I__6520 (
            .O(N__28266),
            .I(N__28259));
    Sp12to4 I__6519 (
            .O(N__28263),
            .I(N__28255));
    InMux I__6518 (
            .O(N__28262),
            .I(N__28252));
    LocalMux I__6517 (
            .O(N__28259),
            .I(N__28249));
    InMux I__6516 (
            .O(N__28258),
            .I(N__28246));
    Span12Mux_h I__6515 (
            .O(N__28255),
            .I(N__28243));
    LocalMux I__6514 (
            .O(N__28252),
            .I(N__28238));
    Span4Mux_h I__6513 (
            .O(N__28249),
            .I(N__28238));
    LocalMux I__6512 (
            .O(N__28246),
            .I(N__28233));
    Span12Mux_v I__6511 (
            .O(N__28243),
            .I(N__28233));
    Odrv4 I__6510 (
            .O(N__28238),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv12 I__6509 (
            .O(N__28233),
            .I(M_this_sprites_address_qZ0Z_3));
    CascadeMux I__6508 (
            .O(N__28228),
            .I(N__28223));
    InMux I__6507 (
            .O(N__28227),
            .I(N__28217));
    InMux I__6506 (
            .O(N__28226),
            .I(N__28214));
    InMux I__6505 (
            .O(N__28223),
            .I(N__28208));
    CascadeMux I__6504 (
            .O(N__28222),
            .I(N__28204));
    InMux I__6503 (
            .O(N__28221),
            .I(N__28200));
    InMux I__6502 (
            .O(N__28220),
            .I(N__28195));
    LocalMux I__6501 (
            .O(N__28217),
            .I(N__28190));
    LocalMux I__6500 (
            .O(N__28214),
            .I(N__28190));
    InMux I__6499 (
            .O(N__28213),
            .I(N__28185));
    InMux I__6498 (
            .O(N__28212),
            .I(N__28185));
    InMux I__6497 (
            .O(N__28211),
            .I(N__28182));
    LocalMux I__6496 (
            .O(N__28208),
            .I(N__28179));
    InMux I__6495 (
            .O(N__28207),
            .I(N__28176));
    InMux I__6494 (
            .O(N__28204),
            .I(N__28171));
    InMux I__6493 (
            .O(N__28203),
            .I(N__28171));
    LocalMux I__6492 (
            .O(N__28200),
            .I(N__28167));
    InMux I__6491 (
            .O(N__28199),
            .I(N__28164));
    InMux I__6490 (
            .O(N__28198),
            .I(N__28157));
    LocalMux I__6489 (
            .O(N__28195),
            .I(N__28150));
    Span4Mux_v I__6488 (
            .O(N__28190),
            .I(N__28150));
    LocalMux I__6487 (
            .O(N__28185),
            .I(N__28150));
    LocalMux I__6486 (
            .O(N__28182),
            .I(N__28145));
    Span4Mux_h I__6485 (
            .O(N__28179),
            .I(N__28145));
    LocalMux I__6484 (
            .O(N__28176),
            .I(N__28140));
    LocalMux I__6483 (
            .O(N__28171),
            .I(N__28140));
    InMux I__6482 (
            .O(N__28170),
            .I(N__28137));
    Span4Mux_v I__6481 (
            .O(N__28167),
            .I(N__28132));
    LocalMux I__6480 (
            .O(N__28164),
            .I(N__28132));
    InMux I__6479 (
            .O(N__28163),
            .I(N__28127));
    InMux I__6478 (
            .O(N__28162),
            .I(N__28127));
    InMux I__6477 (
            .O(N__28161),
            .I(N__28124));
    InMux I__6476 (
            .O(N__28160),
            .I(N__28121));
    LocalMux I__6475 (
            .O(N__28157),
            .I(N__28116));
    Span4Mux_v I__6474 (
            .O(N__28150),
            .I(N__28116));
    Sp12to4 I__6473 (
            .O(N__28145),
            .I(N__28111));
    Span12Mux_h I__6472 (
            .O(N__28140),
            .I(N__28111));
    LocalMux I__6471 (
            .O(N__28137),
            .I(N__28104));
    Span4Mux_h I__6470 (
            .O(N__28132),
            .I(N__28104));
    LocalMux I__6469 (
            .O(N__28127),
            .I(N__28104));
    LocalMux I__6468 (
            .O(N__28124),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__6467 (
            .O(N__28121),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__6466 (
            .O(N__28116),
            .I(M_this_state_qZ0Z_2));
    Odrv12 I__6465 (
            .O(N__28111),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__6464 (
            .O(N__28104),
            .I(M_this_state_qZ0Z_2));
    InMux I__6463 (
            .O(N__28093),
            .I(N__28090));
    LocalMux I__6462 (
            .O(N__28090),
            .I(N__28087));
    Span4Mux_h I__6461 (
            .O(N__28087),
            .I(N__28084));
    Odrv4 I__6460 (
            .O(N__28084),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3 ));
    CascadeMux I__6459 (
            .O(N__28081),
            .I(M_this_state_d88_1_cascade_));
    InMux I__6458 (
            .O(N__28078),
            .I(N__28069));
    InMux I__6457 (
            .O(N__28077),
            .I(N__28069));
    InMux I__6456 (
            .O(N__28076),
            .I(N__28064));
    InMux I__6455 (
            .O(N__28075),
            .I(N__28064));
    InMux I__6454 (
            .O(N__28074),
            .I(N__28061));
    LocalMux I__6453 (
            .O(N__28069),
            .I(N__28056));
    LocalMux I__6452 (
            .O(N__28064),
            .I(N__28056));
    LocalMux I__6451 (
            .O(N__28061),
            .I(N__28053));
    Odrv4 I__6450 (
            .O(N__28056),
            .I(\this_vga_signals.N_390_0 ));
    Odrv12 I__6449 (
            .O(N__28053),
            .I(\this_vga_signals.N_390_0 ));
    CascadeMux I__6448 (
            .O(N__28048),
            .I(M_this_state_d88_12_cascade_));
    CascadeMux I__6447 (
            .O(N__28045),
            .I(N_507_cascade_));
    InMux I__6446 (
            .O(N__28042),
            .I(N__28037));
    InMux I__6445 (
            .O(N__28041),
            .I(N__28032));
    CascadeMux I__6444 (
            .O(N__28040),
            .I(N__28028));
    LocalMux I__6443 (
            .O(N__28037),
            .I(N__28024));
    InMux I__6442 (
            .O(N__28036),
            .I(N__28021));
    InMux I__6441 (
            .O(N__28035),
            .I(N__28018));
    LocalMux I__6440 (
            .O(N__28032),
            .I(N__28014));
    InMux I__6439 (
            .O(N__28031),
            .I(N__28011));
    InMux I__6438 (
            .O(N__28028),
            .I(N__28006));
    InMux I__6437 (
            .O(N__28027),
            .I(N__28006));
    Span4Mux_h I__6436 (
            .O(N__28024),
            .I(N__28001));
    LocalMux I__6435 (
            .O(N__28021),
            .I(N__28001));
    LocalMux I__6434 (
            .O(N__28018),
            .I(N__27998));
    InMux I__6433 (
            .O(N__28017),
            .I(N__27995));
    Span4Mux_h I__6432 (
            .O(N__28014),
            .I(N__27991));
    LocalMux I__6431 (
            .O(N__28011),
            .I(N__27982));
    LocalMux I__6430 (
            .O(N__28006),
            .I(N__27982));
    Span4Mux_v I__6429 (
            .O(N__28001),
            .I(N__27982));
    Span4Mux_h I__6428 (
            .O(N__27998),
            .I(N__27982));
    LocalMux I__6427 (
            .O(N__27995),
            .I(N__27979));
    InMux I__6426 (
            .O(N__27994),
            .I(N__27976));
    Span4Mux_h I__6425 (
            .O(N__27991),
            .I(N__27973));
    Span4Mux_h I__6424 (
            .O(N__27982),
            .I(N__27970));
    Odrv12 I__6423 (
            .O(N__27979),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__6422 (
            .O(N__27976),
            .I(M_this_state_qZ0Z_12));
    Odrv4 I__6421 (
            .O(N__27973),
            .I(M_this_state_qZ0Z_12));
    Odrv4 I__6420 (
            .O(N__27970),
            .I(M_this_state_qZ0Z_12));
    InMux I__6419 (
            .O(N__27961),
            .I(N__27957));
    InMux I__6418 (
            .O(N__27960),
            .I(N__27954));
    LocalMux I__6417 (
            .O(N__27957),
            .I(N__27951));
    LocalMux I__6416 (
            .O(N__27954),
            .I(\this_vga_signals.N_293_1 ));
    Odrv4 I__6415 (
            .O(N__27951),
            .I(\this_vga_signals.N_293_1 ));
    CascadeMux I__6414 (
            .O(N__27946),
            .I(N__27941));
    InMux I__6413 (
            .O(N__27945),
            .I(N__27937));
    CascadeMux I__6412 (
            .O(N__27944),
            .I(N__27932));
    InMux I__6411 (
            .O(N__27941),
            .I(N__27929));
    InMux I__6410 (
            .O(N__27940),
            .I(N__27926));
    LocalMux I__6409 (
            .O(N__27937),
            .I(N__27921));
    InMux I__6408 (
            .O(N__27936),
            .I(N__27916));
    InMux I__6407 (
            .O(N__27935),
            .I(N__27916));
    InMux I__6406 (
            .O(N__27932),
            .I(N__27913));
    LocalMux I__6405 (
            .O(N__27929),
            .I(N__27910));
    LocalMux I__6404 (
            .O(N__27926),
            .I(N__27907));
    InMux I__6403 (
            .O(N__27925),
            .I(N__27902));
    InMux I__6402 (
            .O(N__27924),
            .I(N__27902));
    Span4Mux_v I__6401 (
            .O(N__27921),
            .I(N__27899));
    LocalMux I__6400 (
            .O(N__27916),
            .I(N__27894));
    LocalMux I__6399 (
            .O(N__27913),
            .I(N__27894));
    Span4Mux_v I__6398 (
            .O(N__27910),
            .I(N__27891));
    Span4Mux_v I__6397 (
            .O(N__27907),
            .I(N__27888));
    LocalMux I__6396 (
            .O(N__27902),
            .I(N__27885));
    Span4Mux_h I__6395 (
            .O(N__27899),
            .I(N__27878));
    Span4Mux_v I__6394 (
            .O(N__27894),
            .I(N__27878));
    Span4Mux_h I__6393 (
            .O(N__27891),
            .I(N__27878));
    Odrv4 I__6392 (
            .O(N__27888),
            .I(M_this_state_qZ0Z_15));
    Odrv12 I__6391 (
            .O(N__27885),
            .I(M_this_state_qZ0Z_15));
    Odrv4 I__6390 (
            .O(N__27878),
            .I(M_this_state_qZ0Z_15));
    InMux I__6389 (
            .O(N__27871),
            .I(N__27868));
    LocalMux I__6388 (
            .O(N__27868),
            .I(N__27865));
    Span4Mux_h I__6387 (
            .O(N__27865),
            .I(N__27861));
    InMux I__6386 (
            .O(N__27864),
            .I(N__27858));
    Span4Mux_v I__6385 (
            .O(N__27861),
            .I(N__27855));
    LocalMux I__6384 (
            .O(N__27858),
            .I(N__27852));
    Odrv4 I__6383 (
            .O(N__27855),
            .I(\this_vga_signals.M_this_map_ram_write_data_1_sqmuxa ));
    Odrv12 I__6382 (
            .O(N__27852),
            .I(\this_vga_signals.M_this_map_ram_write_data_1_sqmuxa ));
    CascadeMux I__6381 (
            .O(N__27847),
            .I(\this_vga_signals.N_293_cascade_ ));
    InMux I__6380 (
            .O(N__27844),
            .I(N__27841));
    LocalMux I__6379 (
            .O(N__27841),
            .I(N__27838));
    Span4Mux_v I__6378 (
            .O(N__27838),
            .I(N__27835));
    Span4Mux_v I__6377 (
            .O(N__27835),
            .I(N__27832));
    Span4Mux_h I__6376 (
            .O(N__27832),
            .I(N__27829));
    Odrv4 I__6375 (
            .O(N__27829),
            .I(M_this_map_ram_read_data_7));
    InMux I__6374 (
            .O(N__27826),
            .I(N__27815));
    InMux I__6373 (
            .O(N__27825),
            .I(N__27812));
    InMux I__6372 (
            .O(N__27824),
            .I(N__27809));
    InMux I__6371 (
            .O(N__27823),
            .I(N__27806));
    InMux I__6370 (
            .O(N__27822),
            .I(N__27795));
    InMux I__6369 (
            .O(N__27821),
            .I(N__27795));
    InMux I__6368 (
            .O(N__27820),
            .I(N__27792));
    InMux I__6367 (
            .O(N__27819),
            .I(N__27789));
    InMux I__6366 (
            .O(N__27818),
            .I(N__27786));
    LocalMux I__6365 (
            .O(N__27815),
            .I(N__27781));
    LocalMux I__6364 (
            .O(N__27812),
            .I(N__27781));
    LocalMux I__6363 (
            .O(N__27809),
            .I(N__27776));
    LocalMux I__6362 (
            .O(N__27806),
            .I(N__27776));
    InMux I__6361 (
            .O(N__27805),
            .I(N__27773));
    InMux I__6360 (
            .O(N__27804),
            .I(N__27770));
    InMux I__6359 (
            .O(N__27803),
            .I(N__27763));
    InMux I__6358 (
            .O(N__27802),
            .I(N__27763));
    InMux I__6357 (
            .O(N__27801),
            .I(N__27763));
    InMux I__6356 (
            .O(N__27800),
            .I(N__27759));
    LocalMux I__6355 (
            .O(N__27795),
            .I(N__27754));
    LocalMux I__6354 (
            .O(N__27792),
            .I(N__27754));
    LocalMux I__6353 (
            .O(N__27789),
            .I(N__27747));
    LocalMux I__6352 (
            .O(N__27786),
            .I(N__27747));
    Span4Mux_v I__6351 (
            .O(N__27781),
            .I(N__27747));
    Span4Mux_h I__6350 (
            .O(N__27776),
            .I(N__27744));
    LocalMux I__6349 (
            .O(N__27773),
            .I(N__27737));
    LocalMux I__6348 (
            .O(N__27770),
            .I(N__27737));
    LocalMux I__6347 (
            .O(N__27763),
            .I(N__27737));
    InMux I__6346 (
            .O(N__27762),
            .I(N__27734));
    LocalMux I__6345 (
            .O(N__27759),
            .I(N__27729));
    Span4Mux_v I__6344 (
            .O(N__27754),
            .I(N__27729));
    Span4Mux_h I__6343 (
            .O(N__27747),
            .I(N__27724));
    Span4Mux_v I__6342 (
            .O(N__27744),
            .I(N__27724));
    Span12Mux_v I__6341 (
            .O(N__27737),
            .I(N__27719));
    LocalMux I__6340 (
            .O(N__27734),
            .I(N__27719));
    Sp12to4 I__6339 (
            .O(N__27729),
            .I(N__27716));
    Span4Mux_h I__6338 (
            .O(N__27724),
            .I(N__27713));
    Span12Mux_h I__6337 (
            .O(N__27719),
            .I(N__27710));
    Odrv12 I__6336 (
            .O(N__27716),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__6335 (
            .O(N__27713),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv12 I__6334 (
            .O(N__27710),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    InMux I__6333 (
            .O(N__27703),
            .I(N__27700));
    LocalMux I__6332 (
            .O(N__27700),
            .I(\this_vga_signals.M_this_external_address_d_8_mZ0Z_5 ));
    CascadeMux I__6331 (
            .O(N__27697),
            .I(N__27694));
    InMux I__6330 (
            .O(N__27694),
            .I(N__27691));
    LocalMux I__6329 (
            .O(N__27691),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_5 ));
    InMux I__6328 (
            .O(N__27688),
            .I(N__27685));
    LocalMux I__6327 (
            .O(N__27685),
            .I(N__27682));
    Odrv12 I__6326 (
            .O(N__27682),
            .I(\this_vga_signals.M_this_external_address_q_mZ0Z_6 ));
    CascadeMux I__6325 (
            .O(N__27679),
            .I(\this_vga_signals.M_this_external_address_d_8_mZ0Z_6_cascade_ ));
    CascadeMux I__6324 (
            .O(N__27676),
            .I(N__27673));
    CascadeBuf I__6323 (
            .O(N__27673),
            .I(N__27670));
    CascadeMux I__6322 (
            .O(N__27670),
            .I(N__27667));
    InMux I__6321 (
            .O(N__27667),
            .I(N__27664));
    LocalMux I__6320 (
            .O(N__27664),
            .I(N__27661));
    Span4Mux_s1_v I__6319 (
            .O(N__27661),
            .I(N__27658));
    Span4Mux_h I__6318 (
            .O(N__27658),
            .I(N__27652));
    InMux I__6317 (
            .O(N__27657),
            .I(N__27649));
    InMux I__6316 (
            .O(N__27656),
            .I(N__27646));
    InMux I__6315 (
            .O(N__27655),
            .I(N__27643));
    Span4Mux_v I__6314 (
            .O(N__27652),
            .I(N__27640));
    LocalMux I__6313 (
            .O(N__27649),
            .I(M_this_map_address_qZ0Z_8));
    LocalMux I__6312 (
            .O(N__27646),
            .I(M_this_map_address_qZ0Z_8));
    LocalMux I__6311 (
            .O(N__27643),
            .I(M_this_map_address_qZ0Z_8));
    Odrv4 I__6310 (
            .O(N__27640),
            .I(M_this_map_address_qZ0Z_8));
    InMux I__6309 (
            .O(N__27631),
            .I(N__27628));
    LocalMux I__6308 (
            .O(N__27628),
            .I(N__27618));
    InMux I__6307 (
            .O(N__27627),
            .I(N__27615));
    InMux I__6306 (
            .O(N__27626),
            .I(N__27612));
    CascadeMux I__6305 (
            .O(N__27625),
            .I(N__27608));
    InMux I__6304 (
            .O(N__27624),
            .I(N__27604));
    InMux I__6303 (
            .O(N__27623),
            .I(N__27600));
    CascadeMux I__6302 (
            .O(N__27622),
            .I(N__27594));
    InMux I__6301 (
            .O(N__27621),
            .I(N__27591));
    Span4Mux_v I__6300 (
            .O(N__27618),
            .I(N__27586));
    LocalMux I__6299 (
            .O(N__27615),
            .I(N__27586));
    LocalMux I__6298 (
            .O(N__27612),
            .I(N__27583));
    InMux I__6297 (
            .O(N__27611),
            .I(N__27578));
    InMux I__6296 (
            .O(N__27608),
            .I(N__27578));
    CascadeMux I__6295 (
            .O(N__27607),
            .I(N__27575));
    LocalMux I__6294 (
            .O(N__27604),
            .I(N__27572));
    InMux I__6293 (
            .O(N__27603),
            .I(N__27569));
    LocalMux I__6292 (
            .O(N__27600),
            .I(N__27566));
    InMux I__6291 (
            .O(N__27599),
            .I(N__27563));
    InMux I__6290 (
            .O(N__27598),
            .I(N__27558));
    InMux I__6289 (
            .O(N__27597),
            .I(N__27558));
    InMux I__6288 (
            .O(N__27594),
            .I(N__27555));
    LocalMux I__6287 (
            .O(N__27591),
            .I(N__27545));
    Span4Mux_h I__6286 (
            .O(N__27586),
            .I(N__27545));
    Span4Mux_v I__6285 (
            .O(N__27583),
            .I(N__27545));
    LocalMux I__6284 (
            .O(N__27578),
            .I(N__27545));
    InMux I__6283 (
            .O(N__27575),
            .I(N__27542));
    Sp12to4 I__6282 (
            .O(N__27572),
            .I(N__27529));
    LocalMux I__6281 (
            .O(N__27569),
            .I(N__27529));
    Sp12to4 I__6280 (
            .O(N__27566),
            .I(N__27529));
    LocalMux I__6279 (
            .O(N__27563),
            .I(N__27529));
    LocalMux I__6278 (
            .O(N__27558),
            .I(N__27529));
    LocalMux I__6277 (
            .O(N__27555),
            .I(N__27529));
    InMux I__6276 (
            .O(N__27554),
            .I(N__27526));
    Span4Mux_v I__6275 (
            .O(N__27545),
            .I(N__27523));
    LocalMux I__6274 (
            .O(N__27542),
            .I(N__27518));
    Span12Mux_v I__6273 (
            .O(N__27529),
            .I(N__27518));
    LocalMux I__6272 (
            .O(N__27526),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__6271 (
            .O(N__27523),
            .I(M_this_state_qZ0Z_4));
    Odrv12 I__6270 (
            .O(N__27518),
            .I(M_this_state_qZ0Z_4));
    CascadeMux I__6269 (
            .O(N__27511),
            .I(N__27508));
    InMux I__6268 (
            .O(N__27508),
            .I(N__27505));
    LocalMux I__6267 (
            .O(N__27505),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_8 ));
    InMux I__6266 (
            .O(N__27502),
            .I(N__27498));
    CascadeMux I__6265 (
            .O(N__27501),
            .I(N__27490));
    LocalMux I__6264 (
            .O(N__27498),
            .I(N__27486));
    InMux I__6263 (
            .O(N__27497),
            .I(N__27483));
    InMux I__6262 (
            .O(N__27496),
            .I(N__27477));
    InMux I__6261 (
            .O(N__27495),
            .I(N__27474));
    InMux I__6260 (
            .O(N__27494),
            .I(N__27471));
    IoInMux I__6259 (
            .O(N__27493),
            .I(N__27468));
    InMux I__6258 (
            .O(N__27490),
            .I(N__27465));
    InMux I__6257 (
            .O(N__27489),
            .I(N__27462));
    Span4Mux_v I__6256 (
            .O(N__27486),
            .I(N__27454));
    LocalMux I__6255 (
            .O(N__27483),
            .I(N__27454));
    InMux I__6254 (
            .O(N__27482),
            .I(N__27445));
    InMux I__6253 (
            .O(N__27481),
            .I(N__27445));
    InMux I__6252 (
            .O(N__27480),
            .I(N__27442));
    LocalMux I__6251 (
            .O(N__27477),
            .I(N__27437));
    LocalMux I__6250 (
            .O(N__27474),
            .I(N__27437));
    LocalMux I__6249 (
            .O(N__27471),
            .I(N__27434));
    LocalMux I__6248 (
            .O(N__27468),
            .I(N__27431));
    LocalMux I__6247 (
            .O(N__27465),
            .I(N__27426));
    LocalMux I__6246 (
            .O(N__27462),
            .I(N__27426));
    InMux I__6245 (
            .O(N__27461),
            .I(N__27419));
    InMux I__6244 (
            .O(N__27460),
            .I(N__27419));
    InMux I__6243 (
            .O(N__27459),
            .I(N__27419));
    Sp12to4 I__6242 (
            .O(N__27454),
            .I(N__27416));
    InMux I__6241 (
            .O(N__27453),
            .I(N__27409));
    InMux I__6240 (
            .O(N__27452),
            .I(N__27409));
    InMux I__6239 (
            .O(N__27451),
            .I(N__27409));
    InMux I__6238 (
            .O(N__27450),
            .I(N__27406));
    LocalMux I__6237 (
            .O(N__27445),
            .I(N__27403));
    LocalMux I__6236 (
            .O(N__27442),
            .I(N__27400));
    Span4Mux_v I__6235 (
            .O(N__27437),
            .I(N__27397));
    Span4Mux_v I__6234 (
            .O(N__27434),
            .I(N__27394));
    IoSpan4Mux I__6233 (
            .O(N__27431),
            .I(N__27391));
    Span12Mux_v I__6232 (
            .O(N__27426),
            .I(N__27388));
    LocalMux I__6231 (
            .O(N__27419),
            .I(N__27383));
    Span12Mux_s9_h I__6230 (
            .O(N__27416),
            .I(N__27383));
    LocalMux I__6229 (
            .O(N__27409),
            .I(N__27374));
    LocalMux I__6228 (
            .O(N__27406),
            .I(N__27374));
    Sp12to4 I__6227 (
            .O(N__27403),
            .I(N__27374));
    Sp12to4 I__6226 (
            .O(N__27400),
            .I(N__27374));
    Span4Mux_h I__6225 (
            .O(N__27397),
            .I(N__27371));
    Span4Mux_h I__6224 (
            .O(N__27394),
            .I(N__27368));
    Span4Mux_s2_h I__6223 (
            .O(N__27391),
            .I(N__27365));
    Span12Mux_h I__6222 (
            .O(N__27388),
            .I(N__27362));
    Span12Mux_h I__6221 (
            .O(N__27383),
            .I(N__27359));
    Span12Mux_v I__6220 (
            .O(N__27374),
            .I(N__27356));
    Span4Mux_h I__6219 (
            .O(N__27371),
            .I(N__27351));
    Span4Mux_v I__6218 (
            .O(N__27368),
            .I(N__27351));
    Span4Mux_h I__6217 (
            .O(N__27365),
            .I(N__27348));
    Odrv12 I__6216 (
            .O(N__27362),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__6215 (
            .O(N__27359),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__6214 (
            .O(N__27356),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__6213 (
            .O(N__27351),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__6212 (
            .O(N__27348),
            .I(M_this_reset_cond_out_0));
    CascadeMux I__6211 (
            .O(N__27337),
            .I(\this_vga_signals.M_this_external_address_d_5Z0Z_13_cascade_ ));
    InMux I__6210 (
            .O(N__27334),
            .I(N__27331));
    LocalMux I__6209 (
            .O(N__27331),
            .I(N__27327));
    CascadeMux I__6208 (
            .O(N__27330),
            .I(N__27324));
    Span4Mux_h I__6207 (
            .O(N__27327),
            .I(N__27321));
    InMux I__6206 (
            .O(N__27324),
            .I(N__27318));
    Odrv4 I__6205 (
            .O(N__27321),
            .I(\this_vga_signals.M_this_state_d_1_sqmuxaZ0 ));
    LocalMux I__6204 (
            .O(N__27318),
            .I(\this_vga_signals.M_this_state_d_1_sqmuxaZ0 ));
    CascadeMux I__6203 (
            .O(N__27313),
            .I(N__27310));
    InMux I__6202 (
            .O(N__27310),
            .I(N__27304));
    InMux I__6201 (
            .O(N__27309),
            .I(N__27304));
    LocalMux I__6200 (
            .O(N__27304),
            .I(\this_vga_signals.M_this_state_d_0_sqmuxaZ0Z_1 ));
    CascadeMux I__6199 (
            .O(N__27301),
            .I(\this_vga_signals.un1_M_this_state_q_21_0_cascade_ ));
    InMux I__6198 (
            .O(N__27298),
            .I(N__27295));
    LocalMux I__6197 (
            .O(N__27295),
            .I(\this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_13 ));
    SRMux I__6196 (
            .O(N__27292),
            .I(N__27256));
    SRMux I__6195 (
            .O(N__27291),
            .I(N__27256));
    SRMux I__6194 (
            .O(N__27290),
            .I(N__27256));
    SRMux I__6193 (
            .O(N__27289),
            .I(N__27256));
    SRMux I__6192 (
            .O(N__27288),
            .I(N__27256));
    SRMux I__6191 (
            .O(N__27287),
            .I(N__27256));
    SRMux I__6190 (
            .O(N__27286),
            .I(N__27256));
    SRMux I__6189 (
            .O(N__27285),
            .I(N__27256));
    SRMux I__6188 (
            .O(N__27284),
            .I(N__27256));
    SRMux I__6187 (
            .O(N__27283),
            .I(N__27256));
    SRMux I__6186 (
            .O(N__27282),
            .I(N__27256));
    SRMux I__6185 (
            .O(N__27281),
            .I(N__27256));
    GlobalMux I__6184 (
            .O(N__27256),
            .I(N__27253));
    gio2CtrlBuf I__6183 (
            .O(N__27253),
            .I(N_989_g));
    InMux I__6182 (
            .O(N__27250),
            .I(N__27247));
    LocalMux I__6181 (
            .O(N__27247),
            .I(N__27243));
    InMux I__6180 (
            .O(N__27246),
            .I(N__27240));
    Odrv4 I__6179 (
            .O(N__27243),
            .I(\this_vga_signals.N_469 ));
    LocalMux I__6178 (
            .O(N__27240),
            .I(\this_vga_signals.N_469 ));
    InMux I__6177 (
            .O(N__27235),
            .I(N__27232));
    LocalMux I__6176 (
            .O(N__27232),
            .I(N__27228));
    InMux I__6175 (
            .O(N__27231),
            .I(N__27223));
    Span4Mux_v I__6174 (
            .O(N__27228),
            .I(N__27220));
    CascadeMux I__6173 (
            .O(N__27227),
            .I(N__27217));
    InMux I__6172 (
            .O(N__27226),
            .I(N__27212));
    LocalMux I__6171 (
            .O(N__27223),
            .I(N__27209));
    Span4Mux_h I__6170 (
            .O(N__27220),
            .I(N__27203));
    InMux I__6169 (
            .O(N__27217),
            .I(N__27200));
    InMux I__6168 (
            .O(N__27216),
            .I(N__27195));
    InMux I__6167 (
            .O(N__27215),
            .I(N__27195));
    LocalMux I__6166 (
            .O(N__27212),
            .I(N__27190));
    Span4Mux_h I__6165 (
            .O(N__27209),
            .I(N__27190));
    InMux I__6164 (
            .O(N__27208),
            .I(N__27185));
    InMux I__6163 (
            .O(N__27207),
            .I(N__27185));
    InMux I__6162 (
            .O(N__27206),
            .I(N__27182));
    Odrv4 I__6161 (
            .O(N__27203),
            .I(M_this_state_qZ0Z_14));
    LocalMux I__6160 (
            .O(N__27200),
            .I(M_this_state_qZ0Z_14));
    LocalMux I__6159 (
            .O(N__27195),
            .I(M_this_state_qZ0Z_14));
    Odrv4 I__6158 (
            .O(N__27190),
            .I(M_this_state_qZ0Z_14));
    LocalMux I__6157 (
            .O(N__27185),
            .I(M_this_state_qZ0Z_14));
    LocalMux I__6156 (
            .O(N__27182),
            .I(M_this_state_qZ0Z_14));
    InMux I__6155 (
            .O(N__27169),
            .I(N__27162));
    InMux I__6154 (
            .O(N__27168),
            .I(N__27162));
    InMux I__6153 (
            .O(N__27167),
            .I(N__27155));
    LocalMux I__6152 (
            .O(N__27162),
            .I(N__27152));
    InMux I__6151 (
            .O(N__27161),
            .I(N__27149));
    InMux I__6150 (
            .O(N__27160),
            .I(N__27146));
    InMux I__6149 (
            .O(N__27159),
            .I(N__27143));
    InMux I__6148 (
            .O(N__27158),
            .I(N__27140));
    LocalMux I__6147 (
            .O(N__27155),
            .I(this_start_data_delay_M_last_q));
    Odrv12 I__6146 (
            .O(N__27152),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__6145 (
            .O(N__27149),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__6144 (
            .O(N__27146),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__6143 (
            .O(N__27143),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__6142 (
            .O(N__27140),
            .I(this_start_data_delay_M_last_q));
    CascadeMux I__6141 (
            .O(N__27127),
            .I(N__27123));
    CascadeMux I__6140 (
            .O(N__27126),
            .I(N__27120));
    InMux I__6139 (
            .O(N__27123),
            .I(N__27115));
    InMux I__6138 (
            .O(N__27120),
            .I(N__27112));
    InMux I__6137 (
            .O(N__27119),
            .I(N__27107));
    InMux I__6136 (
            .O(N__27118),
            .I(N__27107));
    LocalMux I__6135 (
            .O(N__27115),
            .I(N__27104));
    LocalMux I__6134 (
            .O(N__27112),
            .I(N__27099));
    LocalMux I__6133 (
            .O(N__27107),
            .I(N__27099));
    Span4Mux_v I__6132 (
            .O(N__27104),
            .I(N__27093));
    Span4Mux_v I__6131 (
            .O(N__27099),
            .I(N__27090));
    CascadeMux I__6130 (
            .O(N__27098),
            .I(N__27087));
    CascadeMux I__6129 (
            .O(N__27097),
            .I(N__27083));
    CascadeMux I__6128 (
            .O(N__27096),
            .I(N__27080));
    Span4Mux_h I__6127 (
            .O(N__27093),
            .I(N__27075));
    Span4Mux_h I__6126 (
            .O(N__27090),
            .I(N__27075));
    InMux I__6125 (
            .O(N__27087),
            .I(N__27070));
    InMux I__6124 (
            .O(N__27086),
            .I(N__27070));
    InMux I__6123 (
            .O(N__27083),
            .I(N__27065));
    InMux I__6122 (
            .O(N__27080),
            .I(N__27065));
    Sp12to4 I__6121 (
            .O(N__27075),
            .I(N__27058));
    LocalMux I__6120 (
            .O(N__27070),
            .I(N__27058));
    LocalMux I__6119 (
            .O(N__27065),
            .I(N__27058));
    Span12Mux_h I__6118 (
            .O(N__27058),
            .I(N__27055));
    Odrv12 I__6117 (
            .O(N__27055),
            .I(port_enb_c));
    InMux I__6116 (
            .O(N__27052),
            .I(N__27046));
    InMux I__6115 (
            .O(N__27051),
            .I(N__27046));
    LocalMux I__6114 (
            .O(N__27046),
            .I(N__27039));
    InMux I__6113 (
            .O(N__27045),
            .I(N__27036));
    InMux I__6112 (
            .O(N__27044),
            .I(N__27031));
    InMux I__6111 (
            .O(N__27043),
            .I(N__27031));
    InMux I__6110 (
            .O(N__27042),
            .I(N__27026));
    Span4Mux_h I__6109 (
            .O(N__27039),
            .I(N__27023));
    LocalMux I__6108 (
            .O(N__27036),
            .I(N__27018));
    LocalMux I__6107 (
            .O(N__27031),
            .I(N__27018));
    InMux I__6106 (
            .O(N__27030),
            .I(N__27013));
    InMux I__6105 (
            .O(N__27029),
            .I(N__27013));
    LocalMux I__6104 (
            .O(N__27026),
            .I(M_this_delay_clk_out_0));
    Odrv4 I__6103 (
            .O(N__27023),
            .I(M_this_delay_clk_out_0));
    Odrv4 I__6102 (
            .O(N__27018),
            .I(M_this_delay_clk_out_0));
    LocalMux I__6101 (
            .O(N__27013),
            .I(M_this_delay_clk_out_0));
    InMux I__6100 (
            .O(N__27004),
            .I(N__26999));
    InMux I__6099 (
            .O(N__27003),
            .I(N__26996));
    CascadeMux I__6098 (
            .O(N__27002),
            .I(N__26992));
    LocalMux I__6097 (
            .O(N__26999),
            .I(N__26988));
    LocalMux I__6096 (
            .O(N__26996),
            .I(N__26985));
    CascadeMux I__6095 (
            .O(N__26995),
            .I(N__26982));
    InMux I__6094 (
            .O(N__26992),
            .I(N__26979));
    CascadeMux I__6093 (
            .O(N__26991),
            .I(N__26975));
    Span4Mux_v I__6092 (
            .O(N__26988),
            .I(N__26969));
    Span4Mux_v I__6091 (
            .O(N__26985),
            .I(N__26969));
    InMux I__6090 (
            .O(N__26982),
            .I(N__26966));
    LocalMux I__6089 (
            .O(N__26979),
            .I(N__26963));
    InMux I__6088 (
            .O(N__26978),
            .I(N__26960));
    InMux I__6087 (
            .O(N__26975),
            .I(N__26957));
    InMux I__6086 (
            .O(N__26974),
            .I(N__26954));
    Span4Mux_h I__6085 (
            .O(N__26969),
            .I(N__26948));
    LocalMux I__6084 (
            .O(N__26966),
            .I(N__26948));
    Span4Mux_v I__6083 (
            .O(N__26963),
            .I(N__26944));
    LocalMux I__6082 (
            .O(N__26960),
            .I(N__26937));
    LocalMux I__6081 (
            .O(N__26957),
            .I(N__26937));
    LocalMux I__6080 (
            .O(N__26954),
            .I(N__26937));
    InMux I__6079 (
            .O(N__26953),
            .I(N__26934));
    Span4Mux_v I__6078 (
            .O(N__26948),
            .I(N__26931));
    InMux I__6077 (
            .O(N__26947),
            .I(N__26928));
    Span4Mux_h I__6076 (
            .O(N__26944),
            .I(N__26921));
    Span4Mux_v I__6075 (
            .O(N__26937),
            .I(N__26921));
    LocalMux I__6074 (
            .O(N__26934),
            .I(N__26921));
    Sp12to4 I__6073 (
            .O(N__26931),
            .I(N__26918));
    LocalMux I__6072 (
            .O(N__26928),
            .I(N__26915));
    Span4Mux_v I__6071 (
            .O(N__26921),
            .I(N__26912));
    Span12Mux_s10_h I__6070 (
            .O(N__26918),
            .I(N__26909));
    Sp12to4 I__6069 (
            .O(N__26915),
            .I(N__26906));
    Sp12to4 I__6068 (
            .O(N__26912),
            .I(N__26903));
    Span12Mux_v I__6067 (
            .O(N__26909),
            .I(N__26900));
    Span12Mux_v I__6066 (
            .O(N__26906),
            .I(N__26895));
    Span12Mux_h I__6065 (
            .O(N__26903),
            .I(N__26895));
    Odrv12 I__6064 (
            .O(N__26900),
            .I(port_address_in_2));
    Odrv12 I__6063 (
            .O(N__26895),
            .I(port_address_in_2));
    InMux I__6062 (
            .O(N__26890),
            .I(N__26886));
    CascadeMux I__6061 (
            .O(N__26889),
            .I(N__26883));
    LocalMux I__6060 (
            .O(N__26886),
            .I(N__26879));
    InMux I__6059 (
            .O(N__26883),
            .I(N__26874));
    InMux I__6058 (
            .O(N__26882),
            .I(N__26870));
    Span4Mux_v I__6057 (
            .O(N__26879),
            .I(N__26867));
    InMux I__6056 (
            .O(N__26878),
            .I(N__26864));
    CascadeMux I__6055 (
            .O(N__26877),
            .I(N__26860));
    LocalMux I__6054 (
            .O(N__26874),
            .I(N__26857));
    InMux I__6053 (
            .O(N__26873),
            .I(N__26853));
    LocalMux I__6052 (
            .O(N__26870),
            .I(N__26846));
    Sp12to4 I__6051 (
            .O(N__26867),
            .I(N__26846));
    LocalMux I__6050 (
            .O(N__26864),
            .I(N__26846));
    InMux I__6049 (
            .O(N__26863),
            .I(N__26843));
    InMux I__6048 (
            .O(N__26860),
            .I(N__26840));
    Span4Mux_v I__6047 (
            .O(N__26857),
            .I(N__26837));
    InMux I__6046 (
            .O(N__26856),
            .I(N__26834));
    LocalMux I__6045 (
            .O(N__26853),
            .I(N__26831));
    Span12Mux_h I__6044 (
            .O(N__26846),
            .I(N__26826));
    LocalMux I__6043 (
            .O(N__26843),
            .I(N__26826));
    LocalMux I__6042 (
            .O(N__26840),
            .I(N__26823));
    Span4Mux_h I__6041 (
            .O(N__26837),
            .I(N__26818));
    LocalMux I__6040 (
            .O(N__26834),
            .I(N__26818));
    Span12Mux_v I__6039 (
            .O(N__26831),
            .I(N__26815));
    Span12Mux_v I__6038 (
            .O(N__26826),
            .I(N__26812));
    Span12Mux_v I__6037 (
            .O(N__26823),
            .I(N__26807));
    Sp12to4 I__6036 (
            .O(N__26818),
            .I(N__26807));
    Odrv12 I__6035 (
            .O(N__26815),
            .I(port_address_in_0));
    Odrv12 I__6034 (
            .O(N__26812),
            .I(port_address_in_0));
    Odrv12 I__6033 (
            .O(N__26807),
            .I(port_address_in_0));
    CascadeMux I__6032 (
            .O(N__26800),
            .I(N__26797));
    InMux I__6031 (
            .O(N__26797),
            .I(N__26793));
    CascadeMux I__6030 (
            .O(N__26796),
            .I(N__26787));
    LocalMux I__6029 (
            .O(N__26793),
            .I(N__26783));
    InMux I__6028 (
            .O(N__26792),
            .I(N__26776));
    InMux I__6027 (
            .O(N__26791),
            .I(N__26776));
    InMux I__6026 (
            .O(N__26790),
            .I(N__26776));
    InMux I__6025 (
            .O(N__26787),
            .I(N__26773));
    InMux I__6024 (
            .O(N__26786),
            .I(N__26770));
    Span4Mux_v I__6023 (
            .O(N__26783),
            .I(N__26766));
    LocalMux I__6022 (
            .O(N__26776),
            .I(N__26759));
    LocalMux I__6021 (
            .O(N__26773),
            .I(N__26759));
    LocalMux I__6020 (
            .O(N__26770),
            .I(N__26759));
    InMux I__6019 (
            .O(N__26769),
            .I(N__26756));
    Sp12to4 I__6018 (
            .O(N__26766),
            .I(N__26753));
    Sp12to4 I__6017 (
            .O(N__26759),
            .I(N__26748));
    LocalMux I__6016 (
            .O(N__26756),
            .I(N__26748));
    Span12Mux_h I__6015 (
            .O(N__26753),
            .I(N__26745));
    Span12Mux_v I__6014 (
            .O(N__26748),
            .I(N__26742));
    Span12Mux_v I__6013 (
            .O(N__26745),
            .I(N__26737));
    Span12Mux_h I__6012 (
            .O(N__26742),
            .I(N__26737));
    Odrv12 I__6011 (
            .O(N__26737),
            .I(port_address_in_3));
    InMux I__6010 (
            .O(N__26734),
            .I(N__26725));
    InMux I__6009 (
            .O(N__26733),
            .I(N__26725));
    InMux I__6008 (
            .O(N__26732),
            .I(N__26725));
    LocalMux I__6007 (
            .O(N__26725),
            .I(N__26721));
    InMux I__6006 (
            .O(N__26724),
            .I(N__26718));
    Span4Mux_h I__6005 (
            .O(N__26721),
            .I(N__26710));
    LocalMux I__6004 (
            .O(N__26718),
            .I(N__26710));
    InMux I__6003 (
            .O(N__26717),
            .I(N__26707));
    InMux I__6002 (
            .O(N__26716),
            .I(N__26704));
    InMux I__6001 (
            .O(N__26715),
            .I(N__26701));
    Span4Mux_h I__6000 (
            .O(N__26710),
            .I(N__26696));
    LocalMux I__5999 (
            .O(N__26707),
            .I(N__26696));
    LocalMux I__5998 (
            .O(N__26704),
            .I(N__26691));
    LocalMux I__5997 (
            .O(N__26701),
            .I(N__26691));
    Span4Mux_v I__5996 (
            .O(N__26696),
            .I(N__26688));
    Span4Mux_v I__5995 (
            .O(N__26691),
            .I(N__26685));
    Sp12to4 I__5994 (
            .O(N__26688),
            .I(N__26680));
    Sp12to4 I__5993 (
            .O(N__26685),
            .I(N__26680));
    Span12Mux_h I__5992 (
            .O(N__26680),
            .I(N__26677));
    Odrv12 I__5991 (
            .O(N__26677),
            .I(port_address_in_1));
    CascadeMux I__5990 (
            .O(N__26674),
            .I(N__26671));
    InMux I__5989 (
            .O(N__26671),
            .I(N__26668));
    LocalMux I__5988 (
            .O(N__26668),
            .I(N__26665));
    Odrv4 I__5987 (
            .O(N__26665),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_10 ));
    InMux I__5986 (
            .O(N__26662),
            .I(N__26659));
    LocalMux I__5985 (
            .O(N__26659),
            .I(\this_vga_signals.M_this_map_address_d_8_mZ0Z_1 ));
    CascadeMux I__5984 (
            .O(N__26656),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_1_cascade_ ));
    InMux I__5983 (
            .O(N__26653),
            .I(N__26650));
    LocalMux I__5982 (
            .O(N__26650),
            .I(un1_M_this_map_address_q_cry_0_c_RNI6GRRZ0));
    CascadeMux I__5981 (
            .O(N__26647),
            .I(N__26644));
    CascadeBuf I__5980 (
            .O(N__26644),
            .I(N__26641));
    CascadeMux I__5979 (
            .O(N__26641),
            .I(N__26638));
    InMux I__5978 (
            .O(N__26638),
            .I(N__26635));
    LocalMux I__5977 (
            .O(N__26635),
            .I(N__26632));
    Span4Mux_v I__5976 (
            .O(N__26632),
            .I(N__26629));
    Span4Mux_h I__5975 (
            .O(N__26629),
            .I(N__26623));
    InMux I__5974 (
            .O(N__26628),
            .I(N__26620));
    InMux I__5973 (
            .O(N__26627),
            .I(N__26617));
    InMux I__5972 (
            .O(N__26626),
            .I(N__26614));
    Span4Mux_v I__5971 (
            .O(N__26623),
            .I(N__26611));
    LocalMux I__5970 (
            .O(N__26620),
            .I(M_this_map_address_qZ0Z_1));
    LocalMux I__5969 (
            .O(N__26617),
            .I(M_this_map_address_qZ0Z_1));
    LocalMux I__5968 (
            .O(N__26614),
            .I(M_this_map_address_qZ0Z_1));
    Odrv4 I__5967 (
            .O(N__26611),
            .I(M_this_map_address_qZ0Z_1));
    CascadeMux I__5966 (
            .O(N__26602),
            .I(\this_vga_signals.M_this_map_address_d_8_mZ0Z_3_cascade_ ));
    InMux I__5965 (
            .O(N__26599),
            .I(N__26596));
    LocalMux I__5964 (
            .O(N__26596),
            .I(un1_M_this_map_address_q_cry_2_c_RNIAMTRZ0));
    CascadeMux I__5963 (
            .O(N__26593),
            .I(N__26590));
    CascadeBuf I__5962 (
            .O(N__26590),
            .I(N__26587));
    CascadeMux I__5961 (
            .O(N__26587),
            .I(N__26584));
    InMux I__5960 (
            .O(N__26584),
            .I(N__26581));
    LocalMux I__5959 (
            .O(N__26581),
            .I(N__26578));
    Span4Mux_s3_v I__5958 (
            .O(N__26578),
            .I(N__26575));
    Span4Mux_h I__5957 (
            .O(N__26575),
            .I(N__26569));
    InMux I__5956 (
            .O(N__26574),
            .I(N__26566));
    InMux I__5955 (
            .O(N__26573),
            .I(N__26563));
    InMux I__5954 (
            .O(N__26572),
            .I(N__26560));
    Span4Mux_v I__5953 (
            .O(N__26569),
            .I(N__26557));
    LocalMux I__5952 (
            .O(N__26566),
            .I(M_this_map_address_qZ0Z_3));
    LocalMux I__5951 (
            .O(N__26563),
            .I(M_this_map_address_qZ0Z_3));
    LocalMux I__5950 (
            .O(N__26560),
            .I(M_this_map_address_qZ0Z_3));
    Odrv4 I__5949 (
            .O(N__26557),
            .I(M_this_map_address_qZ0Z_3));
    InMux I__5948 (
            .O(N__26548),
            .I(N__26545));
    LocalMux I__5947 (
            .O(N__26545),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_3 ));
    InMux I__5946 (
            .O(N__26542),
            .I(N__26539));
    LocalMux I__5945 (
            .O(N__26539),
            .I(\this_vga_signals.M_this_map_address_d_8_mZ0Z_4 ));
    CascadeMux I__5944 (
            .O(N__26536),
            .I(N__26533));
    InMux I__5943 (
            .O(N__26533),
            .I(N__26530));
    LocalMux I__5942 (
            .O(N__26530),
            .I(N__26527));
    Odrv4 I__5941 (
            .O(N__26527),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_4 ));
    InMux I__5940 (
            .O(N__26524),
            .I(N__26521));
    LocalMux I__5939 (
            .O(N__26521),
            .I(un1_M_this_map_address_q_cry_3_c_RNICPURZ0));
    CascadeMux I__5938 (
            .O(N__26518),
            .I(N__26515));
    CascadeBuf I__5937 (
            .O(N__26515),
            .I(N__26512));
    CascadeMux I__5936 (
            .O(N__26512),
            .I(N__26509));
    InMux I__5935 (
            .O(N__26509),
            .I(N__26506));
    LocalMux I__5934 (
            .O(N__26506),
            .I(N__26503));
    Span4Mux_s3_v I__5933 (
            .O(N__26503),
            .I(N__26500));
    Span4Mux_h I__5932 (
            .O(N__26500),
            .I(N__26494));
    InMux I__5931 (
            .O(N__26499),
            .I(N__26489));
    InMux I__5930 (
            .O(N__26498),
            .I(N__26489));
    InMux I__5929 (
            .O(N__26497),
            .I(N__26486));
    Span4Mux_v I__5928 (
            .O(N__26494),
            .I(N__26483));
    LocalMux I__5927 (
            .O(N__26489),
            .I(M_this_map_address_qZ0Z_4));
    LocalMux I__5926 (
            .O(N__26486),
            .I(M_this_map_address_qZ0Z_4));
    Odrv4 I__5925 (
            .O(N__26483),
            .I(M_this_map_address_qZ0Z_4));
    InMux I__5924 (
            .O(N__26476),
            .I(N__26468));
    InMux I__5923 (
            .O(N__26475),
            .I(N__26465));
    InMux I__5922 (
            .O(N__26474),
            .I(N__26459));
    InMux I__5921 (
            .O(N__26473),
            .I(N__26454));
    InMux I__5920 (
            .O(N__26472),
            .I(N__26454));
    InMux I__5919 (
            .O(N__26471),
            .I(N__26450));
    LocalMux I__5918 (
            .O(N__26468),
            .I(N__26445));
    LocalMux I__5917 (
            .O(N__26465),
            .I(N__26445));
    InMux I__5916 (
            .O(N__26464),
            .I(N__26442));
    InMux I__5915 (
            .O(N__26463),
            .I(N__26437));
    InMux I__5914 (
            .O(N__26462),
            .I(N__26437));
    LocalMux I__5913 (
            .O(N__26459),
            .I(N__26433));
    LocalMux I__5912 (
            .O(N__26454),
            .I(N__26430));
    InMux I__5911 (
            .O(N__26453),
            .I(N__26427));
    LocalMux I__5910 (
            .O(N__26450),
            .I(N__26420));
    Span4Mux_h I__5909 (
            .O(N__26445),
            .I(N__26420));
    LocalMux I__5908 (
            .O(N__26442),
            .I(N__26417));
    LocalMux I__5907 (
            .O(N__26437),
            .I(N__26414));
    InMux I__5906 (
            .O(N__26436),
            .I(N__26411));
    Span4Mux_h I__5905 (
            .O(N__26433),
            .I(N__26404));
    Span4Mux_v I__5904 (
            .O(N__26430),
            .I(N__26404));
    LocalMux I__5903 (
            .O(N__26427),
            .I(N__26404));
    InMux I__5902 (
            .O(N__26426),
            .I(N__26401));
    CascadeMux I__5901 (
            .O(N__26425),
            .I(N__26396));
    Span4Mux_v I__5900 (
            .O(N__26420),
            .I(N__26393));
    Span4Mux_v I__5899 (
            .O(N__26417),
            .I(N__26386));
    Span4Mux_h I__5898 (
            .O(N__26414),
            .I(N__26386));
    LocalMux I__5897 (
            .O(N__26411),
            .I(N__26386));
    Span4Mux_v I__5896 (
            .O(N__26404),
            .I(N__26381));
    LocalMux I__5895 (
            .O(N__26401),
            .I(N__26381));
    InMux I__5894 (
            .O(N__26400),
            .I(N__26378));
    InMux I__5893 (
            .O(N__26399),
            .I(N__26373));
    InMux I__5892 (
            .O(N__26396),
            .I(N__26373));
    Odrv4 I__5891 (
            .O(N__26393),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__5890 (
            .O(N__26386),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__5889 (
            .O(N__26381),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__5888 (
            .O(N__26378),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__5887 (
            .O(N__26373),
            .I(M_this_state_qZ0Z_3));
    CascadeMux I__5886 (
            .O(N__26362),
            .I(N__26357));
    InMux I__5885 (
            .O(N__26361),
            .I(N__26354));
    InMux I__5884 (
            .O(N__26360),
            .I(N__26351));
    InMux I__5883 (
            .O(N__26357),
            .I(N__26348));
    LocalMux I__5882 (
            .O(N__26354),
            .I(N__26345));
    LocalMux I__5881 (
            .O(N__26351),
            .I(N__26340));
    LocalMux I__5880 (
            .O(N__26348),
            .I(N__26340));
    Odrv4 I__5879 (
            .O(N__26345),
            .I(un1_M_this_state_q_12_0));
    Odrv4 I__5878 (
            .O(N__26340),
            .I(un1_M_this_state_q_12_0));
    InMux I__5877 (
            .O(N__26335),
            .I(N__26332));
    LocalMux I__5876 (
            .O(N__26332),
            .I(\this_vga_signals.M_this_map_address_d_5_mZ0Z_8 ));
    InMux I__5875 (
            .O(N__26329),
            .I(N__26317));
    InMux I__5874 (
            .O(N__26328),
            .I(N__26317));
    InMux I__5873 (
            .O(N__26327),
            .I(N__26317));
    InMux I__5872 (
            .O(N__26326),
            .I(N__26310));
    InMux I__5871 (
            .O(N__26325),
            .I(N__26310));
    InMux I__5870 (
            .O(N__26324),
            .I(N__26310));
    LocalMux I__5869 (
            .O(N__26317),
            .I(N__26303));
    LocalMux I__5868 (
            .O(N__26310),
            .I(N__26300));
    InMux I__5867 (
            .O(N__26309),
            .I(N__26297));
    InMux I__5866 (
            .O(N__26308),
            .I(N__26290));
    InMux I__5865 (
            .O(N__26307),
            .I(N__26290));
    InMux I__5864 (
            .O(N__26306),
            .I(N__26290));
    Odrv4 I__5863 (
            .O(N__26303),
            .I(\this_vga_signals.un1_M_this_map_ram_write_en_0 ));
    Odrv4 I__5862 (
            .O(N__26300),
            .I(\this_vga_signals.un1_M_this_map_ram_write_en_0 ));
    LocalMux I__5861 (
            .O(N__26297),
            .I(\this_vga_signals.un1_M_this_map_ram_write_en_0 ));
    LocalMux I__5860 (
            .O(N__26290),
            .I(\this_vga_signals.un1_M_this_map_ram_write_en_0 ));
    InMux I__5859 (
            .O(N__26281),
            .I(N__26278));
    LocalMux I__5858 (
            .O(N__26278),
            .I(un1_M_this_map_address_q_cry_7_c_RNIK53SZ0));
    InMux I__5857 (
            .O(N__26275),
            .I(N__26272));
    LocalMux I__5856 (
            .O(N__26272),
            .I(\this_vga_signals.M_this_external_address_d_5Z0Z_14 ));
    InMux I__5855 (
            .O(N__26269),
            .I(N__26266));
    LocalMux I__5854 (
            .O(N__26266),
            .I(\this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_14 ));
    CascadeMux I__5853 (
            .O(N__26263),
            .I(N__26260));
    CascadeBuf I__5852 (
            .O(N__26260),
            .I(N__26257));
    CascadeMux I__5851 (
            .O(N__26257),
            .I(N__26254));
    CascadeBuf I__5850 (
            .O(N__26254),
            .I(N__26251));
    CascadeMux I__5849 (
            .O(N__26251),
            .I(N__26248));
    CascadeBuf I__5848 (
            .O(N__26248),
            .I(N__26245));
    CascadeMux I__5847 (
            .O(N__26245),
            .I(N__26242));
    CascadeBuf I__5846 (
            .O(N__26242),
            .I(N__26239));
    CascadeMux I__5845 (
            .O(N__26239),
            .I(N__26236));
    CascadeBuf I__5844 (
            .O(N__26236),
            .I(N__26233));
    CascadeMux I__5843 (
            .O(N__26233),
            .I(N__26230));
    CascadeBuf I__5842 (
            .O(N__26230),
            .I(N__26227));
    CascadeMux I__5841 (
            .O(N__26227),
            .I(N__26224));
    CascadeBuf I__5840 (
            .O(N__26224),
            .I(N__26221));
    CascadeMux I__5839 (
            .O(N__26221),
            .I(N__26218));
    CascadeBuf I__5838 (
            .O(N__26218),
            .I(N__26215));
    CascadeMux I__5837 (
            .O(N__26215),
            .I(N__26212));
    CascadeBuf I__5836 (
            .O(N__26212),
            .I(N__26209));
    CascadeMux I__5835 (
            .O(N__26209),
            .I(N__26206));
    CascadeBuf I__5834 (
            .O(N__26206),
            .I(N__26203));
    CascadeMux I__5833 (
            .O(N__26203),
            .I(N__26200));
    CascadeBuf I__5832 (
            .O(N__26200),
            .I(N__26197));
    CascadeMux I__5831 (
            .O(N__26197),
            .I(N__26194));
    CascadeBuf I__5830 (
            .O(N__26194),
            .I(N__26191));
    CascadeMux I__5829 (
            .O(N__26191),
            .I(N__26188));
    CascadeBuf I__5828 (
            .O(N__26188),
            .I(N__26185));
    CascadeMux I__5827 (
            .O(N__26185),
            .I(N__26182));
    CascadeBuf I__5826 (
            .O(N__26182),
            .I(N__26179));
    CascadeMux I__5825 (
            .O(N__26179),
            .I(N__26176));
    CascadeBuf I__5824 (
            .O(N__26176),
            .I(N__26173));
    CascadeMux I__5823 (
            .O(N__26173),
            .I(N__26170));
    InMux I__5822 (
            .O(N__26170),
            .I(N__26167));
    LocalMux I__5821 (
            .O(N__26167),
            .I(N__26162));
    CascadeMux I__5820 (
            .O(N__26166),
            .I(N__26159));
    InMux I__5819 (
            .O(N__26165),
            .I(N__26156));
    Span4Mux_s1_v I__5818 (
            .O(N__26162),
            .I(N__26153));
    InMux I__5817 (
            .O(N__26159),
            .I(N__26149));
    LocalMux I__5816 (
            .O(N__26156),
            .I(N__26146));
    Sp12to4 I__5815 (
            .O(N__26153),
            .I(N__26143));
    InMux I__5814 (
            .O(N__26152),
            .I(N__26140));
    LocalMux I__5813 (
            .O(N__26149),
            .I(N__26135));
    Span4Mux_h I__5812 (
            .O(N__26146),
            .I(N__26135));
    Span12Mux_v I__5811 (
            .O(N__26143),
            .I(N__26132));
    LocalMux I__5810 (
            .O(N__26140),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv4 I__5809 (
            .O(N__26135),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv12 I__5808 (
            .O(N__26132),
            .I(M_this_sprites_address_qZ0Z_4));
    InMux I__5807 (
            .O(N__26125),
            .I(N__26122));
    LocalMux I__5806 (
            .O(N__26122),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4 ));
    CascadeMux I__5805 (
            .O(N__26119),
            .I(N__26116));
    CascadeBuf I__5804 (
            .O(N__26116),
            .I(N__26113));
    CascadeMux I__5803 (
            .O(N__26113),
            .I(N__26110));
    InMux I__5802 (
            .O(N__26110),
            .I(N__26107));
    LocalMux I__5801 (
            .O(N__26107),
            .I(N__26104));
    Span4Mux_h I__5800 (
            .O(N__26104),
            .I(N__26101));
    Span4Mux_h I__5799 (
            .O(N__26101),
            .I(N__26097));
    InMux I__5798 (
            .O(N__26100),
            .I(N__26093));
    Span4Mux_v I__5797 (
            .O(N__26097),
            .I(N__26089));
    InMux I__5796 (
            .O(N__26096),
            .I(N__26086));
    LocalMux I__5795 (
            .O(N__26093),
            .I(N__26083));
    InMux I__5794 (
            .O(N__26092),
            .I(N__26080));
    Span4Mux_v I__5793 (
            .O(N__26089),
            .I(N__26077));
    LocalMux I__5792 (
            .O(N__26086),
            .I(M_this_map_address_qZ0Z_0));
    Odrv4 I__5791 (
            .O(N__26083),
            .I(M_this_map_address_qZ0Z_0));
    LocalMux I__5790 (
            .O(N__26080),
            .I(M_this_map_address_qZ0Z_0));
    Odrv4 I__5789 (
            .O(N__26077),
            .I(M_this_map_address_qZ0Z_0));
    InMux I__5788 (
            .O(N__26068),
            .I(N__26065));
    LocalMux I__5787 (
            .O(N__26065),
            .I(\this_vga_signals.M_this_map_address_d_8_mZ0Z_0 ));
    CascadeMux I__5786 (
            .O(N__26062),
            .I(N__26059));
    CascadeBuf I__5785 (
            .O(N__26059),
            .I(N__26056));
    CascadeMux I__5784 (
            .O(N__26056),
            .I(N__26053));
    CascadeBuf I__5783 (
            .O(N__26053),
            .I(N__26050));
    CascadeMux I__5782 (
            .O(N__26050),
            .I(N__26047));
    CascadeBuf I__5781 (
            .O(N__26047),
            .I(N__26044));
    CascadeMux I__5780 (
            .O(N__26044),
            .I(N__26041));
    CascadeBuf I__5779 (
            .O(N__26041),
            .I(N__26038));
    CascadeMux I__5778 (
            .O(N__26038),
            .I(N__26035));
    CascadeBuf I__5777 (
            .O(N__26035),
            .I(N__26032));
    CascadeMux I__5776 (
            .O(N__26032),
            .I(N__26029));
    CascadeBuf I__5775 (
            .O(N__26029),
            .I(N__26026));
    CascadeMux I__5774 (
            .O(N__26026),
            .I(N__26023));
    CascadeBuf I__5773 (
            .O(N__26023),
            .I(N__26020));
    CascadeMux I__5772 (
            .O(N__26020),
            .I(N__26017));
    CascadeBuf I__5771 (
            .O(N__26017),
            .I(N__26014));
    CascadeMux I__5770 (
            .O(N__26014),
            .I(N__26011));
    CascadeBuf I__5769 (
            .O(N__26011),
            .I(N__26008));
    CascadeMux I__5768 (
            .O(N__26008),
            .I(N__26005));
    CascadeBuf I__5767 (
            .O(N__26005),
            .I(N__26002));
    CascadeMux I__5766 (
            .O(N__26002),
            .I(N__25999));
    CascadeBuf I__5765 (
            .O(N__25999),
            .I(N__25996));
    CascadeMux I__5764 (
            .O(N__25996),
            .I(N__25993));
    CascadeBuf I__5763 (
            .O(N__25993),
            .I(N__25990));
    CascadeMux I__5762 (
            .O(N__25990),
            .I(N__25987));
    CascadeBuf I__5761 (
            .O(N__25987),
            .I(N__25984));
    CascadeMux I__5760 (
            .O(N__25984),
            .I(N__25981));
    CascadeBuf I__5759 (
            .O(N__25981),
            .I(N__25978));
    CascadeMux I__5758 (
            .O(N__25978),
            .I(N__25975));
    CascadeBuf I__5757 (
            .O(N__25975),
            .I(N__25972));
    CascadeMux I__5756 (
            .O(N__25972),
            .I(N__25969));
    InMux I__5755 (
            .O(N__25969),
            .I(N__25966));
    LocalMux I__5754 (
            .O(N__25966),
            .I(N__25963));
    Span4Mux_s3_v I__5753 (
            .O(N__25963),
            .I(N__25958));
    InMux I__5752 (
            .O(N__25962),
            .I(N__25955));
    InMux I__5751 (
            .O(N__25961),
            .I(N__25952));
    Span4Mux_v I__5750 (
            .O(N__25958),
            .I(N__25948));
    LocalMux I__5749 (
            .O(N__25955),
            .I(N__25943));
    LocalMux I__5748 (
            .O(N__25952),
            .I(N__25943));
    InMux I__5747 (
            .O(N__25951),
            .I(N__25940));
    Span4Mux_v I__5746 (
            .O(N__25948),
            .I(N__25937));
    Span4Mux_v I__5745 (
            .O(N__25943),
            .I(N__25934));
    LocalMux I__5744 (
            .O(N__25940),
            .I(N__25929));
    Sp12to4 I__5743 (
            .O(N__25937),
            .I(N__25929));
    Odrv4 I__5742 (
            .O(N__25934),
            .I(M_this_sprites_address_qZ0Z_0));
    Odrv12 I__5741 (
            .O(N__25929),
            .I(M_this_sprites_address_qZ0Z_0));
    InMux I__5740 (
            .O(N__25924),
            .I(N__25921));
    LocalMux I__5739 (
            .O(N__25921),
            .I(N__25918));
    Odrv4 I__5738 (
            .O(N__25918),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0 ));
    InMux I__5737 (
            .O(N__25915),
            .I(N__25912));
    LocalMux I__5736 (
            .O(N__25912),
            .I(N__25909));
    Span4Mux_h I__5735 (
            .O(N__25909),
            .I(N__25906));
    Odrv4 I__5734 (
            .O(N__25906),
            .I(\this_vga_signals.N_291 ));
    CascadeMux I__5733 (
            .O(N__25903),
            .I(N__25899));
    InMux I__5732 (
            .O(N__25902),
            .I(N__25895));
    InMux I__5731 (
            .O(N__25899),
            .I(N__25892));
    InMux I__5730 (
            .O(N__25898),
            .I(N__25889));
    LocalMux I__5729 (
            .O(N__25895),
            .I(\this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1 ));
    LocalMux I__5728 (
            .O(N__25892),
            .I(\this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1 ));
    LocalMux I__5727 (
            .O(N__25889),
            .I(\this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1 ));
    CascadeMux I__5726 (
            .O(N__25882),
            .I(N__25878));
    InMux I__5725 (
            .O(N__25881),
            .I(N__25873));
    InMux I__5724 (
            .O(N__25878),
            .I(N__25866));
    InMux I__5723 (
            .O(N__25877),
            .I(N__25866));
    InMux I__5722 (
            .O(N__25876),
            .I(N__25866));
    LocalMux I__5721 (
            .O(N__25873),
            .I(N__25861));
    LocalMux I__5720 (
            .O(N__25866),
            .I(N__25861));
    Span12Mux_v I__5719 (
            .O(N__25861),
            .I(N__25858));
    Span12Mux_h I__5718 (
            .O(N__25858),
            .I(N__25855));
    Odrv12 I__5717 (
            .O(N__25855),
            .I(port_address_in_5));
    InMux I__5716 (
            .O(N__25852),
            .I(N__25843));
    InMux I__5715 (
            .O(N__25851),
            .I(N__25843));
    InMux I__5714 (
            .O(N__25850),
            .I(N__25843));
    LocalMux I__5713 (
            .O(N__25843),
            .I(N__25840));
    Span4Mux_v I__5712 (
            .O(N__25840),
            .I(N__25836));
    InMux I__5711 (
            .O(N__25839),
            .I(N__25833));
    Span4Mux_h I__5710 (
            .O(N__25836),
            .I(N__25830));
    LocalMux I__5709 (
            .O(N__25833),
            .I(N__25827));
    Span4Mux_h I__5708 (
            .O(N__25830),
            .I(N__25824));
    Span12Mux_h I__5707 (
            .O(N__25827),
            .I(N__25821));
    Odrv4 I__5706 (
            .O(N__25824),
            .I(port_address_in_6));
    Odrv12 I__5705 (
            .O(N__25821),
            .I(port_address_in_6));
    CascadeMux I__5704 (
            .O(N__25816),
            .I(\this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_4_cascade_ ));
    InMux I__5703 (
            .O(N__25813),
            .I(N__25804));
    InMux I__5702 (
            .O(N__25812),
            .I(N__25804));
    InMux I__5701 (
            .O(N__25811),
            .I(N__25801));
    InMux I__5700 (
            .O(N__25810),
            .I(N__25796));
    InMux I__5699 (
            .O(N__25809),
            .I(N__25796));
    LocalMux I__5698 (
            .O(N__25804),
            .I(\this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0 ));
    LocalMux I__5697 (
            .O(N__25801),
            .I(\this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0 ));
    LocalMux I__5696 (
            .O(N__25796),
            .I(\this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0 ));
    InMux I__5695 (
            .O(N__25789),
            .I(N__25786));
    LocalMux I__5694 (
            .O(N__25786),
            .I(N__25783));
    Span4Mux_v I__5693 (
            .O(N__25783),
            .I(N__25779));
    InMux I__5692 (
            .O(N__25782),
            .I(N__25776));
    Span4Mux_h I__5691 (
            .O(N__25779),
            .I(N__25771));
    LocalMux I__5690 (
            .O(N__25776),
            .I(N__25771));
    Odrv4 I__5689 (
            .O(N__25771),
            .I(\this_vga_signals.N_444_1 ));
    InMux I__5688 (
            .O(N__25768),
            .I(N__25765));
    LocalMux I__5687 (
            .O(N__25765),
            .I(N__25761));
    CascadeMux I__5686 (
            .O(N__25764),
            .I(N__25758));
    Span4Mux_h I__5685 (
            .O(N__25761),
            .I(N__25755));
    InMux I__5684 (
            .O(N__25758),
            .I(N__25752));
    Odrv4 I__5683 (
            .O(N__25755),
            .I(this_vga_signals_M_this_state_q_ns_i_o2_0_14));
    LocalMux I__5682 (
            .O(N__25752),
            .I(this_vga_signals_M_this_state_q_ns_i_o2_0_14));
    InMux I__5681 (
            .O(N__25747),
            .I(N__25743));
    InMux I__5680 (
            .O(N__25746),
            .I(N__25740));
    LocalMux I__5679 (
            .O(N__25743),
            .I(N__25735));
    LocalMux I__5678 (
            .O(N__25740),
            .I(N__25735));
    Odrv4 I__5677 (
            .O(N__25735),
            .I(M_this_state_q_fastZ0Z_14));
    InMux I__5676 (
            .O(N__25732),
            .I(N__25729));
    LocalMux I__5675 (
            .O(N__25729),
            .I(N__25720));
    InMux I__5674 (
            .O(N__25728),
            .I(N__25717));
    InMux I__5673 (
            .O(N__25727),
            .I(N__25709));
    InMux I__5672 (
            .O(N__25726),
            .I(N__25709));
    InMux I__5671 (
            .O(N__25725),
            .I(N__25709));
    CascadeMux I__5670 (
            .O(N__25724),
            .I(N__25705));
    InMux I__5669 (
            .O(N__25723),
            .I(N__25702));
    Span4Mux_v I__5668 (
            .O(N__25720),
            .I(N__25699));
    LocalMux I__5667 (
            .O(N__25717),
            .I(N__25696));
    InMux I__5666 (
            .O(N__25716),
            .I(N__25693));
    LocalMux I__5665 (
            .O(N__25709),
            .I(N__25690));
    InMux I__5664 (
            .O(N__25708),
            .I(N__25687));
    InMux I__5663 (
            .O(N__25705),
            .I(N__25684));
    LocalMux I__5662 (
            .O(N__25702),
            .I(N__25680));
    Sp12to4 I__5661 (
            .O(N__25699),
            .I(N__25673));
    Sp12to4 I__5660 (
            .O(N__25696),
            .I(N__25673));
    LocalMux I__5659 (
            .O(N__25693),
            .I(N__25673));
    Span4Mux_v I__5658 (
            .O(N__25690),
            .I(N__25670));
    LocalMux I__5657 (
            .O(N__25687),
            .I(N__25667));
    LocalMux I__5656 (
            .O(N__25684),
            .I(N__25664));
    CascadeMux I__5655 (
            .O(N__25683),
            .I(N__25660));
    Span12Mux_v I__5654 (
            .O(N__25680),
            .I(N__25655));
    Span12Mux_v I__5653 (
            .O(N__25673),
            .I(N__25655));
    Span4Mux_h I__5652 (
            .O(N__25670),
            .I(N__25648));
    Span4Mux_h I__5651 (
            .O(N__25667),
            .I(N__25648));
    Span4Mux_v I__5650 (
            .O(N__25664),
            .I(N__25648));
    InMux I__5649 (
            .O(N__25663),
            .I(N__25645));
    InMux I__5648 (
            .O(N__25660),
            .I(N__25642));
    Odrv12 I__5647 (
            .O(N__25655),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__5646 (
            .O(N__25648),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__5645 (
            .O(N__25645),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__5644 (
            .O(N__25642),
            .I(M_this_sprites_address_qZ0Z_12));
    CascadeMux I__5643 (
            .O(N__25633),
            .I(N__25630));
    InMux I__5642 (
            .O(N__25630),
            .I(N__25627));
    LocalMux I__5641 (
            .O(N__25627),
            .I(N__25624));
    Span4Mux_v I__5640 (
            .O(N__25624),
            .I(N__25621));
    Odrv4 I__5639 (
            .O(N__25621),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_12 ));
    CascadeMux I__5638 (
            .O(N__25618),
            .I(N__25615));
    CascadeBuf I__5637 (
            .O(N__25615),
            .I(N__25612));
    CascadeMux I__5636 (
            .O(N__25612),
            .I(N__25609));
    CascadeBuf I__5635 (
            .O(N__25609),
            .I(N__25606));
    CascadeMux I__5634 (
            .O(N__25606),
            .I(N__25603));
    CascadeBuf I__5633 (
            .O(N__25603),
            .I(N__25600));
    CascadeMux I__5632 (
            .O(N__25600),
            .I(N__25597));
    CascadeBuf I__5631 (
            .O(N__25597),
            .I(N__25594));
    CascadeMux I__5630 (
            .O(N__25594),
            .I(N__25591));
    CascadeBuf I__5629 (
            .O(N__25591),
            .I(N__25588));
    CascadeMux I__5628 (
            .O(N__25588),
            .I(N__25585));
    CascadeBuf I__5627 (
            .O(N__25585),
            .I(N__25582));
    CascadeMux I__5626 (
            .O(N__25582),
            .I(N__25579));
    CascadeBuf I__5625 (
            .O(N__25579),
            .I(N__25576));
    CascadeMux I__5624 (
            .O(N__25576),
            .I(N__25573));
    CascadeBuf I__5623 (
            .O(N__25573),
            .I(N__25570));
    CascadeMux I__5622 (
            .O(N__25570),
            .I(N__25567));
    CascadeBuf I__5621 (
            .O(N__25567),
            .I(N__25564));
    CascadeMux I__5620 (
            .O(N__25564),
            .I(N__25561));
    CascadeBuf I__5619 (
            .O(N__25561),
            .I(N__25558));
    CascadeMux I__5618 (
            .O(N__25558),
            .I(N__25555));
    CascadeBuf I__5617 (
            .O(N__25555),
            .I(N__25552));
    CascadeMux I__5616 (
            .O(N__25552),
            .I(N__25549));
    CascadeBuf I__5615 (
            .O(N__25549),
            .I(N__25546));
    CascadeMux I__5614 (
            .O(N__25546),
            .I(N__25543));
    CascadeBuf I__5613 (
            .O(N__25543),
            .I(N__25540));
    CascadeMux I__5612 (
            .O(N__25540),
            .I(N__25537));
    CascadeBuf I__5611 (
            .O(N__25537),
            .I(N__25534));
    CascadeMux I__5610 (
            .O(N__25534),
            .I(N__25531));
    CascadeBuf I__5609 (
            .O(N__25531),
            .I(N__25528));
    CascadeMux I__5608 (
            .O(N__25528),
            .I(N__25525));
    InMux I__5607 (
            .O(N__25525),
            .I(N__25522));
    LocalMux I__5606 (
            .O(N__25522),
            .I(N__25519));
    Span4Mux_h I__5605 (
            .O(N__25519),
            .I(N__25515));
    InMux I__5604 (
            .O(N__25518),
            .I(N__25511));
    Sp12to4 I__5603 (
            .O(N__25515),
            .I(N__25508));
    InMux I__5602 (
            .O(N__25514),
            .I(N__25505));
    LocalMux I__5601 (
            .O(N__25511),
            .I(N__25502));
    Span12Mux_s6_v I__5600 (
            .O(N__25508),
            .I(N__25498));
    LocalMux I__5599 (
            .O(N__25505),
            .I(N__25495));
    Span4Mux_v I__5598 (
            .O(N__25502),
            .I(N__25492));
    InMux I__5597 (
            .O(N__25501),
            .I(N__25489));
    Span12Mux_v I__5596 (
            .O(N__25498),
            .I(N__25486));
    Odrv12 I__5595 (
            .O(N__25495),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv4 I__5594 (
            .O(N__25492),
            .I(M_this_sprites_address_qZ0Z_1));
    LocalMux I__5593 (
            .O(N__25489),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv12 I__5592 (
            .O(N__25486),
            .I(M_this_sprites_address_qZ0Z_1));
    CascadeMux I__5591 (
            .O(N__25477),
            .I(N_389_0_cascade_));
    InMux I__5590 (
            .O(N__25474),
            .I(N__25471));
    LocalMux I__5589 (
            .O(N__25471),
            .I(N__25468));
    Span4Mux_h I__5588 (
            .O(N__25468),
            .I(N__25465));
    Odrv4 I__5587 (
            .O(N__25465),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1 ));
    InMux I__5586 (
            .O(N__25462),
            .I(N__25458));
    InMux I__5585 (
            .O(N__25461),
            .I(N__25455));
    LocalMux I__5584 (
            .O(N__25458),
            .I(N__25452));
    LocalMux I__5583 (
            .O(N__25455),
            .I(M_this_state_q_fastZ0Z_15));
    Odrv12 I__5582 (
            .O(N__25452),
            .I(M_this_state_q_fastZ0Z_15));
    CascadeMux I__5581 (
            .O(N__25447),
            .I(N__25442));
    InMux I__5580 (
            .O(N__25446),
            .I(N__25439));
    InMux I__5579 (
            .O(N__25445),
            .I(N__25436));
    InMux I__5578 (
            .O(N__25442),
            .I(N__25433));
    LocalMux I__5577 (
            .O(N__25439),
            .I(N__25428));
    LocalMux I__5576 (
            .O(N__25436),
            .I(N__25428));
    LocalMux I__5575 (
            .O(N__25433),
            .I(N__25425));
    Span4Mux_v I__5574 (
            .O(N__25428),
            .I(N__25420));
    Span4Mux_h I__5573 (
            .O(N__25425),
            .I(N__25417));
    InMux I__5572 (
            .O(N__25424),
            .I(N__25412));
    InMux I__5571 (
            .O(N__25423),
            .I(N__25412));
    Odrv4 I__5570 (
            .O(N__25420),
            .I(N_297));
    Odrv4 I__5569 (
            .O(N__25417),
            .I(N_297));
    LocalMux I__5568 (
            .O(N__25412),
            .I(N_297));
    CascadeMux I__5567 (
            .O(N__25405),
            .I(N__25402));
    InMux I__5566 (
            .O(N__25402),
            .I(N__25399));
    LocalMux I__5565 (
            .O(N__25399),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_9 ));
    InMux I__5564 (
            .O(N__25396),
            .I(N__25393));
    LocalMux I__5563 (
            .O(N__25393),
            .I(N__25387));
    InMux I__5562 (
            .O(N__25392),
            .I(N__25384));
    InMux I__5561 (
            .O(N__25391),
            .I(N__25374));
    InMux I__5560 (
            .O(N__25390),
            .I(N__25374));
    Span4Mux_h I__5559 (
            .O(N__25387),
            .I(N__25369));
    LocalMux I__5558 (
            .O(N__25384),
            .I(N__25369));
    InMux I__5557 (
            .O(N__25383),
            .I(N__25364));
    InMux I__5556 (
            .O(N__25382),
            .I(N__25364));
    CascadeMux I__5555 (
            .O(N__25381),
            .I(N__25361));
    InMux I__5554 (
            .O(N__25380),
            .I(N__25358));
    InMux I__5553 (
            .O(N__25379),
            .I(N__25355));
    LocalMux I__5552 (
            .O(N__25374),
            .I(N__25348));
    Span4Mux_v I__5551 (
            .O(N__25369),
            .I(N__25348));
    LocalMux I__5550 (
            .O(N__25364),
            .I(N__25348));
    InMux I__5549 (
            .O(N__25361),
            .I(N__25345));
    LocalMux I__5548 (
            .O(N__25358),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__5547 (
            .O(N__25355),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__5546 (
            .O(N__25348),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__5545 (
            .O(N__25345),
            .I(M_this_state_qZ0Z_9));
    CascadeMux I__5544 (
            .O(N__25336),
            .I(\this_vga_signals.M_this_state_q_ns_0_a3_sxZ0Z_9_cascade_ ));
    InMux I__5543 (
            .O(N__25333),
            .I(N__25327));
    InMux I__5542 (
            .O(N__25332),
            .I(N__25327));
    LocalMux I__5541 (
            .O(N__25327),
            .I(N__25324));
    Span4Mux_v I__5540 (
            .O(N__25324),
            .I(N__25321));
    Span4Mux_v I__5539 (
            .O(N__25321),
            .I(N__25318));
    Span4Mux_h I__5538 (
            .O(N__25318),
            .I(N__25315));
    Span4Mux_h I__5537 (
            .O(N__25315),
            .I(N__25312));
    Odrv4 I__5536 (
            .O(N__25312),
            .I(port_address_in_4));
    InMux I__5535 (
            .O(N__25309),
            .I(N__25305));
    InMux I__5534 (
            .O(N__25308),
            .I(N__25302));
    LocalMux I__5533 (
            .O(N__25305),
            .I(N__25299));
    LocalMux I__5532 (
            .O(N__25302),
            .I(N__25296));
    Span4Mux_h I__5531 (
            .O(N__25299),
            .I(N__25291));
    Span4Mux_h I__5530 (
            .O(N__25296),
            .I(N__25291));
    Span4Mux_v I__5529 (
            .O(N__25291),
            .I(N__25288));
    Sp12to4 I__5528 (
            .O(N__25288),
            .I(N__25284));
    InMux I__5527 (
            .O(N__25287),
            .I(N__25281));
    Span12Mux_h I__5526 (
            .O(N__25284),
            .I(N__25278));
    LocalMux I__5525 (
            .O(N__25281),
            .I(N__25275));
    Odrv12 I__5524 (
            .O(N__25278),
            .I(port_rw_in));
    Odrv12 I__5523 (
            .O(N__25275),
            .I(port_rw_in));
    CascadeMux I__5522 (
            .O(N__25270),
            .I(N__25266));
    CascadeMux I__5521 (
            .O(N__25269),
            .I(N__25263));
    InMux I__5520 (
            .O(N__25266),
            .I(N__25258));
    InMux I__5519 (
            .O(N__25263),
            .I(N__25258));
    LocalMux I__5518 (
            .O(N__25258),
            .I(N__25255));
    Span12Mux_h I__5517 (
            .O(N__25255),
            .I(N__25252));
    Span12Mux_v I__5516 (
            .O(N__25252),
            .I(N__25249));
    Odrv12 I__5515 (
            .O(N__25249),
            .I(port_address_in_7));
    InMux I__5514 (
            .O(N__25246),
            .I(N__25243));
    LocalMux I__5513 (
            .O(N__25243),
            .I(un1_M_this_map_address_q_cry_6_c_RNII22SZ0));
    InMux I__5512 (
            .O(N__25240),
            .I(un1_M_this_map_address_q_cry_6));
    InMux I__5511 (
            .O(N__25237),
            .I(bfn_19_23_0_));
    CascadeMux I__5510 (
            .O(N__25234),
            .I(N__25231));
    CascadeBuf I__5509 (
            .O(N__25231),
            .I(N__25228));
    CascadeMux I__5508 (
            .O(N__25228),
            .I(N__25225));
    InMux I__5507 (
            .O(N__25225),
            .I(N__25222));
    LocalMux I__5506 (
            .O(N__25222),
            .I(N__25219));
    Span4Mux_h I__5505 (
            .O(N__25219),
            .I(N__25215));
    InMux I__5504 (
            .O(N__25218),
            .I(N__25211));
    Sp12to4 I__5503 (
            .O(N__25215),
            .I(N__25207));
    InMux I__5502 (
            .O(N__25214),
            .I(N__25204));
    LocalMux I__5501 (
            .O(N__25211),
            .I(N__25201));
    InMux I__5500 (
            .O(N__25210),
            .I(N__25198));
    Span12Mux_s9_v I__5499 (
            .O(N__25207),
            .I(N__25195));
    LocalMux I__5498 (
            .O(N__25204),
            .I(M_this_map_address_qZ0Z_9));
    Odrv12 I__5497 (
            .O(N__25201),
            .I(M_this_map_address_qZ0Z_9));
    LocalMux I__5496 (
            .O(N__25198),
            .I(M_this_map_address_qZ0Z_9));
    Odrv12 I__5495 (
            .O(N__25195),
            .I(M_this_map_address_qZ0Z_9));
    InMux I__5494 (
            .O(N__25186),
            .I(un1_M_this_map_address_q_cry_8));
    InMux I__5493 (
            .O(N__25183),
            .I(N__25180));
    LocalMux I__5492 (
            .O(N__25180),
            .I(un1_M_this_map_address_q_cry_8_c_RNIM84SZ0));
    InMux I__5491 (
            .O(N__25177),
            .I(N__25174));
    LocalMux I__5490 (
            .O(N__25174),
            .I(\this_vga_signals.M_this_map_address_d_5_mZ0Z_7 ));
    CascadeMux I__5489 (
            .O(N__25171),
            .I(N__25168));
    CascadeBuf I__5488 (
            .O(N__25168),
            .I(N__25165));
    CascadeMux I__5487 (
            .O(N__25165),
            .I(N__25162));
    InMux I__5486 (
            .O(N__25162),
            .I(N__25158));
    CascadeMux I__5485 (
            .O(N__25161),
            .I(N__25153));
    LocalMux I__5484 (
            .O(N__25158),
            .I(N__25150));
    InMux I__5483 (
            .O(N__25157),
            .I(N__25147));
    InMux I__5482 (
            .O(N__25156),
            .I(N__25144));
    InMux I__5481 (
            .O(N__25153),
            .I(N__25141));
    Span12Mux_s9_v I__5480 (
            .O(N__25150),
            .I(N__25138));
    LocalMux I__5479 (
            .O(N__25147),
            .I(M_this_map_address_qZ0Z_7));
    LocalMux I__5478 (
            .O(N__25144),
            .I(M_this_map_address_qZ0Z_7));
    LocalMux I__5477 (
            .O(N__25141),
            .I(M_this_map_address_qZ0Z_7));
    Odrv12 I__5476 (
            .O(N__25138),
            .I(M_this_map_address_qZ0Z_7));
    CascadeMux I__5475 (
            .O(N__25129),
            .I(N__25126));
    InMux I__5474 (
            .O(N__25126),
            .I(N__25123));
    LocalMux I__5473 (
            .O(N__25123),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_7 ));
    CascadeMux I__5472 (
            .O(N__25120),
            .I(N__25117));
    CascadeBuf I__5471 (
            .O(N__25117),
            .I(N__25113));
    CascadeMux I__5470 (
            .O(N__25116),
            .I(N__25110));
    CascadeMux I__5469 (
            .O(N__25113),
            .I(N__25107));
    InMux I__5468 (
            .O(N__25110),
            .I(N__25104));
    InMux I__5467 (
            .O(N__25107),
            .I(N__25101));
    LocalMux I__5466 (
            .O(N__25104),
            .I(N__25098));
    LocalMux I__5465 (
            .O(N__25101),
            .I(N__25094));
    Span4Mux_h I__5464 (
            .O(N__25098),
            .I(N__25090));
    CascadeMux I__5463 (
            .O(N__25097),
            .I(N__25087));
    Span4Mux_s2_v I__5462 (
            .O(N__25094),
            .I(N__25084));
    CascadeMux I__5461 (
            .O(N__25093),
            .I(N__25081));
    Span4Mux_v I__5460 (
            .O(N__25090),
            .I(N__25077));
    InMux I__5459 (
            .O(N__25087),
            .I(N__25074));
    Span4Mux_h I__5458 (
            .O(N__25084),
            .I(N__25071));
    InMux I__5457 (
            .O(N__25081),
            .I(N__25066));
    InMux I__5456 (
            .O(N__25080),
            .I(N__25066));
    Span4Mux_h I__5455 (
            .O(N__25077),
            .I(N__25063));
    LocalMux I__5454 (
            .O(N__25074),
            .I(N__25058));
    Span4Mux_v I__5453 (
            .O(N__25071),
            .I(N__25058));
    LocalMux I__5452 (
            .O(N__25066),
            .I(M_this_ppu_map_addr_2));
    Odrv4 I__5451 (
            .O(N__25063),
            .I(M_this_ppu_map_addr_2));
    Odrv4 I__5450 (
            .O(N__25058),
            .I(M_this_ppu_map_addr_2));
    InMux I__5449 (
            .O(N__25051),
            .I(N__25046));
    InMux I__5448 (
            .O(N__25050),
            .I(N__25041));
    InMux I__5447 (
            .O(N__25049),
            .I(N__25041));
    LocalMux I__5446 (
            .O(N__25046),
            .I(\this_ppu.un1_M_haddress_q_c5 ));
    LocalMux I__5445 (
            .O(N__25041),
            .I(\this_ppu.un1_M_haddress_q_c5 ));
    SRMux I__5444 (
            .O(N__25036),
            .I(N__25031));
    SRMux I__5443 (
            .O(N__25035),
            .I(N__25027));
    SRMux I__5442 (
            .O(N__25034),
            .I(N__25024));
    LocalMux I__5441 (
            .O(N__25031),
            .I(N__25021));
    SRMux I__5440 (
            .O(N__25030),
            .I(N__25018));
    LocalMux I__5439 (
            .O(N__25027),
            .I(N__25015));
    LocalMux I__5438 (
            .O(N__25024),
            .I(N__25012));
    Span4Mux_v I__5437 (
            .O(N__25021),
            .I(N__25007));
    LocalMux I__5436 (
            .O(N__25018),
            .I(N__25007));
    Span4Mux_h I__5435 (
            .O(N__25015),
            .I(N__25004));
    Span4Mux_h I__5434 (
            .O(N__25012),
            .I(N__25001));
    Span4Mux_v I__5433 (
            .O(N__25007),
            .I(N__24998));
    Odrv4 I__5432 (
            .O(N__25004),
            .I(\this_ppu.M_last_q_RNI21NK5 ));
    Odrv4 I__5431 (
            .O(N__25001),
            .I(\this_ppu.M_last_q_RNI21NK5 ));
    Odrv4 I__5430 (
            .O(N__24998),
            .I(\this_ppu.M_last_q_RNI21NK5 ));
    InMux I__5429 (
            .O(N__24991),
            .I(N__24988));
    LocalMux I__5428 (
            .O(N__24988),
            .I(N__24985));
    Odrv12 I__5427 (
            .O(N__24985),
            .I(\this_reset_cond.M_stage_qZ0Z_6 ));
    InMux I__5426 (
            .O(N__24982),
            .I(N__24979));
    LocalMux I__5425 (
            .O(N__24979),
            .I(N__24976));
    Odrv12 I__5424 (
            .O(N__24976),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    CascadeMux I__5423 (
            .O(N__24973),
            .I(N__24970));
    CascadeBuf I__5422 (
            .O(N__24970),
            .I(N__24967));
    CascadeMux I__5421 (
            .O(N__24967),
            .I(N__24964));
    CascadeBuf I__5420 (
            .O(N__24964),
            .I(N__24961));
    CascadeMux I__5419 (
            .O(N__24961),
            .I(N__24958));
    CascadeBuf I__5418 (
            .O(N__24958),
            .I(N__24955));
    CascadeMux I__5417 (
            .O(N__24955),
            .I(N__24952));
    CascadeBuf I__5416 (
            .O(N__24952),
            .I(N__24949));
    CascadeMux I__5415 (
            .O(N__24949),
            .I(N__24946));
    CascadeBuf I__5414 (
            .O(N__24946),
            .I(N__24943));
    CascadeMux I__5413 (
            .O(N__24943),
            .I(N__24940));
    CascadeBuf I__5412 (
            .O(N__24940),
            .I(N__24937));
    CascadeMux I__5411 (
            .O(N__24937),
            .I(N__24934));
    CascadeBuf I__5410 (
            .O(N__24934),
            .I(N__24931));
    CascadeMux I__5409 (
            .O(N__24931),
            .I(N__24928));
    CascadeBuf I__5408 (
            .O(N__24928),
            .I(N__24925));
    CascadeMux I__5407 (
            .O(N__24925),
            .I(N__24922));
    CascadeBuf I__5406 (
            .O(N__24922),
            .I(N__24919));
    CascadeMux I__5405 (
            .O(N__24919),
            .I(N__24916));
    CascadeBuf I__5404 (
            .O(N__24916),
            .I(N__24913));
    CascadeMux I__5403 (
            .O(N__24913),
            .I(N__24910));
    CascadeBuf I__5402 (
            .O(N__24910),
            .I(N__24907));
    CascadeMux I__5401 (
            .O(N__24907),
            .I(N__24904));
    CascadeBuf I__5400 (
            .O(N__24904),
            .I(N__24901));
    CascadeMux I__5399 (
            .O(N__24901),
            .I(N__24898));
    CascadeBuf I__5398 (
            .O(N__24898),
            .I(N__24895));
    CascadeMux I__5397 (
            .O(N__24895),
            .I(N__24892));
    CascadeBuf I__5396 (
            .O(N__24892),
            .I(N__24889));
    CascadeMux I__5395 (
            .O(N__24889),
            .I(N__24886));
    CascadeBuf I__5394 (
            .O(N__24886),
            .I(N__24883));
    CascadeMux I__5393 (
            .O(N__24883),
            .I(N__24880));
    InMux I__5392 (
            .O(N__24880),
            .I(N__24877));
    LocalMux I__5391 (
            .O(N__24877),
            .I(N__24874));
    Span4Mux_s1_v I__5390 (
            .O(N__24874),
            .I(N__24870));
    CascadeMux I__5389 (
            .O(N__24873),
            .I(N__24867));
    Sp12to4 I__5388 (
            .O(N__24870),
            .I(N__24863));
    InMux I__5387 (
            .O(N__24867),
            .I(N__24860));
    InMux I__5386 (
            .O(N__24866),
            .I(N__24856));
    Span12Mux_s5_v I__5385 (
            .O(N__24863),
            .I(N__24853));
    LocalMux I__5384 (
            .O(N__24860),
            .I(N__24850));
    InMux I__5383 (
            .O(N__24859),
            .I(N__24847));
    LocalMux I__5382 (
            .O(N__24856),
            .I(N__24842));
    Span12Mux_v I__5381 (
            .O(N__24853),
            .I(N__24842));
    Odrv4 I__5380 (
            .O(N__24850),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__5379 (
            .O(N__24847),
            .I(M_this_sprites_address_qZ0Z_5));
    Odrv12 I__5378 (
            .O(N__24842),
            .I(M_this_sprites_address_qZ0Z_5));
    InMux I__5377 (
            .O(N__24835),
            .I(N__24832));
    LocalMux I__5376 (
            .O(N__24832),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5 ));
    InMux I__5375 (
            .O(N__24829),
            .I(N__24826));
    LocalMux I__5374 (
            .O(N__24826),
            .I(N__24823));
    Odrv4 I__5373 (
            .O(N__24823),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_6 ));
    CascadeMux I__5372 (
            .O(N__24820),
            .I(\this_vga_signals.M_this_map_address_d_5_mZ0Z_6_cascade_ ));
    InMux I__5371 (
            .O(N__24817),
            .I(N__24814));
    LocalMux I__5370 (
            .O(N__24814),
            .I(M_this_map_address_q_RNICF7V6Z0Z_0));
    InMux I__5369 (
            .O(N__24811),
            .I(un1_M_this_map_address_q_cry_0));
    CascadeMux I__5368 (
            .O(N__24808),
            .I(N__24805));
    CascadeBuf I__5367 (
            .O(N__24805),
            .I(N__24802));
    CascadeMux I__5366 (
            .O(N__24802),
            .I(N__24799));
    InMux I__5365 (
            .O(N__24799),
            .I(N__24796));
    LocalMux I__5364 (
            .O(N__24796),
            .I(N__24793));
    Span4Mux_s2_v I__5363 (
            .O(N__24793),
            .I(N__24790));
    Span4Mux_h I__5362 (
            .O(N__24790),
            .I(N__24787));
    Span4Mux_h I__5361 (
            .O(N__24787),
            .I(N__24781));
    InMux I__5360 (
            .O(N__24786),
            .I(N__24776));
    InMux I__5359 (
            .O(N__24785),
            .I(N__24776));
    InMux I__5358 (
            .O(N__24784),
            .I(N__24773));
    Span4Mux_v I__5357 (
            .O(N__24781),
            .I(N__24770));
    LocalMux I__5356 (
            .O(N__24776),
            .I(M_this_map_address_qZ0Z_2));
    LocalMux I__5355 (
            .O(N__24773),
            .I(M_this_map_address_qZ0Z_2));
    Odrv4 I__5354 (
            .O(N__24770),
            .I(M_this_map_address_qZ0Z_2));
    InMux I__5353 (
            .O(N__24763),
            .I(N__24760));
    LocalMux I__5352 (
            .O(N__24760),
            .I(un1_M_this_map_address_q_cry_1_c_RNI8JSRZ0));
    InMux I__5351 (
            .O(N__24757),
            .I(un1_M_this_map_address_q_cry_1));
    InMux I__5350 (
            .O(N__24754),
            .I(un1_M_this_map_address_q_cry_2));
    InMux I__5349 (
            .O(N__24751),
            .I(un1_M_this_map_address_q_cry_3));
    CascadeMux I__5348 (
            .O(N__24748),
            .I(N__24745));
    CascadeBuf I__5347 (
            .O(N__24745),
            .I(N__24742));
    CascadeMux I__5346 (
            .O(N__24742),
            .I(N__24739));
    InMux I__5345 (
            .O(N__24739),
            .I(N__24736));
    LocalMux I__5344 (
            .O(N__24736),
            .I(N__24733));
    Sp12to4 I__5343 (
            .O(N__24733),
            .I(N__24727));
    InMux I__5342 (
            .O(N__24732),
            .I(N__24724));
    InMux I__5341 (
            .O(N__24731),
            .I(N__24721));
    InMux I__5340 (
            .O(N__24730),
            .I(N__24718));
    Span12Mux_s11_v I__5339 (
            .O(N__24727),
            .I(N__24715));
    LocalMux I__5338 (
            .O(N__24724),
            .I(M_this_map_address_qZ0Z_5));
    LocalMux I__5337 (
            .O(N__24721),
            .I(M_this_map_address_qZ0Z_5));
    LocalMux I__5336 (
            .O(N__24718),
            .I(M_this_map_address_qZ0Z_5));
    Odrv12 I__5335 (
            .O(N__24715),
            .I(M_this_map_address_qZ0Z_5));
    InMux I__5334 (
            .O(N__24706),
            .I(N__24703));
    LocalMux I__5333 (
            .O(N__24703),
            .I(un1_M_this_map_address_q_cry_4_c_RNIESVRZ0));
    InMux I__5332 (
            .O(N__24700),
            .I(un1_M_this_map_address_q_cry_4));
    CascadeMux I__5331 (
            .O(N__24697),
            .I(N__24694));
    CascadeBuf I__5330 (
            .O(N__24694),
            .I(N__24691));
    CascadeMux I__5329 (
            .O(N__24691),
            .I(N__24688));
    InMux I__5328 (
            .O(N__24688),
            .I(N__24685));
    LocalMux I__5327 (
            .O(N__24685),
            .I(N__24682));
    Span4Mux_v I__5326 (
            .O(N__24682),
            .I(N__24679));
    Sp12to4 I__5325 (
            .O(N__24679),
            .I(N__24673));
    InMux I__5324 (
            .O(N__24678),
            .I(N__24670));
    InMux I__5323 (
            .O(N__24677),
            .I(N__24667));
    InMux I__5322 (
            .O(N__24676),
            .I(N__24664));
    Span12Mux_h I__5321 (
            .O(N__24673),
            .I(N__24661));
    LocalMux I__5320 (
            .O(N__24670),
            .I(M_this_map_address_qZ0Z_6));
    LocalMux I__5319 (
            .O(N__24667),
            .I(M_this_map_address_qZ0Z_6));
    LocalMux I__5318 (
            .O(N__24664),
            .I(M_this_map_address_qZ0Z_6));
    Odrv12 I__5317 (
            .O(N__24661),
            .I(M_this_map_address_qZ0Z_6));
    InMux I__5316 (
            .O(N__24652),
            .I(N__24649));
    LocalMux I__5315 (
            .O(N__24649),
            .I(un1_M_this_map_address_q_cry_5_c_RNIGV0SZ0));
    InMux I__5314 (
            .O(N__24646),
            .I(un1_M_this_map_address_q_cry_5));
    CascadeMux I__5313 (
            .O(N__24643),
            .I(\this_vga_signals.M_this_state_d_1_sqmuxaZ0_cascade_ ));
    CascadeMux I__5312 (
            .O(N__24640),
            .I(N__24637));
    InMux I__5311 (
            .O(N__24637),
            .I(N__24634));
    LocalMux I__5310 (
            .O(N__24634),
            .I(N__24631));
    Span4Mux_v I__5309 (
            .O(N__24631),
            .I(N__24628));
    Odrv4 I__5308 (
            .O(N__24628),
            .I(\this_vga_signals.N_399_0 ));
    InMux I__5307 (
            .O(N__24625),
            .I(N__24622));
    LocalMux I__5306 (
            .O(N__24622),
            .I(\this_vga_signals.M_this_map_address_d_5_mZ0Z_5 ));
    CascadeMux I__5305 (
            .O(N__24619),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_5_cascade_ ));
    CascadeMux I__5304 (
            .O(N__24616),
            .I(N__24613));
    InMux I__5303 (
            .O(N__24613),
            .I(N__24610));
    LocalMux I__5302 (
            .O(N__24610),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_0 ));
    CascadeMux I__5301 (
            .O(N__24607),
            .I(N__24604));
    InMux I__5300 (
            .O(N__24604),
            .I(N__24601));
    LocalMux I__5299 (
            .O(N__24601),
            .I(N__24598));
    Odrv4 I__5298 (
            .O(N__24598),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_11 ));
    InMux I__5297 (
            .O(N__24595),
            .I(N__24591));
    InMux I__5296 (
            .O(N__24594),
            .I(N__24588));
    LocalMux I__5295 (
            .O(N__24591),
            .I(N__24585));
    LocalMux I__5294 (
            .O(N__24588),
            .I(N__24582));
    Odrv12 I__5293 (
            .O(N__24585),
            .I(\this_vga_signals.N_446_1 ));
    Odrv4 I__5292 (
            .O(N__24582),
            .I(\this_vga_signals.N_446_1 ));
    InMux I__5291 (
            .O(N__24577),
            .I(N__24572));
    InMux I__5290 (
            .O(N__24576),
            .I(N__24569));
    CascadeMux I__5289 (
            .O(N__24575),
            .I(N__24563));
    LocalMux I__5288 (
            .O(N__24572),
            .I(N__24556));
    LocalMux I__5287 (
            .O(N__24569),
            .I(N__24556));
    InMux I__5286 (
            .O(N__24568),
            .I(N__24553));
    InMux I__5285 (
            .O(N__24567),
            .I(N__24550));
    InMux I__5284 (
            .O(N__24566),
            .I(N__24543));
    InMux I__5283 (
            .O(N__24563),
            .I(N__24543));
    InMux I__5282 (
            .O(N__24562),
            .I(N__24543));
    InMux I__5281 (
            .O(N__24561),
            .I(N__24540));
    Span4Mux_h I__5280 (
            .O(N__24556),
            .I(N__24537));
    LocalMux I__5279 (
            .O(N__24553),
            .I(N__24532));
    LocalMux I__5278 (
            .O(N__24550),
            .I(N__24532));
    LocalMux I__5277 (
            .O(N__24543),
            .I(N__24529));
    LocalMux I__5276 (
            .O(N__24540),
            .I(N__24526));
    Span4Mux_h I__5275 (
            .O(N__24537),
            .I(N__24520));
    Span12Mux_h I__5274 (
            .O(N__24532),
            .I(N__24517));
    Span4Mux_h I__5273 (
            .O(N__24529),
            .I(N__24514));
    Span4Mux_h I__5272 (
            .O(N__24526),
            .I(N__24511));
    InMux I__5271 (
            .O(N__24525),
            .I(N__24508));
    InMux I__5270 (
            .O(N__24524),
            .I(N__24505));
    InMux I__5269 (
            .O(N__24523),
            .I(N__24502));
    Odrv4 I__5268 (
            .O(N__24520),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv12 I__5267 (
            .O(N__24517),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv4 I__5266 (
            .O(N__24514),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv4 I__5265 (
            .O(N__24511),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__5264 (
            .O(N__24508),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__5263 (
            .O(N__24505),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__5262 (
            .O(N__24502),
            .I(M_this_sprites_address_qZ0Z_11));
    InMux I__5261 (
            .O(N__24487),
            .I(N__24484));
    LocalMux I__5260 (
            .O(N__24484),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11 ));
    CascadeMux I__5259 (
            .O(N__24481),
            .I(N__24477));
    InMux I__5258 (
            .O(N__24480),
            .I(N__24470));
    InMux I__5257 (
            .O(N__24477),
            .I(N__24462));
    InMux I__5256 (
            .O(N__24476),
            .I(N__24459));
    InMux I__5255 (
            .O(N__24475),
            .I(N__24456));
    InMux I__5254 (
            .O(N__24474),
            .I(N__24449));
    InMux I__5253 (
            .O(N__24473),
            .I(N__24449));
    LocalMux I__5252 (
            .O(N__24470),
            .I(N__24446));
    InMux I__5251 (
            .O(N__24469),
            .I(N__24443));
    InMux I__5250 (
            .O(N__24468),
            .I(N__24440));
    CascadeMux I__5249 (
            .O(N__24467),
            .I(N__24437));
    CascadeMux I__5248 (
            .O(N__24466),
            .I(N__24432));
    InMux I__5247 (
            .O(N__24465),
            .I(N__24428));
    LocalMux I__5246 (
            .O(N__24462),
            .I(N__24423));
    LocalMux I__5245 (
            .O(N__24459),
            .I(N__24423));
    LocalMux I__5244 (
            .O(N__24456),
            .I(N__24420));
    InMux I__5243 (
            .O(N__24455),
            .I(N__24414));
    InMux I__5242 (
            .O(N__24454),
            .I(N__24414));
    LocalMux I__5241 (
            .O(N__24449),
            .I(N__24407));
    Span4Mux_h I__5240 (
            .O(N__24446),
            .I(N__24407));
    LocalMux I__5239 (
            .O(N__24443),
            .I(N__24407));
    LocalMux I__5238 (
            .O(N__24440),
            .I(N__24404));
    InMux I__5237 (
            .O(N__24437),
            .I(N__24400));
    InMux I__5236 (
            .O(N__24436),
            .I(N__24397));
    InMux I__5235 (
            .O(N__24435),
            .I(N__24390));
    InMux I__5234 (
            .O(N__24432),
            .I(N__24390));
    InMux I__5233 (
            .O(N__24431),
            .I(N__24390));
    LocalMux I__5232 (
            .O(N__24428),
            .I(N__24387));
    Span4Mux_h I__5231 (
            .O(N__24423),
            .I(N__24382));
    Span4Mux_h I__5230 (
            .O(N__24420),
            .I(N__24382));
    InMux I__5229 (
            .O(N__24419),
            .I(N__24379));
    LocalMux I__5228 (
            .O(N__24414),
            .I(N__24372));
    Span4Mux_v I__5227 (
            .O(N__24407),
            .I(N__24372));
    Span4Mux_h I__5226 (
            .O(N__24404),
            .I(N__24372));
    InMux I__5225 (
            .O(N__24403),
            .I(N__24369));
    LocalMux I__5224 (
            .O(N__24400),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__5223 (
            .O(N__24397),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__5222 (
            .O(N__24390),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__5221 (
            .O(N__24387),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__5220 (
            .O(N__24382),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__5219 (
            .O(N__24379),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__5218 (
            .O(N__24372),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__5217 (
            .O(N__24369),
            .I(M_this_state_qZ0Z_1));
    CascadeMux I__5216 (
            .O(N__24352),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_ ));
    InMux I__5215 (
            .O(N__24349),
            .I(N__24346));
    LocalMux I__5214 (
            .O(N__24346),
            .I(N__24343));
    Odrv4 I__5213 (
            .O(N__24343),
            .I(un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0));
    CascadeMux I__5212 (
            .O(N__24340),
            .I(N__24337));
    CascadeBuf I__5211 (
            .O(N__24337),
            .I(N__24334));
    CascadeMux I__5210 (
            .O(N__24334),
            .I(N__24331));
    CascadeBuf I__5209 (
            .O(N__24331),
            .I(N__24328));
    CascadeMux I__5208 (
            .O(N__24328),
            .I(N__24325));
    CascadeBuf I__5207 (
            .O(N__24325),
            .I(N__24322));
    CascadeMux I__5206 (
            .O(N__24322),
            .I(N__24319));
    CascadeBuf I__5205 (
            .O(N__24319),
            .I(N__24316));
    CascadeMux I__5204 (
            .O(N__24316),
            .I(N__24313));
    CascadeBuf I__5203 (
            .O(N__24313),
            .I(N__24310));
    CascadeMux I__5202 (
            .O(N__24310),
            .I(N__24307));
    CascadeBuf I__5201 (
            .O(N__24307),
            .I(N__24304));
    CascadeMux I__5200 (
            .O(N__24304),
            .I(N__24301));
    CascadeBuf I__5199 (
            .O(N__24301),
            .I(N__24298));
    CascadeMux I__5198 (
            .O(N__24298),
            .I(N__24295));
    CascadeBuf I__5197 (
            .O(N__24295),
            .I(N__24292));
    CascadeMux I__5196 (
            .O(N__24292),
            .I(N__24289));
    CascadeBuf I__5195 (
            .O(N__24289),
            .I(N__24286));
    CascadeMux I__5194 (
            .O(N__24286),
            .I(N__24283));
    CascadeBuf I__5193 (
            .O(N__24283),
            .I(N__24280));
    CascadeMux I__5192 (
            .O(N__24280),
            .I(N__24277));
    CascadeBuf I__5191 (
            .O(N__24277),
            .I(N__24274));
    CascadeMux I__5190 (
            .O(N__24274),
            .I(N__24271));
    CascadeBuf I__5189 (
            .O(N__24271),
            .I(N__24268));
    CascadeMux I__5188 (
            .O(N__24268),
            .I(N__24265));
    CascadeBuf I__5187 (
            .O(N__24265),
            .I(N__24262));
    CascadeMux I__5186 (
            .O(N__24262),
            .I(N__24259));
    CascadeBuf I__5185 (
            .O(N__24259),
            .I(N__24256));
    CascadeMux I__5184 (
            .O(N__24256),
            .I(N__24253));
    CascadeBuf I__5183 (
            .O(N__24253),
            .I(N__24250));
    CascadeMux I__5182 (
            .O(N__24250),
            .I(N__24247));
    InMux I__5181 (
            .O(N__24247),
            .I(N__24244));
    LocalMux I__5180 (
            .O(N__24244),
            .I(N__24241));
    Span4Mux_h I__5179 (
            .O(N__24241),
            .I(N__24237));
    InMux I__5178 (
            .O(N__24240),
            .I(N__24234));
    Sp12to4 I__5177 (
            .O(N__24237),
            .I(N__24229));
    LocalMux I__5176 (
            .O(N__24234),
            .I(N__24226));
    InMux I__5175 (
            .O(N__24233),
            .I(N__24221));
    InMux I__5174 (
            .O(N__24232),
            .I(N__24221));
    Span12Mux_v I__5173 (
            .O(N__24229),
            .I(N__24218));
    Odrv4 I__5172 (
            .O(N__24226),
            .I(M_this_sprites_address_qZ0Z_7));
    LocalMux I__5171 (
            .O(N__24221),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv12 I__5170 (
            .O(N__24218),
            .I(M_this_sprites_address_qZ0Z_7));
    InMux I__5169 (
            .O(N__24211),
            .I(N__24208));
    LocalMux I__5168 (
            .O(N__24208),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_7 ));
    InMux I__5167 (
            .O(N__24205),
            .I(N__24202));
    LocalMux I__5166 (
            .O(N__24202),
            .I(N__24199));
    Odrv4 I__5165 (
            .O(N__24199),
            .I(un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0));
    CascadeMux I__5164 (
            .O(N__24196),
            .I(N__24193));
    InMux I__5163 (
            .O(N__24193),
            .I(N__24190));
    LocalMux I__5162 (
            .O(N__24190),
            .I(N__24187));
    Span4Mux_h I__5161 (
            .O(N__24187),
            .I(N__24184));
    Odrv4 I__5160 (
            .O(N__24184),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_4 ));
    InMux I__5159 (
            .O(N__24181),
            .I(N__24176));
    InMux I__5158 (
            .O(N__24180),
            .I(N__24165));
    InMux I__5157 (
            .O(N__24179),
            .I(N__24165));
    LocalMux I__5156 (
            .O(N__24176),
            .I(N__24162));
    InMux I__5155 (
            .O(N__24175),
            .I(N__24159));
    InMux I__5154 (
            .O(N__24174),
            .I(N__24152));
    InMux I__5153 (
            .O(N__24173),
            .I(N__24152));
    InMux I__5152 (
            .O(N__24172),
            .I(N__24152));
    InMux I__5151 (
            .O(N__24171),
            .I(N__24144));
    InMux I__5150 (
            .O(N__24170),
            .I(N__24144));
    LocalMux I__5149 (
            .O(N__24165),
            .I(N__24139));
    Span4Mux_v I__5148 (
            .O(N__24162),
            .I(N__24132));
    LocalMux I__5147 (
            .O(N__24159),
            .I(N__24132));
    LocalMux I__5146 (
            .O(N__24152),
            .I(N__24132));
    InMux I__5145 (
            .O(N__24151),
            .I(N__24129));
    InMux I__5144 (
            .O(N__24150),
            .I(N__24124));
    InMux I__5143 (
            .O(N__24149),
            .I(N__24124));
    LocalMux I__5142 (
            .O(N__24144),
            .I(N__24121));
    InMux I__5141 (
            .O(N__24143),
            .I(N__24116));
    InMux I__5140 (
            .O(N__24142),
            .I(N__24116));
    Odrv4 I__5139 (
            .O(N__24139),
            .I(\this_vga_signals.un1_M_this_state_q_19_0 ));
    Odrv4 I__5138 (
            .O(N__24132),
            .I(\this_vga_signals.un1_M_this_state_q_19_0 ));
    LocalMux I__5137 (
            .O(N__24129),
            .I(\this_vga_signals.un1_M_this_state_q_19_0 ));
    LocalMux I__5136 (
            .O(N__24124),
            .I(\this_vga_signals.un1_M_this_state_q_19_0 ));
    Odrv4 I__5135 (
            .O(N__24121),
            .I(\this_vga_signals.un1_M_this_state_q_19_0 ));
    LocalMux I__5134 (
            .O(N__24116),
            .I(\this_vga_signals.un1_M_this_state_q_19_0 ));
    CascadeMux I__5133 (
            .O(N__24103),
            .I(\this_vga_signals.N_294_cascade_ ));
    CascadeMux I__5132 (
            .O(N__24100),
            .I(\this_vga_signals.un1_M_this_state_q_14Z0Z_1_cascade_ ));
    CascadeMux I__5131 (
            .O(N__24097),
            .I(N__24092));
    InMux I__5130 (
            .O(N__24096),
            .I(N__24089));
    InMux I__5129 (
            .O(N__24095),
            .I(N__24086));
    InMux I__5128 (
            .O(N__24092),
            .I(N__24083));
    LocalMux I__5127 (
            .O(N__24089),
            .I(un1_M_this_state_q_14_0));
    LocalMux I__5126 (
            .O(N__24086),
            .I(un1_M_this_state_q_14_0));
    LocalMux I__5125 (
            .O(N__24083),
            .I(un1_M_this_state_q_14_0));
    CascadeMux I__5124 (
            .O(N__24076),
            .I(N__24073));
    InMux I__5123 (
            .O(N__24073),
            .I(N__24069));
    InMux I__5122 (
            .O(N__24072),
            .I(N__24066));
    LocalMux I__5121 (
            .O(N__24069),
            .I(this_vga_signals_un23_i_a2_1_1));
    LocalMux I__5120 (
            .O(N__24066),
            .I(this_vga_signals_un23_i_a2_1_1));
    InMux I__5119 (
            .O(N__24061),
            .I(N__24058));
    LocalMux I__5118 (
            .O(N__24058),
            .I(N__24055));
    Odrv4 I__5117 (
            .O(N__24055),
            .I(un23_i_a2_1));
    InMux I__5116 (
            .O(N__24052),
            .I(N__24049));
    LocalMux I__5115 (
            .O(N__24049),
            .I(N__24046));
    Odrv4 I__5114 (
            .O(N__24046),
            .I(\this_vga_signals.N_486 ));
    InMux I__5113 (
            .O(N__24043),
            .I(N__24039));
    CascadeMux I__5112 (
            .O(N__24042),
            .I(N__24036));
    LocalMux I__5111 (
            .O(N__24039),
            .I(N__24033));
    InMux I__5110 (
            .O(N__24036),
            .I(N__24030));
    Span4Mux_v I__5109 (
            .O(N__24033),
            .I(N__24027));
    LocalMux I__5108 (
            .O(N__24030),
            .I(N__24024));
    Odrv4 I__5107 (
            .O(N__24027),
            .I(\this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_5 ));
    Odrv4 I__5106 (
            .O(N__24024),
            .I(\this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_5 ));
    CascadeMux I__5105 (
            .O(N__24019),
            .I(\this_vga_signals.N_486_cascade_ ));
    InMux I__5104 (
            .O(N__24016),
            .I(N__24013));
    LocalMux I__5103 (
            .O(N__24013),
            .I(N__24009));
    InMux I__5102 (
            .O(N__24012),
            .I(N__24006));
    Span4Mux_v I__5101 (
            .O(N__24009),
            .I(N__24001));
    LocalMux I__5100 (
            .O(N__24006),
            .I(N__24001));
    Span4Mux_v I__5099 (
            .O(N__24001),
            .I(N__23998));
    Odrv4 I__5098 (
            .O(N__23998),
            .I(\this_vga_signals.N_438_1 ));
    CascadeMux I__5097 (
            .O(N__23995),
            .I(N__23992));
    InMux I__5096 (
            .O(N__23992),
            .I(N__23989));
    LocalMux I__5095 (
            .O(N__23989),
            .I(N__23986));
    Odrv12 I__5094 (
            .O(N__23986),
            .I(this_vga_signals_M_this_state_q_ns_i_o2_0_12));
    InMux I__5093 (
            .O(N__23983),
            .I(N__23977));
    InMux I__5092 (
            .O(N__23982),
            .I(N__23977));
    LocalMux I__5091 (
            .O(N__23977),
            .I(N__23972));
    InMux I__5090 (
            .O(N__23976),
            .I(N__23969));
    InMux I__5089 (
            .O(N__23975),
            .I(N__23966));
    Odrv4 I__5088 (
            .O(N__23972),
            .I(\this_ppu.un1_M_haddress_q_c2 ));
    LocalMux I__5087 (
            .O(N__23969),
            .I(\this_ppu.un1_M_haddress_q_c2 ));
    LocalMux I__5086 (
            .O(N__23966),
            .I(\this_ppu.un1_M_haddress_q_c2 ));
    CascadeMux I__5085 (
            .O(N__23959),
            .I(N__23955));
    CascadeMux I__5084 (
            .O(N__23958),
            .I(N__23952));
    CascadeBuf I__5083 (
            .O(N__23955),
            .I(N__23949));
    InMux I__5082 (
            .O(N__23952),
            .I(N__23946));
    CascadeMux I__5081 (
            .O(N__23949),
            .I(N__23943));
    LocalMux I__5080 (
            .O(N__23946),
            .I(N__23940));
    InMux I__5079 (
            .O(N__23943),
            .I(N__23937));
    Span4Mux_h I__5078 (
            .O(N__23940),
            .I(N__23934));
    LocalMux I__5077 (
            .O(N__23937),
            .I(N__23931));
    Span4Mux_v I__5076 (
            .O(N__23934),
            .I(N__23927));
    Span4Mux_s2_v I__5075 (
            .O(N__23931),
            .I(N__23924));
    CascadeMux I__5074 (
            .O(N__23930),
            .I(N__23921));
    Span4Mux_v I__5073 (
            .O(N__23927),
            .I(N__23916));
    Span4Mux_h I__5072 (
            .O(N__23924),
            .I(N__23913));
    InMux I__5071 (
            .O(N__23921),
            .I(N__23908));
    InMux I__5070 (
            .O(N__23920),
            .I(N__23908));
    InMux I__5069 (
            .O(N__23919),
            .I(N__23905));
    Span4Mux_h I__5068 (
            .O(N__23916),
            .I(N__23900));
    Span4Mux_v I__5067 (
            .O(N__23913),
            .I(N__23900));
    LocalMux I__5066 (
            .O(N__23908),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__5065 (
            .O(N__23905),
            .I(M_this_ppu_map_addr_0));
    Odrv4 I__5064 (
            .O(N__23900),
            .I(M_this_ppu_map_addr_0));
    InMux I__5063 (
            .O(N__23893),
            .I(N__23890));
    LocalMux I__5062 (
            .O(N__23890),
            .I(N__23887));
    Span4Mux_v I__5061 (
            .O(N__23887),
            .I(N__23882));
    InMux I__5060 (
            .O(N__23886),
            .I(N__23878));
    InMux I__5059 (
            .O(N__23885),
            .I(N__23875));
    Span4Mux_h I__5058 (
            .O(N__23882),
            .I(N__23872));
    InMux I__5057 (
            .O(N__23881),
            .I(N__23869));
    LocalMux I__5056 (
            .O(N__23878),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    LocalMux I__5055 (
            .O(N__23875),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    Odrv4 I__5054 (
            .O(N__23872),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    LocalMux I__5053 (
            .O(N__23869),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    CascadeMux I__5052 (
            .O(N__23860),
            .I(N__23857));
    CascadeBuf I__5051 (
            .O(N__23857),
            .I(N__23854));
    CascadeMux I__5050 (
            .O(N__23854),
            .I(N__23851));
    InMux I__5049 (
            .O(N__23851),
            .I(N__23848));
    LocalMux I__5048 (
            .O(N__23848),
            .I(N__23845));
    Span4Mux_h I__5047 (
            .O(N__23845),
            .I(N__23842));
    Span4Mux_h I__5046 (
            .O(N__23842),
            .I(N__23839));
    Odrv4 I__5045 (
            .O(N__23839),
            .I(this_ppu_M_vaddress_q_i_6));
    InMux I__5044 (
            .O(N__23836),
            .I(N__23833));
    LocalMux I__5043 (
            .O(N__23833),
            .I(N__23830));
    Span4Mux_h I__5042 (
            .O(N__23830),
            .I(N__23827));
    Odrv4 I__5041 (
            .O(N__23827),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_6 ));
    CascadeMux I__5040 (
            .O(N__23824),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6_cascade_ ));
    InMux I__5039 (
            .O(N__23821),
            .I(N__23818));
    LocalMux I__5038 (
            .O(N__23818),
            .I(N__23815));
    Odrv4 I__5037 (
            .O(N__23815),
            .I(un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0));
    CascadeMux I__5036 (
            .O(N__23812),
            .I(N__23809));
    CascadeBuf I__5035 (
            .O(N__23809),
            .I(N__23806));
    CascadeMux I__5034 (
            .O(N__23806),
            .I(N__23803));
    CascadeBuf I__5033 (
            .O(N__23803),
            .I(N__23800));
    CascadeMux I__5032 (
            .O(N__23800),
            .I(N__23797));
    CascadeBuf I__5031 (
            .O(N__23797),
            .I(N__23794));
    CascadeMux I__5030 (
            .O(N__23794),
            .I(N__23791));
    CascadeBuf I__5029 (
            .O(N__23791),
            .I(N__23788));
    CascadeMux I__5028 (
            .O(N__23788),
            .I(N__23785));
    CascadeBuf I__5027 (
            .O(N__23785),
            .I(N__23782));
    CascadeMux I__5026 (
            .O(N__23782),
            .I(N__23779));
    CascadeBuf I__5025 (
            .O(N__23779),
            .I(N__23776));
    CascadeMux I__5024 (
            .O(N__23776),
            .I(N__23773));
    CascadeBuf I__5023 (
            .O(N__23773),
            .I(N__23770));
    CascadeMux I__5022 (
            .O(N__23770),
            .I(N__23767));
    CascadeBuf I__5021 (
            .O(N__23767),
            .I(N__23764));
    CascadeMux I__5020 (
            .O(N__23764),
            .I(N__23761));
    CascadeBuf I__5019 (
            .O(N__23761),
            .I(N__23758));
    CascadeMux I__5018 (
            .O(N__23758),
            .I(N__23755));
    CascadeBuf I__5017 (
            .O(N__23755),
            .I(N__23752));
    CascadeMux I__5016 (
            .O(N__23752),
            .I(N__23749));
    CascadeBuf I__5015 (
            .O(N__23749),
            .I(N__23746));
    CascadeMux I__5014 (
            .O(N__23746),
            .I(N__23743));
    CascadeBuf I__5013 (
            .O(N__23743),
            .I(N__23740));
    CascadeMux I__5012 (
            .O(N__23740),
            .I(N__23737));
    CascadeBuf I__5011 (
            .O(N__23737),
            .I(N__23734));
    CascadeMux I__5010 (
            .O(N__23734),
            .I(N__23731));
    CascadeBuf I__5009 (
            .O(N__23731),
            .I(N__23728));
    CascadeMux I__5008 (
            .O(N__23728),
            .I(N__23725));
    CascadeBuf I__5007 (
            .O(N__23725),
            .I(N__23722));
    CascadeMux I__5006 (
            .O(N__23722),
            .I(N__23719));
    InMux I__5005 (
            .O(N__23719),
            .I(N__23716));
    LocalMux I__5004 (
            .O(N__23716),
            .I(N__23713));
    Span4Mux_v I__5003 (
            .O(N__23713),
            .I(N__23708));
    InMux I__5002 (
            .O(N__23712),
            .I(N__23705));
    InMux I__5001 (
            .O(N__23711),
            .I(N__23702));
    Span4Mux_v I__5000 (
            .O(N__23708),
            .I(N__23699));
    LocalMux I__4999 (
            .O(N__23705),
            .I(N__23696));
    LocalMux I__4998 (
            .O(N__23702),
            .I(N__23692));
    Sp12to4 I__4997 (
            .O(N__23699),
            .I(N__23689));
    Span4Mux_v I__4996 (
            .O(N__23696),
            .I(N__23686));
    InMux I__4995 (
            .O(N__23695),
            .I(N__23683));
    Sp12to4 I__4994 (
            .O(N__23692),
            .I(N__23678));
    Span12Mux_h I__4993 (
            .O(N__23689),
            .I(N__23678));
    Odrv4 I__4992 (
            .O(N__23686),
            .I(M_this_sprites_address_qZ0Z_6));
    LocalMux I__4991 (
            .O(N__23683),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv12 I__4990 (
            .O(N__23678),
            .I(M_this_sprites_address_qZ0Z_6));
    CascadeMux I__4989 (
            .O(N__23671),
            .I(N__23668));
    InMux I__4988 (
            .O(N__23668),
            .I(N__23665));
    LocalMux I__4987 (
            .O(N__23665),
            .I(N__23662));
    Span4Mux_v I__4986 (
            .O(N__23662),
            .I(N__23659));
    Odrv4 I__4985 (
            .O(N__23659),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_0 ));
    CascadeMux I__4984 (
            .O(N__23656),
            .I(N__23653));
    InMux I__4983 (
            .O(N__23653),
            .I(N__23650));
    LocalMux I__4982 (
            .O(N__23650),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_5 ));
    InMux I__4981 (
            .O(N__23647),
            .I(N__23644));
    LocalMux I__4980 (
            .O(N__23644),
            .I(N__23641));
    Odrv4 I__4979 (
            .O(N__23641),
            .I(un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0));
    CascadeMux I__4978 (
            .O(N__23638),
            .I(N__23635));
    InMux I__4977 (
            .O(N__23635),
            .I(N__23632));
    LocalMux I__4976 (
            .O(N__23632),
            .I(N__23629));
    Odrv4 I__4975 (
            .O(N__23629),
            .I(\this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_6 ));
    CascadeMux I__4974 (
            .O(N__23626),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_2_cascade_ ));
    InMux I__4973 (
            .O(N__23623),
            .I(N__23620));
    LocalMux I__4972 (
            .O(N__23620),
            .I(\this_vga_signals.M_this_map_address_d_8_mZ0Z_2 ));
    InMux I__4971 (
            .O(N__23617),
            .I(N__23614));
    LocalMux I__4970 (
            .O(N__23614),
            .I(N__23611));
    Span4Mux_h I__4969 (
            .O(N__23611),
            .I(N__23608));
    Odrv4 I__4968 (
            .O(N__23608),
            .I(\this_vga_signals.M_this_map_address_q_mZ0Z_9 ));
    CascadeMux I__4967 (
            .O(N__23605),
            .I(N__23602));
    InMux I__4966 (
            .O(N__23602),
            .I(N__23599));
    LocalMux I__4965 (
            .O(N__23599),
            .I(\this_vga_signals.M_this_map_address_d_5_mZ0Z_9 ));
    CascadeMux I__4964 (
            .O(N__23596),
            .I(N__23592));
    CascadeMux I__4963 (
            .O(N__23595),
            .I(N__23589));
    InMux I__4962 (
            .O(N__23592),
            .I(N__23586));
    CascadeBuf I__4961 (
            .O(N__23589),
            .I(N__23583));
    LocalMux I__4960 (
            .O(N__23586),
            .I(N__23580));
    CascadeMux I__4959 (
            .O(N__23583),
            .I(N__23577));
    Span4Mux_h I__4958 (
            .O(N__23580),
            .I(N__23574));
    InMux I__4957 (
            .O(N__23577),
            .I(N__23571));
    Span4Mux_h I__4956 (
            .O(N__23574),
            .I(N__23566));
    LocalMux I__4955 (
            .O(N__23571),
            .I(N__23563));
    InMux I__4954 (
            .O(N__23570),
            .I(N__23560));
    InMux I__4953 (
            .O(N__23569),
            .I(N__23557));
    Sp12to4 I__4952 (
            .O(N__23566),
            .I(N__23552));
    Span12Mux_h I__4951 (
            .O(N__23563),
            .I(N__23552));
    LocalMux I__4950 (
            .O(N__23560),
            .I(M_this_ppu_map_addr_1));
    LocalMux I__4949 (
            .O(N__23557),
            .I(M_this_ppu_map_addr_1));
    Odrv12 I__4948 (
            .O(N__23552),
            .I(M_this_ppu_map_addr_1));
    CascadeMux I__4947 (
            .O(N__23545),
            .I(N__23542));
    CascadeBuf I__4946 (
            .O(N__23542),
            .I(N__23539));
    CascadeMux I__4945 (
            .O(N__23539),
            .I(N__23536));
    CascadeBuf I__4944 (
            .O(N__23536),
            .I(N__23533));
    CascadeMux I__4943 (
            .O(N__23533),
            .I(N__23530));
    CascadeBuf I__4942 (
            .O(N__23530),
            .I(N__23527));
    CascadeMux I__4941 (
            .O(N__23527),
            .I(N__23524));
    CascadeBuf I__4940 (
            .O(N__23524),
            .I(N__23521));
    CascadeMux I__4939 (
            .O(N__23521),
            .I(N__23518));
    CascadeBuf I__4938 (
            .O(N__23518),
            .I(N__23515));
    CascadeMux I__4937 (
            .O(N__23515),
            .I(N__23512));
    CascadeBuf I__4936 (
            .O(N__23512),
            .I(N__23509));
    CascadeMux I__4935 (
            .O(N__23509),
            .I(N__23506));
    CascadeBuf I__4934 (
            .O(N__23506),
            .I(N__23503));
    CascadeMux I__4933 (
            .O(N__23503),
            .I(N__23500));
    CascadeBuf I__4932 (
            .O(N__23500),
            .I(N__23497));
    CascadeMux I__4931 (
            .O(N__23497),
            .I(N__23494));
    CascadeBuf I__4930 (
            .O(N__23494),
            .I(N__23491));
    CascadeMux I__4929 (
            .O(N__23491),
            .I(N__23488));
    CascadeBuf I__4928 (
            .O(N__23488),
            .I(N__23485));
    CascadeMux I__4927 (
            .O(N__23485),
            .I(N__23482));
    CascadeBuf I__4926 (
            .O(N__23482),
            .I(N__23479));
    CascadeMux I__4925 (
            .O(N__23479),
            .I(N__23476));
    CascadeBuf I__4924 (
            .O(N__23476),
            .I(N__23473));
    CascadeMux I__4923 (
            .O(N__23473),
            .I(N__23470));
    CascadeBuf I__4922 (
            .O(N__23470),
            .I(N__23467));
    CascadeMux I__4921 (
            .O(N__23467),
            .I(N__23464));
    CascadeBuf I__4920 (
            .O(N__23464),
            .I(N__23461));
    CascadeMux I__4919 (
            .O(N__23461),
            .I(N__23458));
    CascadeBuf I__4918 (
            .O(N__23458),
            .I(N__23455));
    CascadeMux I__4917 (
            .O(N__23455),
            .I(N__23451));
    CascadeMux I__4916 (
            .O(N__23454),
            .I(N__23448));
    InMux I__4915 (
            .O(N__23451),
            .I(N__23445));
    InMux I__4914 (
            .O(N__23448),
            .I(N__23442));
    LocalMux I__4913 (
            .O(N__23445),
            .I(N__23439));
    LocalMux I__4912 (
            .O(N__23442),
            .I(N__23435));
    Span4Mux_v I__4911 (
            .O(N__23439),
            .I(N__23432));
    CascadeMux I__4910 (
            .O(N__23438),
            .I(N__23429));
    Sp12to4 I__4909 (
            .O(N__23435),
            .I(N__23423));
    Span4Mux_h I__4908 (
            .O(N__23432),
            .I(N__23420));
    InMux I__4907 (
            .O(N__23429),
            .I(N__23417));
    InMux I__4906 (
            .O(N__23428),
            .I(N__23414));
    InMux I__4905 (
            .O(N__23427),
            .I(N__23409));
    InMux I__4904 (
            .O(N__23426),
            .I(N__23409));
    Span12Mux_v I__4903 (
            .O(N__23423),
            .I(N__23406));
    Span4Mux_h I__4902 (
            .O(N__23420),
            .I(N__23403));
    LocalMux I__4901 (
            .O(N__23417),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__4900 (
            .O(N__23414),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__4899 (
            .O(N__23409),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__4898 (
            .O(N__23406),
            .I(M_this_ppu_vram_addr_2));
    Odrv4 I__4897 (
            .O(N__23403),
            .I(M_this_ppu_vram_addr_2));
    InMux I__4896 (
            .O(N__23392),
            .I(N__23389));
    LocalMux I__4895 (
            .O(N__23389),
            .I(un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0));
    InMux I__4894 (
            .O(N__23386),
            .I(N__23383));
    LocalMux I__4893 (
            .O(N__23383),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12 ));
    InMux I__4892 (
            .O(N__23380),
            .I(N__23377));
    LocalMux I__4891 (
            .O(N__23377),
            .I(un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0));
    InMux I__4890 (
            .O(N__23374),
            .I(N__23371));
    LocalMux I__4889 (
            .O(N__23371),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13 ));
    CascadeMux I__4888 (
            .O(N__23368),
            .I(N__23365));
    InMux I__4887 (
            .O(N__23365),
            .I(N__23362));
    LocalMux I__4886 (
            .O(N__23362),
            .I(N__23359));
    Odrv4 I__4885 (
            .O(N__23359),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_13 ));
    InMux I__4884 (
            .O(N__23356),
            .I(N__23353));
    LocalMux I__4883 (
            .O(N__23353),
            .I(un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0));
    CascadeMux I__4882 (
            .O(N__23350),
            .I(N__23344));
    CascadeMux I__4881 (
            .O(N__23349),
            .I(N__23341));
    CascadeMux I__4880 (
            .O(N__23348),
            .I(N__23336));
    CascadeMux I__4879 (
            .O(N__23347),
            .I(N__23333));
    InMux I__4878 (
            .O(N__23344),
            .I(N__23330));
    InMux I__4877 (
            .O(N__23341),
            .I(N__23327));
    CascadeMux I__4876 (
            .O(N__23340),
            .I(N__23324));
    CascadeMux I__4875 (
            .O(N__23339),
            .I(N__23320));
    InMux I__4874 (
            .O(N__23336),
            .I(N__23316));
    InMux I__4873 (
            .O(N__23333),
            .I(N__23313));
    LocalMux I__4872 (
            .O(N__23330),
            .I(N__23310));
    LocalMux I__4871 (
            .O(N__23327),
            .I(N__23307));
    InMux I__4870 (
            .O(N__23324),
            .I(N__23300));
    InMux I__4869 (
            .O(N__23323),
            .I(N__23300));
    InMux I__4868 (
            .O(N__23320),
            .I(N__23300));
    CascadeMux I__4867 (
            .O(N__23319),
            .I(N__23297));
    LocalMux I__4866 (
            .O(N__23316),
            .I(N__23294));
    LocalMux I__4865 (
            .O(N__23313),
            .I(N__23290));
    Span4Mux_v I__4864 (
            .O(N__23310),
            .I(N__23285));
    Span4Mux_v I__4863 (
            .O(N__23307),
            .I(N__23285));
    LocalMux I__4862 (
            .O(N__23300),
            .I(N__23282));
    InMux I__4861 (
            .O(N__23297),
            .I(N__23279));
    Span4Mux_h I__4860 (
            .O(N__23294),
            .I(N__23276));
    InMux I__4859 (
            .O(N__23293),
            .I(N__23273));
    Span12Mux_v I__4858 (
            .O(N__23290),
            .I(N__23268));
    Span4Mux_h I__4857 (
            .O(N__23285),
            .I(N__23263));
    Span4Mux_v I__4856 (
            .O(N__23282),
            .I(N__23263));
    LocalMux I__4855 (
            .O(N__23279),
            .I(N__23260));
    Span4Mux_h I__4854 (
            .O(N__23276),
            .I(N__23255));
    LocalMux I__4853 (
            .O(N__23273),
            .I(N__23255));
    InMux I__4852 (
            .O(N__23272),
            .I(N__23252));
    InMux I__4851 (
            .O(N__23271),
            .I(N__23249));
    Odrv12 I__4850 (
            .O(N__23268),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__4849 (
            .O(N__23263),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__4848 (
            .O(N__23260),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__4847 (
            .O(N__23255),
            .I(M_this_sprites_address_qZ0Z_13));
    LocalMux I__4846 (
            .O(N__23252),
            .I(M_this_sprites_address_qZ0Z_13));
    LocalMux I__4845 (
            .O(N__23249),
            .I(M_this_sprites_address_qZ0Z_13));
    InMux I__4844 (
            .O(N__23236),
            .I(N__23233));
    LocalMux I__4843 (
            .O(N__23233),
            .I(N__23230));
    Odrv12 I__4842 (
            .O(N__23230),
            .I(\this_vga_signals.M_this_state_q_ns_0_o2_0_0_0 ));
    CascadeMux I__4841 (
            .O(N__23227),
            .I(\this_vga_signals.M_this_state_q_ns_0_o2_0_1Z0Z_0_cascade_ ));
    InMux I__4840 (
            .O(N__23224),
            .I(N__23221));
    LocalMux I__4839 (
            .O(N__23221),
            .I(N__23218));
    Odrv12 I__4838 (
            .O(N__23218),
            .I(M_this_sprites_address_q_RNI1DGI7Z0Z_0));
    InMux I__4837 (
            .O(N__23215),
            .I(N__23212));
    LocalMux I__4836 (
            .O(N__23212),
            .I(N__23209));
    Span12Mux_h I__4835 (
            .O(N__23209),
            .I(N__23206));
    Odrv12 I__4834 (
            .O(N__23206),
            .I(M_this_map_ram_read_data_5));
    CascadeMux I__4833 (
            .O(N__23203),
            .I(N__23200));
    InMux I__4832 (
            .O(N__23200),
            .I(N__23193));
    CascadeMux I__4831 (
            .O(N__23199),
            .I(N__23189));
    InMux I__4830 (
            .O(N__23198),
            .I(N__23186));
    InMux I__4829 (
            .O(N__23197),
            .I(N__23180));
    InMux I__4828 (
            .O(N__23196),
            .I(N__23180));
    LocalMux I__4827 (
            .O(N__23193),
            .I(N__23177));
    InMux I__4826 (
            .O(N__23192),
            .I(N__23174));
    InMux I__4825 (
            .O(N__23189),
            .I(N__23171));
    LocalMux I__4824 (
            .O(N__23186),
            .I(N__23168));
    InMux I__4823 (
            .O(N__23185),
            .I(N__23165));
    LocalMux I__4822 (
            .O(N__23180),
            .I(N__23162));
    Span4Mux_h I__4821 (
            .O(N__23177),
            .I(N__23154));
    LocalMux I__4820 (
            .O(N__23174),
            .I(N__23154));
    LocalMux I__4819 (
            .O(N__23171),
            .I(N__23154));
    Span4Mux_v I__4818 (
            .O(N__23168),
            .I(N__23149));
    LocalMux I__4817 (
            .O(N__23165),
            .I(N__23149));
    Span4Mux_v I__4816 (
            .O(N__23162),
            .I(N__23146));
    InMux I__4815 (
            .O(N__23161),
            .I(N__23143));
    Span4Mux_h I__4814 (
            .O(N__23154),
            .I(N__23140));
    Span4Mux_h I__4813 (
            .O(N__23149),
            .I(N__23137));
    Sp12to4 I__4812 (
            .O(N__23146),
            .I(N__23132));
    LocalMux I__4811 (
            .O(N__23143),
            .I(N__23132));
    Span4Mux_v I__4810 (
            .O(N__23140),
            .I(N__23129));
    Sp12to4 I__4809 (
            .O(N__23137),
            .I(N__23124));
    Span12Mux_h I__4808 (
            .O(N__23132),
            .I(N__23124));
    Odrv4 I__4807 (
            .O(N__23129),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    Odrv12 I__4806 (
            .O(N__23124),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    InMux I__4805 (
            .O(N__23119),
            .I(un1_M_this_sprites_address_q_cry_5));
    InMux I__4804 (
            .O(N__23116),
            .I(un1_M_this_sprites_address_q_cry_6));
    CascadeMux I__4803 (
            .O(N__23113),
            .I(N__23110));
    CascadeBuf I__4802 (
            .O(N__23110),
            .I(N__23107));
    CascadeMux I__4801 (
            .O(N__23107),
            .I(N__23104));
    CascadeBuf I__4800 (
            .O(N__23104),
            .I(N__23101));
    CascadeMux I__4799 (
            .O(N__23101),
            .I(N__23098));
    CascadeBuf I__4798 (
            .O(N__23098),
            .I(N__23095));
    CascadeMux I__4797 (
            .O(N__23095),
            .I(N__23092));
    CascadeBuf I__4796 (
            .O(N__23092),
            .I(N__23089));
    CascadeMux I__4795 (
            .O(N__23089),
            .I(N__23086));
    CascadeBuf I__4794 (
            .O(N__23086),
            .I(N__23083));
    CascadeMux I__4793 (
            .O(N__23083),
            .I(N__23080));
    CascadeBuf I__4792 (
            .O(N__23080),
            .I(N__23077));
    CascadeMux I__4791 (
            .O(N__23077),
            .I(N__23074));
    CascadeBuf I__4790 (
            .O(N__23074),
            .I(N__23071));
    CascadeMux I__4789 (
            .O(N__23071),
            .I(N__23068));
    CascadeBuf I__4788 (
            .O(N__23068),
            .I(N__23065));
    CascadeMux I__4787 (
            .O(N__23065),
            .I(N__23062));
    CascadeBuf I__4786 (
            .O(N__23062),
            .I(N__23059));
    CascadeMux I__4785 (
            .O(N__23059),
            .I(N__23056));
    CascadeBuf I__4784 (
            .O(N__23056),
            .I(N__23053));
    CascadeMux I__4783 (
            .O(N__23053),
            .I(N__23050));
    CascadeBuf I__4782 (
            .O(N__23050),
            .I(N__23047));
    CascadeMux I__4781 (
            .O(N__23047),
            .I(N__23044));
    CascadeBuf I__4780 (
            .O(N__23044),
            .I(N__23041));
    CascadeMux I__4779 (
            .O(N__23041),
            .I(N__23038));
    CascadeBuf I__4778 (
            .O(N__23038),
            .I(N__23035));
    CascadeMux I__4777 (
            .O(N__23035),
            .I(N__23032));
    CascadeBuf I__4776 (
            .O(N__23032),
            .I(N__23029));
    CascadeMux I__4775 (
            .O(N__23029),
            .I(N__23026));
    CascadeBuf I__4774 (
            .O(N__23026),
            .I(N__23023));
    CascadeMux I__4773 (
            .O(N__23023),
            .I(N__23020));
    InMux I__4772 (
            .O(N__23020),
            .I(N__23017));
    LocalMux I__4771 (
            .O(N__23017),
            .I(N__23014));
    Span4Mux_s1_v I__4770 (
            .O(N__23014),
            .I(N__23011));
    Sp12to4 I__4769 (
            .O(N__23011),
            .I(N__23006));
    InMux I__4768 (
            .O(N__23010),
            .I(N__23003));
    InMux I__4767 (
            .O(N__23009),
            .I(N__22999));
    Span12Mux_h I__4766 (
            .O(N__23006),
            .I(N__22996));
    LocalMux I__4765 (
            .O(N__23003),
            .I(N__22993));
    InMux I__4764 (
            .O(N__23002),
            .I(N__22990));
    LocalMux I__4763 (
            .O(N__22999),
            .I(N__22985));
    Span12Mux_v I__4762 (
            .O(N__22996),
            .I(N__22985));
    Odrv4 I__4761 (
            .O(N__22993),
            .I(M_this_sprites_address_qZ0Z_8));
    LocalMux I__4760 (
            .O(N__22990),
            .I(M_this_sprites_address_qZ0Z_8));
    Odrv12 I__4759 (
            .O(N__22985),
            .I(M_this_sprites_address_qZ0Z_8));
    InMux I__4758 (
            .O(N__22978),
            .I(N__22975));
    LocalMux I__4757 (
            .O(N__22975),
            .I(N__22972));
    Odrv4 I__4756 (
            .O(N__22972),
            .I(un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0));
    InMux I__4755 (
            .O(N__22969),
            .I(bfn_18_18_0_));
    CascadeMux I__4754 (
            .O(N__22966),
            .I(N__22963));
    CascadeBuf I__4753 (
            .O(N__22963),
            .I(N__22960));
    CascadeMux I__4752 (
            .O(N__22960),
            .I(N__22957));
    CascadeBuf I__4751 (
            .O(N__22957),
            .I(N__22954));
    CascadeMux I__4750 (
            .O(N__22954),
            .I(N__22951));
    CascadeBuf I__4749 (
            .O(N__22951),
            .I(N__22948));
    CascadeMux I__4748 (
            .O(N__22948),
            .I(N__22945));
    CascadeBuf I__4747 (
            .O(N__22945),
            .I(N__22942));
    CascadeMux I__4746 (
            .O(N__22942),
            .I(N__22939));
    CascadeBuf I__4745 (
            .O(N__22939),
            .I(N__22936));
    CascadeMux I__4744 (
            .O(N__22936),
            .I(N__22933));
    CascadeBuf I__4743 (
            .O(N__22933),
            .I(N__22930));
    CascadeMux I__4742 (
            .O(N__22930),
            .I(N__22927));
    CascadeBuf I__4741 (
            .O(N__22927),
            .I(N__22924));
    CascadeMux I__4740 (
            .O(N__22924),
            .I(N__22921));
    CascadeBuf I__4739 (
            .O(N__22921),
            .I(N__22918));
    CascadeMux I__4738 (
            .O(N__22918),
            .I(N__22915));
    CascadeBuf I__4737 (
            .O(N__22915),
            .I(N__22912));
    CascadeMux I__4736 (
            .O(N__22912),
            .I(N__22909));
    CascadeBuf I__4735 (
            .O(N__22909),
            .I(N__22906));
    CascadeMux I__4734 (
            .O(N__22906),
            .I(N__22903));
    CascadeBuf I__4733 (
            .O(N__22903),
            .I(N__22900));
    CascadeMux I__4732 (
            .O(N__22900),
            .I(N__22897));
    CascadeBuf I__4731 (
            .O(N__22897),
            .I(N__22894));
    CascadeMux I__4730 (
            .O(N__22894),
            .I(N__22891));
    CascadeBuf I__4729 (
            .O(N__22891),
            .I(N__22888));
    CascadeMux I__4728 (
            .O(N__22888),
            .I(N__22885));
    CascadeBuf I__4727 (
            .O(N__22885),
            .I(N__22882));
    CascadeMux I__4726 (
            .O(N__22882),
            .I(N__22879));
    CascadeBuf I__4725 (
            .O(N__22879),
            .I(N__22876));
    CascadeMux I__4724 (
            .O(N__22876),
            .I(N__22873));
    InMux I__4723 (
            .O(N__22873),
            .I(N__22870));
    LocalMux I__4722 (
            .O(N__22870),
            .I(N__22867));
    Span4Mux_h I__4721 (
            .O(N__22867),
            .I(N__22864));
    Span4Mux_h I__4720 (
            .O(N__22864),
            .I(N__22861));
    Span4Mux_h I__4719 (
            .O(N__22861),
            .I(N__22856));
    InMux I__4718 (
            .O(N__22860),
            .I(N__22852));
    InMux I__4717 (
            .O(N__22859),
            .I(N__22849));
    Sp12to4 I__4716 (
            .O(N__22856),
            .I(N__22846));
    InMux I__4715 (
            .O(N__22855),
            .I(N__22843));
    LocalMux I__4714 (
            .O(N__22852),
            .I(N__22836));
    LocalMux I__4713 (
            .O(N__22849),
            .I(N__22836));
    Span12Mux_s11_v I__4712 (
            .O(N__22846),
            .I(N__22836));
    LocalMux I__4711 (
            .O(N__22843),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv12 I__4710 (
            .O(N__22836),
            .I(M_this_sprites_address_qZ0Z_9));
    InMux I__4709 (
            .O(N__22831),
            .I(N__22828));
    LocalMux I__4708 (
            .O(N__22828),
            .I(N__22825));
    Odrv12 I__4707 (
            .O(N__22825),
            .I(un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0));
    InMux I__4706 (
            .O(N__22822),
            .I(un1_M_this_sprites_address_q_cry_8));
    CascadeMux I__4705 (
            .O(N__22819),
            .I(N__22816));
    CascadeBuf I__4704 (
            .O(N__22816),
            .I(N__22813));
    CascadeMux I__4703 (
            .O(N__22813),
            .I(N__22810));
    CascadeBuf I__4702 (
            .O(N__22810),
            .I(N__22807));
    CascadeMux I__4701 (
            .O(N__22807),
            .I(N__22804));
    CascadeBuf I__4700 (
            .O(N__22804),
            .I(N__22801));
    CascadeMux I__4699 (
            .O(N__22801),
            .I(N__22798));
    CascadeBuf I__4698 (
            .O(N__22798),
            .I(N__22795));
    CascadeMux I__4697 (
            .O(N__22795),
            .I(N__22792));
    CascadeBuf I__4696 (
            .O(N__22792),
            .I(N__22789));
    CascadeMux I__4695 (
            .O(N__22789),
            .I(N__22786));
    CascadeBuf I__4694 (
            .O(N__22786),
            .I(N__22783));
    CascadeMux I__4693 (
            .O(N__22783),
            .I(N__22780));
    CascadeBuf I__4692 (
            .O(N__22780),
            .I(N__22777));
    CascadeMux I__4691 (
            .O(N__22777),
            .I(N__22774));
    CascadeBuf I__4690 (
            .O(N__22774),
            .I(N__22771));
    CascadeMux I__4689 (
            .O(N__22771),
            .I(N__22768));
    CascadeBuf I__4688 (
            .O(N__22768),
            .I(N__22765));
    CascadeMux I__4687 (
            .O(N__22765),
            .I(N__22762));
    CascadeBuf I__4686 (
            .O(N__22762),
            .I(N__22759));
    CascadeMux I__4685 (
            .O(N__22759),
            .I(N__22756));
    CascadeBuf I__4684 (
            .O(N__22756),
            .I(N__22753));
    CascadeMux I__4683 (
            .O(N__22753),
            .I(N__22750));
    CascadeBuf I__4682 (
            .O(N__22750),
            .I(N__22747));
    CascadeMux I__4681 (
            .O(N__22747),
            .I(N__22744));
    CascadeBuf I__4680 (
            .O(N__22744),
            .I(N__22741));
    CascadeMux I__4679 (
            .O(N__22741),
            .I(N__22738));
    CascadeBuf I__4678 (
            .O(N__22738),
            .I(N__22735));
    CascadeMux I__4677 (
            .O(N__22735),
            .I(N__22732));
    CascadeBuf I__4676 (
            .O(N__22732),
            .I(N__22729));
    CascadeMux I__4675 (
            .O(N__22729),
            .I(N__22726));
    InMux I__4674 (
            .O(N__22726),
            .I(N__22723));
    LocalMux I__4673 (
            .O(N__22723),
            .I(N__22720));
    Span4Mux_s2_v I__4672 (
            .O(N__22720),
            .I(N__22716));
    InMux I__4671 (
            .O(N__22719),
            .I(N__22712));
    Span4Mux_v I__4670 (
            .O(N__22716),
            .I(N__22709));
    InMux I__4669 (
            .O(N__22715),
            .I(N__22705));
    LocalMux I__4668 (
            .O(N__22712),
            .I(N__22702));
    Sp12to4 I__4667 (
            .O(N__22709),
            .I(N__22699));
    InMux I__4666 (
            .O(N__22708),
            .I(N__22696));
    LocalMux I__4665 (
            .O(N__22705),
            .I(N__22691));
    Span4Mux_h I__4664 (
            .O(N__22702),
            .I(N__22691));
    Span12Mux_h I__4663 (
            .O(N__22699),
            .I(N__22688));
    LocalMux I__4662 (
            .O(N__22696),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv4 I__4661 (
            .O(N__22691),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv12 I__4660 (
            .O(N__22688),
            .I(M_this_sprites_address_qZ0Z_10));
    InMux I__4659 (
            .O(N__22681),
            .I(N__22678));
    LocalMux I__4658 (
            .O(N__22678),
            .I(un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0));
    InMux I__4657 (
            .O(N__22675),
            .I(un1_M_this_sprites_address_q_cry_9));
    InMux I__4656 (
            .O(N__22672),
            .I(un1_M_this_sprites_address_q_cry_10));
    InMux I__4655 (
            .O(N__22669),
            .I(un1_M_this_sprites_address_q_cry_11));
    InMux I__4654 (
            .O(N__22666),
            .I(un1_M_this_sprites_address_q_cry_12));
    CascadeMux I__4653 (
            .O(N__22663),
            .I(N__22659));
    InMux I__4652 (
            .O(N__22662),
            .I(N__22656));
    InMux I__4651 (
            .O(N__22659),
            .I(N__22650));
    LocalMux I__4650 (
            .O(N__22656),
            .I(N__22647));
    InMux I__4649 (
            .O(N__22655),
            .I(N__22640));
    InMux I__4648 (
            .O(N__22654),
            .I(N__22640));
    InMux I__4647 (
            .O(N__22653),
            .I(N__22640));
    LocalMux I__4646 (
            .O(N__22650),
            .I(N__22637));
    Odrv4 I__4645 (
            .O(N__22647),
            .I(\this_vga_signals.M_this_state_q_ns_15 ));
    LocalMux I__4644 (
            .O(N__22640),
            .I(\this_vga_signals.M_this_state_q_ns_15 ));
    Odrv4 I__4643 (
            .O(N__22637),
            .I(\this_vga_signals.M_this_state_q_ns_15 ));
    InMux I__4642 (
            .O(N__22630),
            .I(N__22627));
    LocalMux I__4641 (
            .O(N__22627),
            .I(N__22624));
    Odrv4 I__4640 (
            .O(N__22624),
            .I(un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0));
    InMux I__4639 (
            .O(N__22621),
            .I(un1_M_this_sprites_address_q_cry_0));
    CascadeMux I__4638 (
            .O(N__22618),
            .I(N__22615));
    CascadeBuf I__4637 (
            .O(N__22615),
            .I(N__22612));
    CascadeMux I__4636 (
            .O(N__22612),
            .I(N__22609));
    CascadeBuf I__4635 (
            .O(N__22609),
            .I(N__22606));
    CascadeMux I__4634 (
            .O(N__22606),
            .I(N__22603));
    CascadeBuf I__4633 (
            .O(N__22603),
            .I(N__22600));
    CascadeMux I__4632 (
            .O(N__22600),
            .I(N__22597));
    CascadeBuf I__4631 (
            .O(N__22597),
            .I(N__22594));
    CascadeMux I__4630 (
            .O(N__22594),
            .I(N__22591));
    CascadeBuf I__4629 (
            .O(N__22591),
            .I(N__22588));
    CascadeMux I__4628 (
            .O(N__22588),
            .I(N__22585));
    CascadeBuf I__4627 (
            .O(N__22585),
            .I(N__22582));
    CascadeMux I__4626 (
            .O(N__22582),
            .I(N__22579));
    CascadeBuf I__4625 (
            .O(N__22579),
            .I(N__22576));
    CascadeMux I__4624 (
            .O(N__22576),
            .I(N__22573));
    CascadeBuf I__4623 (
            .O(N__22573),
            .I(N__22570));
    CascadeMux I__4622 (
            .O(N__22570),
            .I(N__22567));
    CascadeBuf I__4621 (
            .O(N__22567),
            .I(N__22564));
    CascadeMux I__4620 (
            .O(N__22564),
            .I(N__22561));
    CascadeBuf I__4619 (
            .O(N__22561),
            .I(N__22558));
    CascadeMux I__4618 (
            .O(N__22558),
            .I(N__22555));
    CascadeBuf I__4617 (
            .O(N__22555),
            .I(N__22552));
    CascadeMux I__4616 (
            .O(N__22552),
            .I(N__22549));
    CascadeBuf I__4615 (
            .O(N__22549),
            .I(N__22546));
    CascadeMux I__4614 (
            .O(N__22546),
            .I(N__22543));
    CascadeBuf I__4613 (
            .O(N__22543),
            .I(N__22540));
    CascadeMux I__4612 (
            .O(N__22540),
            .I(N__22537));
    CascadeBuf I__4611 (
            .O(N__22537),
            .I(N__22534));
    CascadeMux I__4610 (
            .O(N__22534),
            .I(N__22531));
    CascadeBuf I__4609 (
            .O(N__22531),
            .I(N__22528));
    CascadeMux I__4608 (
            .O(N__22528),
            .I(N__22525));
    InMux I__4607 (
            .O(N__22525),
            .I(N__22522));
    LocalMux I__4606 (
            .O(N__22522),
            .I(N__22519));
    Span4Mux_v I__4605 (
            .O(N__22519),
            .I(N__22516));
    Span4Mux_h I__4604 (
            .O(N__22516),
            .I(N__22512));
    InMux I__4603 (
            .O(N__22515),
            .I(N__22509));
    Sp12to4 I__4602 (
            .O(N__22512),
            .I(N__22504));
    LocalMux I__4601 (
            .O(N__22509),
            .I(N__22501));
    InMux I__4600 (
            .O(N__22508),
            .I(N__22496));
    InMux I__4599 (
            .O(N__22507),
            .I(N__22496));
    Span12Mux_v I__4598 (
            .O(N__22504),
            .I(N__22493));
    Odrv4 I__4597 (
            .O(N__22501),
            .I(M_this_sprites_address_qZ0Z_2));
    LocalMux I__4596 (
            .O(N__22496),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv12 I__4595 (
            .O(N__22493),
            .I(M_this_sprites_address_qZ0Z_2));
    InMux I__4594 (
            .O(N__22486),
            .I(N__22483));
    LocalMux I__4593 (
            .O(N__22483),
            .I(N__22480));
    Odrv4 I__4592 (
            .O(N__22480),
            .I(un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0));
    InMux I__4591 (
            .O(N__22477),
            .I(un1_M_this_sprites_address_q_cry_1));
    InMux I__4590 (
            .O(N__22474),
            .I(N__22471));
    LocalMux I__4589 (
            .O(N__22471),
            .I(N__22468));
    Odrv4 I__4588 (
            .O(N__22468),
            .I(un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0));
    InMux I__4587 (
            .O(N__22465),
            .I(un1_M_this_sprites_address_q_cry_2));
    InMux I__4586 (
            .O(N__22462),
            .I(un1_M_this_sprites_address_q_cry_3));
    InMux I__4585 (
            .O(N__22459),
            .I(un1_M_this_sprites_address_q_cry_4));
    CascadeMux I__4584 (
            .O(N__22456),
            .I(N__22453));
    InMux I__4583 (
            .O(N__22453),
            .I(N__22450));
    LocalMux I__4582 (
            .O(N__22450),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_1 ));
    InMux I__4581 (
            .O(N__22447),
            .I(N__22444));
    LocalMux I__4580 (
            .O(N__22444),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9 ));
    CascadeMux I__4579 (
            .O(N__22441),
            .I(N__22438));
    InMux I__4578 (
            .O(N__22438),
            .I(N__22435));
    LocalMux I__4577 (
            .O(N__22435),
            .I(N__22432));
    Odrv4 I__4576 (
            .O(N__22432),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_9 ));
    CascadeMux I__4575 (
            .O(N__22429),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2_cascade_ ));
    InMux I__4574 (
            .O(N__22426),
            .I(N__22423));
    LocalMux I__4573 (
            .O(N__22423),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_2 ));
    CascadeMux I__4572 (
            .O(N__22420),
            .I(N__22417));
    InMux I__4571 (
            .O(N__22417),
            .I(N__22414));
    LocalMux I__4570 (
            .O(N__22414),
            .I(N__22411));
    Odrv4 I__4569 (
            .O(N__22411),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_3 ));
    CascadeMux I__4568 (
            .O(N__22408),
            .I(N__22405));
    InMux I__4567 (
            .O(N__22405),
            .I(N__22402));
    LocalMux I__4566 (
            .O(N__22402),
            .I(N__22399));
    Span4Mux_v I__4565 (
            .O(N__22399),
            .I(N__22396));
    Odrv4 I__4564 (
            .O(N__22396),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_10 ));
    InMux I__4563 (
            .O(N__22393),
            .I(N__22390));
    LocalMux I__4562 (
            .O(N__22390),
            .I(M_this_state_q_RNIMJ231Z0Z_8));
    CascadeMux I__4561 (
            .O(N__22387),
            .I(N__22384));
    InMux I__4560 (
            .O(N__22384),
            .I(N__22381));
    LocalMux I__4559 (
            .O(N__22381),
            .I(\this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_3 ));
    InMux I__4558 (
            .O(N__22378),
            .I(N__22375));
    LocalMux I__4557 (
            .O(N__22375),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10 ));
    CascadeMux I__4556 (
            .O(N__22372),
            .I(N__22369));
    CascadeBuf I__4555 (
            .O(N__22369),
            .I(N__22366));
    CascadeMux I__4554 (
            .O(N__22366),
            .I(N__22363));
    CascadeBuf I__4553 (
            .O(N__22363),
            .I(N__22360));
    CascadeMux I__4552 (
            .O(N__22360),
            .I(N__22357));
    CascadeBuf I__4551 (
            .O(N__22357),
            .I(N__22354));
    CascadeMux I__4550 (
            .O(N__22354),
            .I(N__22351));
    CascadeBuf I__4549 (
            .O(N__22351),
            .I(N__22348));
    CascadeMux I__4548 (
            .O(N__22348),
            .I(N__22345));
    CascadeBuf I__4547 (
            .O(N__22345),
            .I(N__22342));
    CascadeMux I__4546 (
            .O(N__22342),
            .I(N__22339));
    CascadeBuf I__4545 (
            .O(N__22339),
            .I(N__22336));
    CascadeMux I__4544 (
            .O(N__22336),
            .I(N__22333));
    CascadeBuf I__4543 (
            .O(N__22333),
            .I(N__22330));
    CascadeMux I__4542 (
            .O(N__22330),
            .I(N__22327));
    CascadeBuf I__4541 (
            .O(N__22327),
            .I(N__22324));
    CascadeMux I__4540 (
            .O(N__22324),
            .I(N__22321));
    CascadeBuf I__4539 (
            .O(N__22321),
            .I(N__22318));
    CascadeMux I__4538 (
            .O(N__22318),
            .I(N__22315));
    CascadeBuf I__4537 (
            .O(N__22315),
            .I(N__22312));
    CascadeMux I__4536 (
            .O(N__22312),
            .I(N__22309));
    CascadeBuf I__4535 (
            .O(N__22309),
            .I(N__22306));
    CascadeMux I__4534 (
            .O(N__22306),
            .I(N__22303));
    CascadeBuf I__4533 (
            .O(N__22303),
            .I(N__22300));
    CascadeMux I__4532 (
            .O(N__22300),
            .I(N__22297));
    CascadeBuf I__4531 (
            .O(N__22297),
            .I(N__22294));
    CascadeMux I__4530 (
            .O(N__22294),
            .I(N__22291));
    CascadeBuf I__4529 (
            .O(N__22291),
            .I(N__22288));
    CascadeMux I__4528 (
            .O(N__22288),
            .I(N__22285));
    CascadeBuf I__4527 (
            .O(N__22285),
            .I(N__22281));
    CascadeMux I__4526 (
            .O(N__22284),
            .I(N__22278));
    CascadeMux I__4525 (
            .O(N__22281),
            .I(N__22275));
    InMux I__4524 (
            .O(N__22278),
            .I(N__22272));
    InMux I__4523 (
            .O(N__22275),
            .I(N__22269));
    LocalMux I__4522 (
            .O(N__22272),
            .I(N__22266));
    LocalMux I__4521 (
            .O(N__22269),
            .I(N__22263));
    Span4Mux_v I__4520 (
            .O(N__22266),
            .I(N__22259));
    Span4Mux_v I__4519 (
            .O(N__22263),
            .I(N__22256));
    InMux I__4518 (
            .O(N__22262),
            .I(N__22253));
    Sp12to4 I__4517 (
            .O(N__22259),
            .I(N__22248));
    Sp12to4 I__4516 (
            .O(N__22256),
            .I(N__22245));
    LocalMux I__4515 (
            .O(N__22253),
            .I(N__22242));
    InMux I__4514 (
            .O(N__22252),
            .I(N__22237));
    InMux I__4513 (
            .O(N__22251),
            .I(N__22237));
    Span12Mux_h I__4512 (
            .O(N__22248),
            .I(N__22232));
    Span12Mux_h I__4511 (
            .O(N__22245),
            .I(N__22232));
    Odrv4 I__4510 (
            .O(N__22242),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__4509 (
            .O(N__22237),
            .I(M_this_ppu_vram_addr_0));
    Odrv12 I__4508 (
            .O(N__22232),
            .I(M_this_ppu_vram_addr_0));
    CEMux I__4507 (
            .O(N__22225),
            .I(N__22221));
    InMux I__4506 (
            .O(N__22224),
            .I(N__22216));
    LocalMux I__4505 (
            .O(N__22221),
            .I(N__22213));
    InMux I__4504 (
            .O(N__22220),
            .I(N__22210));
    InMux I__4503 (
            .O(N__22219),
            .I(N__22207));
    LocalMux I__4502 (
            .O(N__22216),
            .I(N__22204));
    Span4Mux_h I__4501 (
            .O(N__22213),
            .I(N__22201));
    LocalMux I__4500 (
            .O(N__22210),
            .I(N__22196));
    LocalMux I__4499 (
            .O(N__22207),
            .I(N__22196));
    Span4Mux_h I__4498 (
            .O(N__22204),
            .I(N__22193));
    Span4Mux_h I__4497 (
            .O(N__22201),
            .I(N__22190));
    Span4Mux_v I__4496 (
            .O(N__22196),
            .I(N__22187));
    Span4Mux_v I__4495 (
            .O(N__22193),
            .I(N__22184));
    Odrv4 I__4494 (
            .O(N__22190),
            .I(M_this_ppu_vram_en_0));
    Odrv4 I__4493 (
            .O(N__22187),
            .I(M_this_ppu_vram_en_0));
    Odrv4 I__4492 (
            .O(N__22184),
            .I(M_this_ppu_vram_en_0));
    CascadeMux I__4491 (
            .O(N__22177),
            .I(N__22174));
    CascadeBuf I__4490 (
            .O(N__22174),
            .I(N__22171));
    CascadeMux I__4489 (
            .O(N__22171),
            .I(N__22168));
    CascadeBuf I__4488 (
            .O(N__22168),
            .I(N__22165));
    CascadeMux I__4487 (
            .O(N__22165),
            .I(N__22162));
    CascadeBuf I__4486 (
            .O(N__22162),
            .I(N__22159));
    CascadeMux I__4485 (
            .O(N__22159),
            .I(N__22156));
    CascadeBuf I__4484 (
            .O(N__22156),
            .I(N__22153));
    CascadeMux I__4483 (
            .O(N__22153),
            .I(N__22150));
    CascadeBuf I__4482 (
            .O(N__22150),
            .I(N__22147));
    CascadeMux I__4481 (
            .O(N__22147),
            .I(N__22144));
    CascadeBuf I__4480 (
            .O(N__22144),
            .I(N__22141));
    CascadeMux I__4479 (
            .O(N__22141),
            .I(N__22138));
    CascadeBuf I__4478 (
            .O(N__22138),
            .I(N__22135));
    CascadeMux I__4477 (
            .O(N__22135),
            .I(N__22132));
    CascadeBuf I__4476 (
            .O(N__22132),
            .I(N__22129));
    CascadeMux I__4475 (
            .O(N__22129),
            .I(N__22126));
    CascadeBuf I__4474 (
            .O(N__22126),
            .I(N__22123));
    CascadeMux I__4473 (
            .O(N__22123),
            .I(N__22120));
    CascadeBuf I__4472 (
            .O(N__22120),
            .I(N__22117));
    CascadeMux I__4471 (
            .O(N__22117),
            .I(N__22114));
    CascadeBuf I__4470 (
            .O(N__22114),
            .I(N__22111));
    CascadeMux I__4469 (
            .O(N__22111),
            .I(N__22108));
    CascadeBuf I__4468 (
            .O(N__22108),
            .I(N__22105));
    CascadeMux I__4467 (
            .O(N__22105),
            .I(N__22102));
    CascadeBuf I__4466 (
            .O(N__22102),
            .I(N__22099));
    CascadeMux I__4465 (
            .O(N__22099),
            .I(N__22096));
    CascadeBuf I__4464 (
            .O(N__22096),
            .I(N__22093));
    CascadeMux I__4463 (
            .O(N__22093),
            .I(N__22090));
    CascadeBuf I__4462 (
            .O(N__22090),
            .I(N__22087));
    CascadeMux I__4461 (
            .O(N__22087),
            .I(N__22083));
    CascadeMux I__4460 (
            .O(N__22086),
            .I(N__22080));
    InMux I__4459 (
            .O(N__22083),
            .I(N__22077));
    InMux I__4458 (
            .O(N__22080),
            .I(N__22073));
    LocalMux I__4457 (
            .O(N__22077),
            .I(N__22070));
    CascadeMux I__4456 (
            .O(N__22076),
            .I(N__22067));
    LocalMux I__4455 (
            .O(N__22073),
            .I(N__22063));
    Span4Mux_s3_v I__4454 (
            .O(N__22070),
            .I(N__22060));
    InMux I__4453 (
            .O(N__22067),
            .I(N__22057));
    CascadeMux I__4452 (
            .O(N__22066),
            .I(N__22054));
    Sp12to4 I__4451 (
            .O(N__22063),
            .I(N__22051));
    Sp12to4 I__4450 (
            .O(N__22060),
            .I(N__22048));
    LocalMux I__4449 (
            .O(N__22057),
            .I(N__22045));
    InMux I__4448 (
            .O(N__22054),
            .I(N__22042));
    Span12Mux_v I__4447 (
            .O(N__22051),
            .I(N__22039));
    Span12Mux_h I__4446 (
            .O(N__22048),
            .I(N__22036));
    Odrv4 I__4445 (
            .O(N__22045),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__4444 (
            .O(N__22042),
            .I(M_this_ppu_vram_addr_1));
    Odrv12 I__4443 (
            .O(N__22039),
            .I(M_this_ppu_vram_addr_1));
    Odrv12 I__4442 (
            .O(N__22036),
            .I(M_this_ppu_vram_addr_1));
    InMux I__4441 (
            .O(N__22027),
            .I(N__22017));
    InMux I__4440 (
            .O(N__22026),
            .I(N__22017));
    InMux I__4439 (
            .O(N__22025),
            .I(N__22012));
    InMux I__4438 (
            .O(N__22024),
            .I(N__22012));
    InMux I__4437 (
            .O(N__22023),
            .I(N__22005));
    InMux I__4436 (
            .O(N__22022),
            .I(N__22002));
    LocalMux I__4435 (
            .O(N__22017),
            .I(N__21998));
    LocalMux I__4434 (
            .O(N__22012),
            .I(N__21995));
    CascadeMux I__4433 (
            .O(N__22011),
            .I(N__21991));
    InMux I__4432 (
            .O(N__22010),
            .I(N__21984));
    InMux I__4431 (
            .O(N__22009),
            .I(N__21979));
    InMux I__4430 (
            .O(N__22008),
            .I(N__21979));
    LocalMux I__4429 (
            .O(N__22005),
            .I(N__21976));
    LocalMux I__4428 (
            .O(N__22002),
            .I(N__21973));
    InMux I__4427 (
            .O(N__22001),
            .I(N__21969));
    Span4Mux_v I__4426 (
            .O(N__21998),
            .I(N__21964));
    Span4Mux_v I__4425 (
            .O(N__21995),
            .I(N__21964));
    InMux I__4424 (
            .O(N__21994),
            .I(N__21961));
    InMux I__4423 (
            .O(N__21991),
            .I(N__21958));
    InMux I__4422 (
            .O(N__21990),
            .I(N__21955));
    InMux I__4421 (
            .O(N__21989),
            .I(N__21948));
    InMux I__4420 (
            .O(N__21988),
            .I(N__21948));
    InMux I__4419 (
            .O(N__21987),
            .I(N__21948));
    LocalMux I__4418 (
            .O(N__21984),
            .I(N__21945));
    LocalMux I__4417 (
            .O(N__21979),
            .I(N__21940));
    Span4Mux_v I__4416 (
            .O(N__21976),
            .I(N__21940));
    Span4Mux_v I__4415 (
            .O(N__21973),
            .I(N__21937));
    InMux I__4414 (
            .O(N__21972),
            .I(N__21934));
    LocalMux I__4413 (
            .O(N__21969),
            .I(N__21929));
    Span4Mux_h I__4412 (
            .O(N__21964),
            .I(N__21929));
    LocalMux I__4411 (
            .O(N__21961),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    LocalMux I__4410 (
            .O(N__21958),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    LocalMux I__4409 (
            .O(N__21955),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    LocalMux I__4408 (
            .O(N__21948),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    Odrv4 I__4407 (
            .O(N__21945),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    Odrv4 I__4406 (
            .O(N__21940),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    Odrv4 I__4405 (
            .O(N__21937),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    LocalMux I__4404 (
            .O(N__21934),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    Odrv4 I__4403 (
            .O(N__21929),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    InMux I__4402 (
            .O(N__21910),
            .I(N__21907));
    LocalMux I__4401 (
            .O(N__21907),
            .I(N__21904));
    Odrv4 I__4400 (
            .O(N__21904),
            .I(M_this_state_q_RNI2S2SZ0Z_13));
    CascadeMux I__4399 (
            .O(N__21901),
            .I(M_this_state_q_RNITS9I4Z0Z_7_cascade_));
    IoInMux I__4398 (
            .O(N__21898),
            .I(N__21895));
    LocalMux I__4397 (
            .O(N__21895),
            .I(N__21892));
    IoSpan4Mux I__4396 (
            .O(N__21892),
            .I(N__21889));
    Span4Mux_s3_h I__4395 (
            .O(N__21889),
            .I(N__21886));
    Sp12to4 I__4394 (
            .O(N__21886),
            .I(N__21883));
    Span12Mux_s11_h I__4393 (
            .O(N__21883),
            .I(N__21880));
    Span12Mux_v I__4392 (
            .O(N__21880),
            .I(N__21877));
    Odrv12 I__4391 (
            .O(N__21877),
            .I(dma_ac0_5_i));
    CascadeMux I__4390 (
            .O(N__21874),
            .I(dma_ac0_5_i_cascade_));
    IoInMux I__4389 (
            .O(N__21871),
            .I(N__21868));
    LocalMux I__4388 (
            .O(N__21868),
            .I(N__21862));
    IoInMux I__4387 (
            .O(N__21867),
            .I(N__21859));
    IoInMux I__4386 (
            .O(N__21866),
            .I(N__21855));
    IoInMux I__4385 (
            .O(N__21865),
            .I(N__21849));
    IoSpan4Mux I__4384 (
            .O(N__21862),
            .I(N__21843));
    LocalMux I__4383 (
            .O(N__21859),
            .I(N__21843));
    IoInMux I__4382 (
            .O(N__21858),
            .I(N__21840));
    LocalMux I__4381 (
            .O(N__21855),
            .I(N__21836));
    IoInMux I__4380 (
            .O(N__21854),
            .I(N__21833));
    IoInMux I__4379 (
            .O(N__21853),
            .I(N__21830));
    IoInMux I__4378 (
            .O(N__21852),
            .I(N__21827));
    LocalMux I__4377 (
            .O(N__21849),
            .I(N__21823));
    IoInMux I__4376 (
            .O(N__21848),
            .I(N__21819));
    IoSpan4Mux I__4375 (
            .O(N__21843),
            .I(N__21814));
    LocalMux I__4374 (
            .O(N__21840),
            .I(N__21814));
    IoInMux I__4373 (
            .O(N__21839),
            .I(N__21811));
    IoSpan4Mux I__4372 (
            .O(N__21836),
            .I(N__21802));
    LocalMux I__4371 (
            .O(N__21833),
            .I(N__21802));
    LocalMux I__4370 (
            .O(N__21830),
            .I(N__21802));
    LocalMux I__4369 (
            .O(N__21827),
            .I(N__21799));
    IoInMux I__4368 (
            .O(N__21826),
            .I(N__21796));
    IoSpan4Mux I__4367 (
            .O(N__21823),
            .I(N__21793));
    IoInMux I__4366 (
            .O(N__21822),
            .I(N__21790));
    LocalMux I__4365 (
            .O(N__21819),
            .I(N__21787));
    IoSpan4Mux I__4364 (
            .O(N__21814),
            .I(N__21782));
    LocalMux I__4363 (
            .O(N__21811),
            .I(N__21782));
    IoInMux I__4362 (
            .O(N__21810),
            .I(N__21779));
    IoInMux I__4361 (
            .O(N__21809),
            .I(N__21776));
    IoSpan4Mux I__4360 (
            .O(N__21802),
            .I(N__21768));
    IoSpan4Mux I__4359 (
            .O(N__21799),
            .I(N__21768));
    LocalMux I__4358 (
            .O(N__21796),
            .I(N__21768));
    IoSpan4Mux I__4357 (
            .O(N__21793),
            .I(N__21763));
    LocalMux I__4356 (
            .O(N__21790),
            .I(N__21763));
    IoSpan4Mux I__4355 (
            .O(N__21787),
            .I(N__21760));
    IoSpan4Mux I__4354 (
            .O(N__21782),
            .I(N__21755));
    LocalMux I__4353 (
            .O(N__21779),
            .I(N__21755));
    LocalMux I__4352 (
            .O(N__21776),
            .I(N__21752));
    IoInMux I__4351 (
            .O(N__21775),
            .I(N__21749));
    IoSpan4Mux I__4350 (
            .O(N__21768),
            .I(N__21744));
    IoSpan4Mux I__4349 (
            .O(N__21763),
            .I(N__21744));
    Span4Mux_s3_h I__4348 (
            .O(N__21760),
            .I(N__21740));
    IoSpan4Mux I__4347 (
            .O(N__21755),
            .I(N__21735));
    IoSpan4Mux I__4346 (
            .O(N__21752),
            .I(N__21735));
    LocalMux I__4345 (
            .O(N__21749),
            .I(N__21731));
    Span4Mux_s0_h I__4344 (
            .O(N__21744),
            .I(N__21728));
    IoInMux I__4343 (
            .O(N__21743),
            .I(N__21725));
    Span4Mux_v I__4342 (
            .O(N__21740),
            .I(N__21722));
    Span4Mux_s3_v I__4341 (
            .O(N__21735),
            .I(N__21719));
    IoInMux I__4340 (
            .O(N__21734),
            .I(N__21716));
    Span12Mux_s9_h I__4339 (
            .O(N__21731),
            .I(N__21713));
    Sp12to4 I__4338 (
            .O(N__21728),
            .I(N__21708));
    LocalMux I__4337 (
            .O(N__21725),
            .I(N__21708));
    Sp12to4 I__4336 (
            .O(N__21722),
            .I(N__21705));
    Sp12to4 I__4335 (
            .O(N__21719),
            .I(N__21700));
    LocalMux I__4334 (
            .O(N__21716),
            .I(N__21700));
    Span12Mux_v I__4333 (
            .O(N__21713),
            .I(N__21695));
    Span12Mux_s9_h I__4332 (
            .O(N__21708),
            .I(N__21695));
    Span12Mux_h I__4331 (
            .O(N__21705),
            .I(N__21690));
    Span12Mux_s5_v I__4330 (
            .O(N__21700),
            .I(N__21690));
    Odrv12 I__4329 (
            .O(N__21695),
            .I(dma_ac0_5_i_i));
    Odrv12 I__4328 (
            .O(N__21690),
            .I(dma_ac0_5_i_i));
    InMux I__4327 (
            .O(N__21685),
            .I(N__21682));
    LocalMux I__4326 (
            .O(N__21682),
            .I(\this_vga_signals.un23_i_a2_4Z0Z_0 ));
    InMux I__4325 (
            .O(N__21679),
            .I(N__21676));
    LocalMux I__4324 (
            .O(N__21676),
            .I(M_this_state_q_RNI6Q0SZ0Z_7));
    InMux I__4323 (
            .O(N__21673),
            .I(N__21670));
    LocalMux I__4322 (
            .O(N__21670),
            .I(N__21667));
    Odrv4 I__4321 (
            .O(N__21667),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8 ));
    CascadeMux I__4320 (
            .O(N__21664),
            .I(N__21661));
    InMux I__4319 (
            .O(N__21661),
            .I(N__21658));
    LocalMux I__4318 (
            .O(N__21658),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_8 ));
    CascadeMux I__4317 (
            .O(N__21655),
            .I(\this_vga_signals.un23_i_a2_x1Z0Z_0_cascade_ ));
    InMux I__4316 (
            .O(N__21652),
            .I(N__21649));
    LocalMux I__4315 (
            .O(N__21649),
            .I(N__21646));
    Span4Mux_v I__4314 (
            .O(N__21646),
            .I(N__21643));
    Span4Mux_v I__4313 (
            .O(N__21643),
            .I(N__21638));
    InMux I__4312 (
            .O(N__21642),
            .I(N__21635));
    InMux I__4311 (
            .O(N__21641),
            .I(N__21632));
    Sp12to4 I__4310 (
            .O(N__21638),
            .I(N__21627));
    LocalMux I__4309 (
            .O(N__21635),
            .I(N__21627));
    LocalMux I__4308 (
            .O(N__21632),
            .I(N__21624));
    Span12Mux_s4_h I__4307 (
            .O(N__21627),
            .I(N__21621));
    Span4Mux_v I__4306 (
            .O(N__21624),
            .I(N__21618));
    Span12Mux_h I__4305 (
            .O(N__21621),
            .I(N__21615));
    Span4Mux_h I__4304 (
            .O(N__21618),
            .I(N__21612));
    Odrv12 I__4303 (
            .O(N__21615),
            .I(dma_ac0Z0Z_5));
    Odrv4 I__4302 (
            .O(N__21612),
            .I(dma_ac0Z0Z_5));
    InMux I__4301 (
            .O(N__21607),
            .I(N__21604));
    LocalMux I__4300 (
            .O(N__21604),
            .I(this_vga_signals_un23_i_a2_1_3));
    InMux I__4299 (
            .O(N__21601),
            .I(N__21598));
    LocalMux I__4298 (
            .O(N__21598),
            .I(this_vga_signals_un23_i_a2_4_2));
    CascadeMux I__4297 (
            .O(N__21595),
            .I(this_vga_signals_un23_i_a2_3_2_cascade_));
    InMux I__4296 (
            .O(N__21592),
            .I(N__21589));
    LocalMux I__4295 (
            .O(N__21589),
            .I(dma_c3_0));
    InMux I__4294 (
            .O(N__21586),
            .I(N__21582));
    InMux I__4293 (
            .O(N__21585),
            .I(N__21579));
    LocalMux I__4292 (
            .O(N__21582),
            .I(dma_axb0));
    LocalMux I__4291 (
            .O(N__21579),
            .I(dma_axb0));
    CascadeMux I__4290 (
            .O(N__21574),
            .I(N__21571));
    CascadeBuf I__4289 (
            .O(N__21571),
            .I(N__21568));
    CascadeMux I__4288 (
            .O(N__21568),
            .I(N__21565));
    InMux I__4287 (
            .O(N__21565),
            .I(N__21562));
    LocalMux I__4286 (
            .O(N__21562),
            .I(N__21559));
    Span4Mux_s2_v I__4285 (
            .O(N__21559),
            .I(N__21556));
    Span4Mux_h I__4284 (
            .O(N__21556),
            .I(N__21552));
    CascadeMux I__4283 (
            .O(N__21555),
            .I(N__21548));
    Span4Mux_h I__4282 (
            .O(N__21552),
            .I(N__21544));
    InMux I__4281 (
            .O(N__21551),
            .I(N__21541));
    InMux I__4280 (
            .O(N__21548),
            .I(N__21538));
    InMux I__4279 (
            .O(N__21547),
            .I(N__21535));
    Span4Mux_v I__4278 (
            .O(N__21544),
            .I(N__21532));
    LocalMux I__4277 (
            .O(N__21541),
            .I(M_this_ppu_map_addr_7));
    LocalMux I__4276 (
            .O(N__21538),
            .I(M_this_ppu_map_addr_7));
    LocalMux I__4275 (
            .O(N__21535),
            .I(M_this_ppu_map_addr_7));
    Odrv4 I__4274 (
            .O(N__21532),
            .I(M_this_ppu_map_addr_7));
    InMux I__4273 (
            .O(N__21523),
            .I(N__21518));
    InMux I__4272 (
            .O(N__21522),
            .I(N__21515));
    InMux I__4271 (
            .O(N__21521),
            .I(N__21512));
    LocalMux I__4270 (
            .O(N__21518),
            .I(\this_ppu.un1_M_vaddress_q_c5 ));
    LocalMux I__4269 (
            .O(N__21515),
            .I(\this_ppu.un1_M_vaddress_q_c5 ));
    LocalMux I__4268 (
            .O(N__21512),
            .I(\this_ppu.un1_M_vaddress_q_c5 ));
    SRMux I__4267 (
            .O(N__21505),
            .I(N__21500));
    SRMux I__4266 (
            .O(N__21504),
            .I(N__21497));
    SRMux I__4265 (
            .O(N__21503),
            .I(N__21494));
    LocalMux I__4264 (
            .O(N__21500),
            .I(N__21489));
    LocalMux I__4263 (
            .O(N__21497),
            .I(N__21484));
    LocalMux I__4262 (
            .O(N__21494),
            .I(N__21484));
    SRMux I__4261 (
            .O(N__21493),
            .I(N__21481));
    SRMux I__4260 (
            .O(N__21492),
            .I(N__21478));
    Span4Mux_h I__4259 (
            .O(N__21489),
            .I(N__21471));
    Span4Mux_v I__4258 (
            .O(N__21484),
            .I(N__21471));
    LocalMux I__4257 (
            .O(N__21481),
            .I(N__21471));
    LocalMux I__4256 (
            .O(N__21478),
            .I(N__21468));
    Span4Mux_h I__4255 (
            .O(N__21471),
            .I(N__21463));
    Span4Mux_v I__4254 (
            .O(N__21468),
            .I(N__21460));
    SRMux I__4253 (
            .O(N__21467),
            .I(N__21457));
    SRMux I__4252 (
            .O(N__21466),
            .I(N__21454));
    Odrv4 I__4251 (
            .O(N__21463),
            .I(\this_ppu.M_last_q_RNIQKTIG ));
    Odrv4 I__4250 (
            .O(N__21460),
            .I(\this_ppu.M_last_q_RNIQKTIG ));
    LocalMux I__4249 (
            .O(N__21457),
            .I(\this_ppu.M_last_q_RNIQKTIG ));
    LocalMux I__4248 (
            .O(N__21454),
            .I(\this_ppu.M_last_q_RNIQKTIG ));
    InMux I__4247 (
            .O(N__21445),
            .I(N__21441));
    InMux I__4246 (
            .O(N__21444),
            .I(N__21438));
    LocalMux I__4245 (
            .O(N__21441),
            .I(\this_ppu.M_vaddress_qZ0Z_7 ));
    LocalMux I__4244 (
            .O(N__21438),
            .I(\this_ppu.M_vaddress_qZ0Z_7 ));
    CascadeMux I__4243 (
            .O(N__21433),
            .I(N__21430));
    CascadeBuf I__4242 (
            .O(N__21430),
            .I(N__21427));
    CascadeMux I__4241 (
            .O(N__21427),
            .I(N__21424));
    InMux I__4240 (
            .O(N__21424),
            .I(N__21421));
    LocalMux I__4239 (
            .O(N__21421),
            .I(N__21418));
    Span12Mux_h I__4238 (
            .O(N__21418),
            .I(N__21415));
    Odrv12 I__4237 (
            .O(N__21415),
            .I(M_this_ppu_map_addr_9));
    IoInMux I__4236 (
            .O(N__21412),
            .I(N__21409));
    LocalMux I__4235 (
            .O(N__21409),
            .I(N__21406));
    IoSpan4Mux I__4234 (
            .O(N__21406),
            .I(N__21403));
    Span4Mux_s0_v I__4233 (
            .O(N__21403),
            .I(N__21400));
    Span4Mux_v I__4232 (
            .O(N__21400),
            .I(N__21397));
    Span4Mux_v I__4231 (
            .O(N__21397),
            .I(N__21394));
    Sp12to4 I__4230 (
            .O(N__21394),
            .I(N__21391));
    Odrv12 I__4229 (
            .O(N__21391),
            .I(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO));
    InMux I__4228 (
            .O(N__21388),
            .I(N__21384));
    InMux I__4227 (
            .O(N__21387),
            .I(N__21380));
    LocalMux I__4226 (
            .O(N__21384),
            .I(N__21376));
    InMux I__4225 (
            .O(N__21383),
            .I(N__21373));
    LocalMux I__4224 (
            .O(N__21380),
            .I(N__21369));
    InMux I__4223 (
            .O(N__21379),
            .I(N__21366));
    Span4Mux_h I__4222 (
            .O(N__21376),
            .I(N__21362));
    LocalMux I__4221 (
            .O(N__21373),
            .I(N__21359));
    InMux I__4220 (
            .O(N__21372),
            .I(N__21356));
    Span4Mux_v I__4219 (
            .O(N__21369),
            .I(N__21350));
    LocalMux I__4218 (
            .O(N__21366),
            .I(N__21350));
    InMux I__4217 (
            .O(N__21365),
            .I(N__21347));
    Span4Mux_v I__4216 (
            .O(N__21362),
            .I(N__21341));
    Span4Mux_h I__4215 (
            .O(N__21359),
            .I(N__21341));
    LocalMux I__4214 (
            .O(N__21356),
            .I(N__21338));
    InMux I__4213 (
            .O(N__21355),
            .I(N__21335));
    Span4Mux_v I__4212 (
            .O(N__21350),
            .I(N__21330));
    LocalMux I__4211 (
            .O(N__21347),
            .I(N__21330));
    InMux I__4210 (
            .O(N__21346),
            .I(N__21327));
    Span4Mux_v I__4209 (
            .O(N__21341),
            .I(N__21322));
    Span4Mux_h I__4208 (
            .O(N__21338),
            .I(N__21322));
    LocalMux I__4207 (
            .O(N__21335),
            .I(N__21319));
    Span4Mux_v I__4206 (
            .O(N__21330),
            .I(N__21314));
    LocalMux I__4205 (
            .O(N__21327),
            .I(N__21314));
    Span4Mux_v I__4204 (
            .O(N__21322),
            .I(N__21309));
    Span4Mux_h I__4203 (
            .O(N__21319),
            .I(N__21309));
    Span4Mux_h I__4202 (
            .O(N__21314),
            .I(N__21306));
    Span4Mux_h I__4201 (
            .O(N__21309),
            .I(N__21301));
    Span4Mux_h I__4200 (
            .O(N__21306),
            .I(N__21301));
    Odrv4 I__4199 (
            .O(N__21301),
            .I(M_this_sprites_ram_write_data_0));
    InMux I__4198 (
            .O(N__21298),
            .I(N__21294));
    InMux I__4197 (
            .O(N__21297),
            .I(N__21290));
    LocalMux I__4196 (
            .O(N__21294),
            .I(N__21286));
    InMux I__4195 (
            .O(N__21293),
            .I(N__21283));
    LocalMux I__4194 (
            .O(N__21290),
            .I(N__21279));
    InMux I__4193 (
            .O(N__21289),
            .I(N__21276));
    Span4Mux_v I__4192 (
            .O(N__21286),
            .I(N__21270));
    LocalMux I__4191 (
            .O(N__21283),
            .I(N__21270));
    InMux I__4190 (
            .O(N__21282),
            .I(N__21267));
    Span4Mux_h I__4189 (
            .O(N__21279),
            .I(N__21264));
    LocalMux I__4188 (
            .O(N__21276),
            .I(N__21261));
    InMux I__4187 (
            .O(N__21275),
            .I(N__21258));
    Span4Mux_v I__4186 (
            .O(N__21270),
            .I(N__21253));
    LocalMux I__4185 (
            .O(N__21267),
            .I(N__21253));
    Span4Mux_v I__4184 (
            .O(N__21264),
            .I(N__21247));
    Span4Mux_h I__4183 (
            .O(N__21261),
            .I(N__21247));
    LocalMux I__4182 (
            .O(N__21258),
            .I(N__21244));
    Span4Mux_v I__4181 (
            .O(N__21253),
            .I(N__21241));
    InMux I__4180 (
            .O(N__21252),
            .I(N__21238));
    Span4Mux_v I__4179 (
            .O(N__21247),
            .I(N__21232));
    Span4Mux_h I__4178 (
            .O(N__21244),
            .I(N__21232));
    Span4Mux_v I__4177 (
            .O(N__21241),
            .I(N__21227));
    LocalMux I__4176 (
            .O(N__21238),
            .I(N__21227));
    InMux I__4175 (
            .O(N__21237),
            .I(N__21224));
    Span4Mux_v I__4174 (
            .O(N__21232),
            .I(N__21219));
    Span4Mux_h I__4173 (
            .O(N__21227),
            .I(N__21219));
    LocalMux I__4172 (
            .O(N__21224),
            .I(N__21216));
    Span4Mux_h I__4171 (
            .O(N__21219),
            .I(N__21213));
    Span12Mux_s10_h I__4170 (
            .O(N__21216),
            .I(N__21210));
    Odrv4 I__4169 (
            .O(N__21213),
            .I(M_this_sprites_ram_write_data_1));
    Odrv12 I__4168 (
            .O(N__21210),
            .I(M_this_sprites_ram_write_data_1));
    CascadeMux I__4167 (
            .O(N__21205),
            .I(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux_cascade_ ));
    InMux I__4166 (
            .O(N__21202),
            .I(N__21199));
    LocalMux I__4165 (
            .O(N__21199),
            .I(N__21192));
    InMux I__4164 (
            .O(N__21198),
            .I(N__21189));
    InMux I__4163 (
            .O(N__21197),
            .I(N__21186));
    InMux I__4162 (
            .O(N__21196),
            .I(N__21183));
    InMux I__4161 (
            .O(N__21195),
            .I(N__21178));
    Span4Mux_v I__4160 (
            .O(N__21192),
            .I(N__21174));
    LocalMux I__4159 (
            .O(N__21189),
            .I(N__21171));
    LocalMux I__4158 (
            .O(N__21186),
            .I(N__21168));
    LocalMux I__4157 (
            .O(N__21183),
            .I(N__21165));
    InMux I__4156 (
            .O(N__21182),
            .I(N__21162));
    InMux I__4155 (
            .O(N__21181),
            .I(N__21159));
    LocalMux I__4154 (
            .O(N__21178),
            .I(N__21156));
    InMux I__4153 (
            .O(N__21177),
            .I(N__21153));
    Sp12to4 I__4152 (
            .O(N__21174),
            .I(N__21146));
    Sp12to4 I__4151 (
            .O(N__21171),
            .I(N__21146));
    Sp12to4 I__4150 (
            .O(N__21168),
            .I(N__21146));
    Sp12to4 I__4149 (
            .O(N__21165),
            .I(N__21143));
    LocalMux I__4148 (
            .O(N__21162),
            .I(N__21140));
    LocalMux I__4147 (
            .O(N__21159),
            .I(N__21137));
    Span12Mux_h I__4146 (
            .O(N__21156),
            .I(N__21134));
    LocalMux I__4145 (
            .O(N__21153),
            .I(N__21131));
    Span12Mux_v I__4144 (
            .O(N__21146),
            .I(N__21126));
    Span12Mux_v I__4143 (
            .O(N__21143),
            .I(N__21126));
    Span12Mux_h I__4142 (
            .O(N__21140),
            .I(N__21121));
    Span12Mux_h I__4141 (
            .O(N__21137),
            .I(N__21121));
    Span12Mux_v I__4140 (
            .O(N__21134),
            .I(N__21116));
    Span12Mux_h I__4139 (
            .O(N__21131),
            .I(N__21116));
    Odrv12 I__4138 (
            .O(N__21126),
            .I(M_this_sprites_ram_write_data_2));
    Odrv12 I__4137 (
            .O(N__21121),
            .I(M_this_sprites_ram_write_data_2));
    Odrv12 I__4136 (
            .O(N__21116),
            .I(M_this_sprites_ram_write_data_2));
    InMux I__4135 (
            .O(N__21109),
            .I(N__21106));
    LocalMux I__4134 (
            .O(N__21106),
            .I(N__21101));
    InMux I__4133 (
            .O(N__21105),
            .I(N__21096));
    InMux I__4132 (
            .O(N__21104),
            .I(N__21096));
    Odrv4 I__4131 (
            .O(N__21101),
            .I(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ));
    LocalMux I__4130 (
            .O(N__21096),
            .I(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ));
    InMux I__4129 (
            .O(N__21091),
            .I(N__21086));
    InMux I__4128 (
            .O(N__21090),
            .I(N__21082));
    InMux I__4127 (
            .O(N__21089),
            .I(N__21078));
    LocalMux I__4126 (
            .O(N__21086),
            .I(N__21074));
    InMux I__4125 (
            .O(N__21085),
            .I(N__21071));
    LocalMux I__4124 (
            .O(N__21082),
            .I(N__21067));
    InMux I__4123 (
            .O(N__21081),
            .I(N__21064));
    LocalMux I__4122 (
            .O(N__21078),
            .I(N__21061));
    InMux I__4121 (
            .O(N__21077),
            .I(N__21058));
    Span4Mux_v I__4120 (
            .O(N__21074),
            .I(N__21053));
    LocalMux I__4119 (
            .O(N__21071),
            .I(N__21053));
    InMux I__4118 (
            .O(N__21070),
            .I(N__21050));
    Span4Mux_h I__4117 (
            .O(N__21067),
            .I(N__21046));
    LocalMux I__4116 (
            .O(N__21064),
            .I(N__21043));
    Span4Mux_v I__4115 (
            .O(N__21061),
            .I(N__21038));
    LocalMux I__4114 (
            .O(N__21058),
            .I(N__21038));
    Span4Mux_v I__4113 (
            .O(N__21053),
            .I(N__21033));
    LocalMux I__4112 (
            .O(N__21050),
            .I(N__21033));
    InMux I__4111 (
            .O(N__21049),
            .I(N__21030));
    Span4Mux_v I__4110 (
            .O(N__21046),
            .I(N__21025));
    Span4Mux_h I__4109 (
            .O(N__21043),
            .I(N__21025));
    Sp12to4 I__4108 (
            .O(N__21038),
            .I(N__21022));
    Span4Mux_v I__4107 (
            .O(N__21033),
            .I(N__21019));
    LocalMux I__4106 (
            .O(N__21030),
            .I(N__21016));
    Span4Mux_h I__4105 (
            .O(N__21025),
            .I(N__21013));
    Span12Mux_v I__4104 (
            .O(N__21022),
            .I(N__21006));
    Sp12to4 I__4103 (
            .O(N__21019),
            .I(N__21006));
    Span12Mux_s8_h I__4102 (
            .O(N__21016),
            .I(N__21006));
    Odrv4 I__4101 (
            .O(N__21013),
            .I(M_this_sprites_ram_write_data_3));
    Odrv12 I__4100 (
            .O(N__21006),
            .I(M_this_sprites_ram_write_data_3));
    CascadeMux I__4099 (
            .O(N__21001),
            .I(N__20995));
    InMux I__4098 (
            .O(N__21000),
            .I(N__20992));
    InMux I__4097 (
            .O(N__20999),
            .I(N__20988));
    InMux I__4096 (
            .O(N__20998),
            .I(N__20983));
    InMux I__4095 (
            .O(N__20995),
            .I(N__20983));
    LocalMux I__4094 (
            .O(N__20992),
            .I(N__20978));
    InMux I__4093 (
            .O(N__20991),
            .I(N__20975));
    LocalMux I__4092 (
            .O(N__20988),
            .I(N__20972));
    LocalMux I__4091 (
            .O(N__20983),
            .I(N__20969));
    InMux I__4090 (
            .O(N__20982),
            .I(N__20964));
    InMux I__4089 (
            .O(N__20981),
            .I(N__20964));
    Span4Mux_v I__4088 (
            .O(N__20978),
            .I(N__20959));
    LocalMux I__4087 (
            .O(N__20975),
            .I(N__20956));
    Span4Mux_v I__4086 (
            .O(N__20972),
            .I(N__20949));
    Span4Mux_h I__4085 (
            .O(N__20969),
            .I(N__20949));
    LocalMux I__4084 (
            .O(N__20964),
            .I(N__20949));
    InMux I__4083 (
            .O(N__20963),
            .I(N__20946));
    InMux I__4082 (
            .O(N__20962),
            .I(N__20943));
    Sp12to4 I__4081 (
            .O(N__20959),
            .I(N__20938));
    Sp12to4 I__4080 (
            .O(N__20956),
            .I(N__20938));
    Span4Mux_h I__4079 (
            .O(N__20949),
            .I(N__20935));
    LocalMux I__4078 (
            .O(N__20946),
            .I(N__20932));
    LocalMux I__4077 (
            .O(N__20943),
            .I(N__20929));
    Odrv12 I__4076 (
            .O(N__20938),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__4075 (
            .O(N__20935),
            .I(M_this_vga_ramdac_en_0));
    Odrv12 I__4074 (
            .O(N__20932),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__4073 (
            .O(N__20929),
            .I(M_this_vga_ramdac_en_0));
    InMux I__4072 (
            .O(N__20920),
            .I(N__20917));
    LocalMux I__4071 (
            .O(N__20917),
            .I(N__20914));
    Span12Mux_h I__4070 (
            .O(N__20914),
            .I(N__20908));
    InMux I__4069 (
            .O(N__20913),
            .I(N__20903));
    InMux I__4068 (
            .O(N__20912),
            .I(N__20903));
    InMux I__4067 (
            .O(N__20911),
            .I(N__20900));
    Odrv12 I__4066 (
            .O(N__20908),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__4065 (
            .O(N__20903),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__4064 (
            .O(N__20900),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    CascadeMux I__4063 (
            .O(N__20893),
            .I(N__20890));
    InMux I__4062 (
            .O(N__20890),
            .I(N__20887));
    LocalMux I__4061 (
            .O(N__20887),
            .I(N__20884));
    Span12Mux_v I__4060 (
            .O(N__20884),
            .I(N__20881));
    Odrv12 I__4059 (
            .O(N__20881),
            .I(M_this_vga_signals_address_5));
    InMux I__4058 (
            .O(N__20878),
            .I(N__20875));
    LocalMux I__4057 (
            .O(N__20875),
            .I(N__20872));
    Span4Mux_h I__4056 (
            .O(N__20872),
            .I(N__20869));
    Odrv4 I__4055 (
            .O(N__20869),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    CEMux I__4054 (
            .O(N__20866),
            .I(N__20863));
    LocalMux I__4053 (
            .O(N__20863),
            .I(N__20859));
    CEMux I__4052 (
            .O(N__20862),
            .I(N__20856));
    Span4Mux_s3_v I__4051 (
            .O(N__20859),
            .I(N__20851));
    LocalMux I__4050 (
            .O(N__20856),
            .I(N__20851));
    Span4Mux_h I__4049 (
            .O(N__20851),
            .I(N__20848));
    Span4Mux_v I__4048 (
            .O(N__20848),
            .I(N__20845));
    Span4Mux_v I__4047 (
            .O(N__20845),
            .I(N__20842));
    Span4Mux_h I__4046 (
            .O(N__20842),
            .I(N__20839));
    Odrv4 I__4045 (
            .O(N__20839),
            .I(\this_sprites_ram.mem_WE_14 ));
    CEMux I__4044 (
            .O(N__20836),
            .I(N__20833));
    LocalMux I__4043 (
            .O(N__20833),
            .I(N__20829));
    CEMux I__4042 (
            .O(N__20832),
            .I(N__20826));
    Span4Mux_v I__4041 (
            .O(N__20829),
            .I(N__20821));
    LocalMux I__4040 (
            .O(N__20826),
            .I(N__20821));
    Span4Mux_h I__4039 (
            .O(N__20821),
            .I(N__20818));
    Span4Mux_v I__4038 (
            .O(N__20818),
            .I(N__20815));
    Span4Mux_h I__4037 (
            .O(N__20815),
            .I(N__20812));
    Odrv4 I__4036 (
            .O(N__20812),
            .I(\this_sprites_ram.mem_WE_12 ));
    InMux I__4035 (
            .O(N__20809),
            .I(N__20805));
    InMux I__4034 (
            .O(N__20808),
            .I(N__20802));
    LocalMux I__4033 (
            .O(N__20805),
            .I(N__20795));
    LocalMux I__4032 (
            .O(N__20802),
            .I(N__20795));
    InMux I__4031 (
            .O(N__20801),
            .I(N__20792));
    InMux I__4030 (
            .O(N__20800),
            .I(N__20789));
    Span4Mux_v I__4029 (
            .O(N__20795),
            .I(N__20781));
    LocalMux I__4028 (
            .O(N__20792),
            .I(N__20781));
    LocalMux I__4027 (
            .O(N__20789),
            .I(N__20781));
    InMux I__4026 (
            .O(N__20788),
            .I(N__20778));
    Span4Mux_v I__4025 (
            .O(N__20781),
            .I(N__20775));
    LocalMux I__4024 (
            .O(N__20778),
            .I(N__20772));
    Span4Mux_h I__4023 (
            .O(N__20775),
            .I(N__20764));
    Span4Mux_v I__4022 (
            .O(N__20772),
            .I(N__20764));
    InMux I__4021 (
            .O(N__20771),
            .I(N__20757));
    InMux I__4020 (
            .O(N__20770),
            .I(N__20757));
    InMux I__4019 (
            .O(N__20769),
            .I(N__20757));
    Odrv4 I__4018 (
            .O(N__20764),
            .I(M_this_sprites_ram_write_en_0));
    LocalMux I__4017 (
            .O(N__20757),
            .I(M_this_sprites_ram_write_en_0));
    CEMux I__4016 (
            .O(N__20752),
            .I(N__20748));
    CEMux I__4015 (
            .O(N__20751),
            .I(N__20745));
    LocalMux I__4014 (
            .O(N__20748),
            .I(N__20742));
    LocalMux I__4013 (
            .O(N__20745),
            .I(N__20739));
    Span4Mux_h I__4012 (
            .O(N__20742),
            .I(N__20736));
    Span4Mux_h I__4011 (
            .O(N__20739),
            .I(N__20733));
    Span4Mux_v I__4010 (
            .O(N__20736),
            .I(N__20730));
    Span4Mux_h I__4009 (
            .O(N__20733),
            .I(N__20727));
    Span4Mux_h I__4008 (
            .O(N__20730),
            .I(N__20724));
    Span4Mux_v I__4007 (
            .O(N__20727),
            .I(N__20721));
    Odrv4 I__4006 (
            .O(N__20724),
            .I(\this_sprites_ram.mem_WE_10 ));
    Odrv4 I__4005 (
            .O(N__20721),
            .I(\this_sprites_ram.mem_WE_10 ));
    InMux I__4004 (
            .O(N__20716),
            .I(N__20713));
    LocalMux I__4003 (
            .O(N__20713),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__4002 (
            .O(N__20710),
            .I(N__20707));
    LocalMux I__4001 (
            .O(N__20707),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    InMux I__4000 (
            .O(N__20704),
            .I(N__20701));
    LocalMux I__3999 (
            .O(N__20701),
            .I(N__20698));
    Span4Mux_h I__3998 (
            .O(N__20698),
            .I(N__20695));
    Span4Mux_v I__3997 (
            .O(N__20695),
            .I(N__20692));
    Span4Mux_h I__3996 (
            .O(N__20692),
            .I(N__20689));
    Odrv4 I__3995 (
            .O(N__20689),
            .I(\this_sprites_ram.mem_out_bus6_1 ));
    InMux I__3994 (
            .O(N__20686),
            .I(N__20683));
    LocalMux I__3993 (
            .O(N__20683),
            .I(N__20680));
    Span4Mux_h I__3992 (
            .O(N__20680),
            .I(N__20677));
    Span4Mux_v I__3991 (
            .O(N__20677),
            .I(N__20674));
    Span4Mux_v I__3990 (
            .O(N__20674),
            .I(N__20671));
    Odrv4 I__3989 (
            .O(N__20671),
            .I(\this_sprites_ram.mem_out_bus2_1 ));
    InMux I__3988 (
            .O(N__20668),
            .I(N__20665));
    LocalMux I__3987 (
            .O(N__20665),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ));
    InMux I__3986 (
            .O(N__20662),
            .I(N__20659));
    LocalMux I__3985 (
            .O(N__20659),
            .I(N__20656));
    Odrv12 I__3984 (
            .O(N__20656),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ));
    InMux I__3983 (
            .O(N__20653),
            .I(N__20650));
    LocalMux I__3982 (
            .O(N__20650),
            .I(N__20647));
    Span4Mux_h I__3981 (
            .O(N__20647),
            .I(N__20644));
    Odrv4 I__3980 (
            .O(N__20644),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ));
    InMux I__3979 (
            .O(N__20641),
            .I(N__20638));
    LocalMux I__3978 (
            .O(N__20638),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2 ));
    InMux I__3977 (
            .O(N__20635),
            .I(N__20632));
    LocalMux I__3976 (
            .O(N__20632),
            .I(N__20629));
    Span4Mux_v I__3975 (
            .O(N__20629),
            .I(N__20626));
    Span4Mux_h I__3974 (
            .O(N__20626),
            .I(N__20623));
    Span4Mux_h I__3973 (
            .O(N__20623),
            .I(N__20620));
    Odrv4 I__3972 (
            .O(N__20620),
            .I(M_this_ppu_vram_data_2));
    InMux I__3971 (
            .O(N__20617),
            .I(N__20614));
    LocalMux I__3970 (
            .O(N__20614),
            .I(N__20609));
    InMux I__3969 (
            .O(N__20613),
            .I(N__20605));
    InMux I__3968 (
            .O(N__20612),
            .I(N__20602));
    Span4Mux_h I__3967 (
            .O(N__20609),
            .I(N__20598));
    InMux I__3966 (
            .O(N__20608),
            .I(N__20595));
    LocalMux I__3965 (
            .O(N__20605),
            .I(N__20590));
    LocalMux I__3964 (
            .O(N__20602),
            .I(N__20590));
    InMux I__3963 (
            .O(N__20601),
            .I(N__20587));
    Odrv4 I__3962 (
            .O(N__20598),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__3961 (
            .O(N__20595),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv12 I__3960 (
            .O(N__20590),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__3959 (
            .O(N__20587),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    InMux I__3958 (
            .O(N__20578),
            .I(N__20573));
    InMux I__3957 (
            .O(N__20577),
            .I(N__20568));
    InMux I__3956 (
            .O(N__20576),
            .I(N__20568));
    LocalMux I__3955 (
            .O(N__20573),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    LocalMux I__3954 (
            .O(N__20568),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    CEMux I__3953 (
            .O(N__20563),
            .I(N__20560));
    LocalMux I__3952 (
            .O(N__20560),
            .I(N__20557));
    Span4Mux_s2_v I__3951 (
            .O(N__20557),
            .I(N__20553));
    CEMux I__3950 (
            .O(N__20556),
            .I(N__20550));
    Sp12to4 I__3949 (
            .O(N__20553),
            .I(N__20545));
    LocalMux I__3948 (
            .O(N__20550),
            .I(N__20545));
    Span12Mux_v I__3947 (
            .O(N__20545),
            .I(N__20542));
    Odrv12 I__3946 (
            .O(N__20542),
            .I(\this_sprites_ram.mem_WE_0 ));
    CascadeMux I__3945 (
            .O(N__20539),
            .I(N__20536));
    CascadeBuf I__3944 (
            .O(N__20536),
            .I(N__20533));
    CascadeMux I__3943 (
            .O(N__20533),
            .I(N__20530));
    InMux I__3942 (
            .O(N__20530),
            .I(N__20526));
    InMux I__3941 (
            .O(N__20529),
            .I(N__20522));
    LocalMux I__3940 (
            .O(N__20526),
            .I(N__20519));
    InMux I__3939 (
            .O(N__20525),
            .I(N__20516));
    LocalMux I__3938 (
            .O(N__20522),
            .I(N__20511));
    Span12Mux_s9_v I__3937 (
            .O(N__20519),
            .I(N__20511));
    LocalMux I__3936 (
            .O(N__20516),
            .I(M_this_ppu_map_addr_6));
    Odrv12 I__3935 (
            .O(N__20511),
            .I(M_this_ppu_map_addr_6));
    CascadeMux I__3934 (
            .O(N__20506),
            .I(N__20503));
    CascadeBuf I__3933 (
            .O(N__20503),
            .I(N__20500));
    CascadeMux I__3932 (
            .O(N__20500),
            .I(N__20497));
    InMux I__3931 (
            .O(N__20497),
            .I(N__20494));
    LocalMux I__3930 (
            .O(N__20494),
            .I(N__20490));
    InMux I__3929 (
            .O(N__20493),
            .I(N__20487));
    Span4Mux_h I__3928 (
            .O(N__20490),
            .I(N__20484));
    LocalMux I__3927 (
            .O(N__20487),
            .I(N__20479));
    Sp12to4 I__3926 (
            .O(N__20484),
            .I(N__20476));
    InMux I__3925 (
            .O(N__20483),
            .I(N__20473));
    InMux I__3924 (
            .O(N__20482),
            .I(N__20470));
    Span4Mux_h I__3923 (
            .O(N__20479),
            .I(N__20467));
    Span12Mux_s10_v I__3922 (
            .O(N__20476),
            .I(N__20464));
    LocalMux I__3921 (
            .O(N__20473),
            .I(M_this_ppu_map_addr_5));
    LocalMux I__3920 (
            .O(N__20470),
            .I(M_this_ppu_map_addr_5));
    Odrv4 I__3919 (
            .O(N__20467),
            .I(M_this_ppu_map_addr_5));
    Odrv12 I__3918 (
            .O(N__20464),
            .I(M_this_ppu_map_addr_5));
    CascadeMux I__3917 (
            .O(N__20455),
            .I(N__20452));
    CascadeBuf I__3916 (
            .O(N__20452),
            .I(N__20449));
    CascadeMux I__3915 (
            .O(N__20449),
            .I(N__20446));
    CascadeBuf I__3914 (
            .O(N__20446),
            .I(N__20443));
    CascadeMux I__3913 (
            .O(N__20443),
            .I(N__20440));
    CascadeBuf I__3912 (
            .O(N__20440),
            .I(N__20437));
    CascadeMux I__3911 (
            .O(N__20437),
            .I(N__20434));
    CascadeBuf I__3910 (
            .O(N__20434),
            .I(N__20431));
    CascadeMux I__3909 (
            .O(N__20431),
            .I(N__20428));
    CascadeBuf I__3908 (
            .O(N__20428),
            .I(N__20425));
    CascadeMux I__3907 (
            .O(N__20425),
            .I(N__20422));
    CascadeBuf I__3906 (
            .O(N__20422),
            .I(N__20419));
    CascadeMux I__3905 (
            .O(N__20419),
            .I(N__20416));
    CascadeBuf I__3904 (
            .O(N__20416),
            .I(N__20413));
    CascadeMux I__3903 (
            .O(N__20413),
            .I(N__20410));
    CascadeBuf I__3902 (
            .O(N__20410),
            .I(N__20407));
    CascadeMux I__3901 (
            .O(N__20407),
            .I(N__20404));
    CascadeBuf I__3900 (
            .O(N__20404),
            .I(N__20401));
    CascadeMux I__3899 (
            .O(N__20401),
            .I(N__20398));
    CascadeBuf I__3898 (
            .O(N__20398),
            .I(N__20395));
    CascadeMux I__3897 (
            .O(N__20395),
            .I(N__20392));
    CascadeBuf I__3896 (
            .O(N__20392),
            .I(N__20389));
    CascadeMux I__3895 (
            .O(N__20389),
            .I(N__20386));
    CascadeBuf I__3894 (
            .O(N__20386),
            .I(N__20383));
    CascadeMux I__3893 (
            .O(N__20383),
            .I(N__20380));
    CascadeBuf I__3892 (
            .O(N__20380),
            .I(N__20377));
    CascadeMux I__3891 (
            .O(N__20377),
            .I(N__20374));
    CascadeBuf I__3890 (
            .O(N__20374),
            .I(N__20371));
    CascadeMux I__3889 (
            .O(N__20371),
            .I(N__20368));
    CascadeBuf I__3888 (
            .O(N__20368),
            .I(N__20365));
    CascadeMux I__3887 (
            .O(N__20365),
            .I(N__20361));
    CascadeMux I__3886 (
            .O(N__20364),
            .I(N__20358));
    InMux I__3885 (
            .O(N__20361),
            .I(N__20353));
    InMux I__3884 (
            .O(N__20358),
            .I(N__20349));
    InMux I__3883 (
            .O(N__20357),
            .I(N__20346));
    CascadeMux I__3882 (
            .O(N__20356),
            .I(N__20343));
    LocalMux I__3881 (
            .O(N__20353),
            .I(N__20340));
    CascadeMux I__3880 (
            .O(N__20352),
            .I(N__20337));
    LocalMux I__3879 (
            .O(N__20349),
            .I(N__20334));
    LocalMux I__3878 (
            .O(N__20346),
            .I(N__20331));
    InMux I__3877 (
            .O(N__20343),
            .I(N__20328));
    Span4Mux_v I__3876 (
            .O(N__20340),
            .I(N__20325));
    InMux I__3875 (
            .O(N__20337),
            .I(N__20322));
    Span4Mux_h I__3874 (
            .O(N__20334),
            .I(N__20315));
    Span4Mux_v I__3873 (
            .O(N__20331),
            .I(N__20315));
    LocalMux I__3872 (
            .O(N__20328),
            .I(N__20315));
    Span4Mux_v I__3871 (
            .O(N__20325),
            .I(N__20312));
    LocalMux I__3870 (
            .O(N__20322),
            .I(M_this_ppu_sprites_addr_5));
    Odrv4 I__3869 (
            .O(N__20315),
            .I(M_this_ppu_sprites_addr_5));
    Odrv4 I__3868 (
            .O(N__20312),
            .I(M_this_ppu_sprites_addr_5));
    InMux I__3867 (
            .O(N__20305),
            .I(N__20300));
    InMux I__3866 (
            .O(N__20304),
            .I(N__20297));
    InMux I__3865 (
            .O(N__20303),
            .I(N__20294));
    LocalMux I__3864 (
            .O(N__20300),
            .I(N__20289));
    LocalMux I__3863 (
            .O(N__20297),
            .I(N__20289));
    LocalMux I__3862 (
            .O(N__20294),
            .I(N__20286));
    Span4Mux_v I__3861 (
            .O(N__20289),
            .I(N__20283));
    Span4Mux_v I__3860 (
            .O(N__20286),
            .I(N__20280));
    Odrv4 I__3859 (
            .O(N__20283),
            .I(\this_ppu.un1_M_vaddress_q_c2 ));
    Odrv4 I__3858 (
            .O(N__20280),
            .I(\this_ppu.un1_M_vaddress_q_c2 ));
    CascadeMux I__3857 (
            .O(N__20275),
            .I(\this_ppu.M_state_q_i_1_cascade_ ));
    InMux I__3856 (
            .O(N__20272),
            .I(N__20269));
    LocalMux I__3855 (
            .O(N__20269),
            .I(\this_ppu.M_last_q_RNIMRAD5_2 ));
    InMux I__3854 (
            .O(N__20266),
            .I(N__20263));
    LocalMux I__3853 (
            .O(N__20263),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_3 ));
    CascadeMux I__3852 (
            .O(N__20260),
            .I(N__20256));
    CascadeMux I__3851 (
            .O(N__20259),
            .I(N__20253));
    InMux I__3850 (
            .O(N__20256),
            .I(N__20250));
    InMux I__3849 (
            .O(N__20253),
            .I(N__20247));
    LocalMux I__3848 (
            .O(N__20250),
            .I(\this_ppu.M_count_qZ1Z_3 ));
    LocalMux I__3847 (
            .O(N__20247),
            .I(\this_ppu.M_count_qZ1Z_3 ));
    CascadeMux I__3846 (
            .O(N__20242),
            .I(N__20239));
    InMux I__3845 (
            .O(N__20239),
            .I(N__20235));
    InMux I__3844 (
            .O(N__20238),
            .I(N__20232));
    LocalMux I__3843 (
            .O(N__20235),
            .I(\this_ppu.M_count_qZ1Z_4 ));
    LocalMux I__3842 (
            .O(N__20232),
            .I(\this_ppu.M_count_qZ1Z_4 ));
    CascadeMux I__3841 (
            .O(N__20227),
            .I(N__20224));
    InMux I__3840 (
            .O(N__20224),
            .I(N__20221));
    LocalMux I__3839 (
            .O(N__20221),
            .I(N__20217));
    InMux I__3838 (
            .O(N__20220),
            .I(N__20214));
    Odrv4 I__3837 (
            .O(N__20217),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    LocalMux I__3836 (
            .O(N__20214),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    InMux I__3835 (
            .O(N__20209),
            .I(N__20206));
    LocalMux I__3834 (
            .O(N__20206),
            .I(\this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4 ));
    InMux I__3833 (
            .O(N__20203),
            .I(N__20199));
    InMux I__3832 (
            .O(N__20202),
            .I(N__20196));
    LocalMux I__3831 (
            .O(N__20199),
            .I(\this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_5 ));
    LocalMux I__3830 (
            .O(N__20196),
            .I(\this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_5 ));
    CascadeMux I__3829 (
            .O(N__20191),
            .I(\this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4_cascade_ ));
    CascadeMux I__3828 (
            .O(N__20188),
            .I(N__20185));
    InMux I__3827 (
            .O(N__20185),
            .I(N__20181));
    InMux I__3826 (
            .O(N__20184),
            .I(N__20178));
    LocalMux I__3825 (
            .O(N__20181),
            .I(N__20170));
    LocalMux I__3824 (
            .O(N__20178),
            .I(N__20170));
    CascadeMux I__3823 (
            .O(N__20177),
            .I(N__20167));
    CascadeMux I__3822 (
            .O(N__20176),
            .I(N__20164));
    CascadeMux I__3821 (
            .O(N__20175),
            .I(N__20161));
    Span4Mux_v I__3820 (
            .O(N__20170),
            .I(N__20156));
    InMux I__3819 (
            .O(N__20167),
            .I(N__20153));
    InMux I__3818 (
            .O(N__20164),
            .I(N__20150));
    InMux I__3817 (
            .O(N__20161),
            .I(N__20145));
    InMux I__3816 (
            .O(N__20160),
            .I(N__20145));
    InMux I__3815 (
            .O(N__20159),
            .I(N__20142));
    Odrv4 I__3814 (
            .O(N__20156),
            .I(\this_ppu.M_state_d_0_sqmuxa_1 ));
    LocalMux I__3813 (
            .O(N__20153),
            .I(\this_ppu.M_state_d_0_sqmuxa_1 ));
    LocalMux I__3812 (
            .O(N__20150),
            .I(\this_ppu.M_state_d_0_sqmuxa_1 ));
    LocalMux I__3811 (
            .O(N__20145),
            .I(\this_ppu.M_state_d_0_sqmuxa_1 ));
    LocalMux I__3810 (
            .O(N__20142),
            .I(\this_ppu.M_state_d_0_sqmuxa_1 ));
    CascadeMux I__3809 (
            .O(N__20131),
            .I(\this_ppu.M_state_d_0_sqmuxa_1_cascade_ ));
    InMux I__3808 (
            .O(N__20128),
            .I(N__20125));
    LocalMux I__3807 (
            .O(N__20125),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_5 ));
    CascadeMux I__3806 (
            .O(N__20122),
            .I(N__20119));
    InMux I__3805 (
            .O(N__20119),
            .I(N__20115));
    InMux I__3804 (
            .O(N__20118),
            .I(N__20112));
    LocalMux I__3803 (
            .O(N__20115),
            .I(\this_ppu.M_count_qZ1Z_5 ));
    LocalMux I__3802 (
            .O(N__20112),
            .I(\this_ppu.M_count_qZ1Z_5 ));
    InMux I__3801 (
            .O(N__20107),
            .I(N__20101));
    InMux I__3800 (
            .O(N__20106),
            .I(N__20101));
    LocalMux I__3799 (
            .O(N__20101),
            .I(N__20088));
    InMux I__3798 (
            .O(N__20100),
            .I(N__20081));
    InMux I__3797 (
            .O(N__20099),
            .I(N__20081));
    InMux I__3796 (
            .O(N__20098),
            .I(N__20081));
    InMux I__3795 (
            .O(N__20097),
            .I(N__20078));
    InMux I__3794 (
            .O(N__20096),
            .I(N__20075));
    InMux I__3793 (
            .O(N__20095),
            .I(N__20072));
    InMux I__3792 (
            .O(N__20094),
            .I(N__20069));
    InMux I__3791 (
            .O(N__20093),
            .I(N__20062));
    InMux I__3790 (
            .O(N__20092),
            .I(N__20062));
    InMux I__3789 (
            .O(N__20091),
            .I(N__20062));
    Span4Mux_h I__3788 (
            .O(N__20088),
            .I(N__20059));
    LocalMux I__3787 (
            .O(N__20081),
            .I(N__20056));
    LocalMux I__3786 (
            .O(N__20078),
            .I(\this_ppu.M_state_q_i_1 ));
    LocalMux I__3785 (
            .O(N__20075),
            .I(\this_ppu.M_state_q_i_1 ));
    LocalMux I__3784 (
            .O(N__20072),
            .I(\this_ppu.M_state_q_i_1 ));
    LocalMux I__3783 (
            .O(N__20069),
            .I(\this_ppu.M_state_q_i_1 ));
    LocalMux I__3782 (
            .O(N__20062),
            .I(\this_ppu.M_state_q_i_1 ));
    Odrv4 I__3781 (
            .O(N__20059),
            .I(\this_ppu.M_state_q_i_1 ));
    Odrv4 I__3780 (
            .O(N__20056),
            .I(\this_ppu.M_state_q_i_1 ));
    CascadeMux I__3779 (
            .O(N__20041),
            .I(N__20037));
    InMux I__3778 (
            .O(N__20040),
            .I(N__20032));
    InMux I__3777 (
            .O(N__20037),
            .I(N__20032));
    LocalMux I__3776 (
            .O(N__20032),
            .I(\this_ppu.M_count_qZ0Z_7 ));
    InMux I__3775 (
            .O(N__20029),
            .I(N__20019));
    InMux I__3774 (
            .O(N__20028),
            .I(N__20016));
    InMux I__3773 (
            .O(N__20027),
            .I(N__20013));
    InMux I__3772 (
            .O(N__20026),
            .I(N__20006));
    InMux I__3771 (
            .O(N__20025),
            .I(N__20006));
    InMux I__3770 (
            .O(N__20024),
            .I(N__20006));
    InMux I__3769 (
            .O(N__20023),
            .I(N__20001));
    InMux I__3768 (
            .O(N__20022),
            .I(N__20001));
    LocalMux I__3767 (
            .O(N__20019),
            .I(\this_ppu.N_82_i ));
    LocalMux I__3766 (
            .O(N__20016),
            .I(\this_ppu.N_82_i ));
    LocalMux I__3765 (
            .O(N__20013),
            .I(\this_ppu.N_82_i ));
    LocalMux I__3764 (
            .O(N__20006),
            .I(\this_ppu.N_82_i ));
    LocalMux I__3763 (
            .O(N__20001),
            .I(\this_ppu.N_82_i ));
    InMux I__3762 (
            .O(N__19990),
            .I(N__19987));
    LocalMux I__3761 (
            .O(N__19987),
            .I(\this_ppu.un1_M_count_q_1_axb_7 ));
    InMux I__3760 (
            .O(N__19984),
            .I(N__19981));
    LocalMux I__3759 (
            .O(N__19981),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__3758 (
            .O(N__19978),
            .I(N__19975));
    LocalMux I__3757 (
            .O(N__19975),
            .I(N__19972));
    Span4Mux_h I__3756 (
            .O(N__19972),
            .I(N__19969));
    Sp12to4 I__3755 (
            .O(N__19969),
            .I(N__19966));
    Span12Mux_v I__3754 (
            .O(N__19966),
            .I(N__19963));
    Odrv12 I__3753 (
            .O(N__19963),
            .I(\this_sprites_ram.mem_out_bus6_2 ));
    InMux I__3752 (
            .O(N__19960),
            .I(N__19957));
    LocalMux I__3751 (
            .O(N__19957),
            .I(N__19954));
    Span4Mux_v I__3750 (
            .O(N__19954),
            .I(N__19951));
    Sp12to4 I__3749 (
            .O(N__19951),
            .I(N__19948));
    Odrv12 I__3748 (
            .O(N__19948),
            .I(\this_sprites_ram.mem_out_bus2_2 ));
    CascadeMux I__3747 (
            .O(N__19945),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_ ));
    InMux I__3746 (
            .O(N__19942),
            .I(N__19939));
    LocalMux I__3745 (
            .O(N__19939),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0 ));
    InMux I__3744 (
            .O(N__19936),
            .I(N__19933));
    LocalMux I__3743 (
            .O(N__19933),
            .I(N__19930));
    Odrv4 I__3742 (
            .O(N__19930),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ));
    InMux I__3741 (
            .O(N__19927),
            .I(N__19924));
    LocalMux I__3740 (
            .O(N__19924),
            .I(N__19921));
    Span4Mux_v I__3739 (
            .O(N__19921),
            .I(N__19918));
    Odrv4 I__3738 (
            .O(N__19918),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ));
    CascadeMux I__3737 (
            .O(N__19915),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ));
    InMux I__3736 (
            .O(N__19912),
            .I(N__19909));
    LocalMux I__3735 (
            .O(N__19909),
            .I(N__19906));
    Span4Mux_v I__3734 (
            .O(N__19906),
            .I(N__19903));
    Sp12to4 I__3733 (
            .O(N__19903),
            .I(N__19900));
    Odrv12 I__3732 (
            .O(N__19900),
            .I(M_this_ppu_vram_data_1));
    InMux I__3731 (
            .O(N__19897),
            .I(N__19894));
    LocalMux I__3730 (
            .O(N__19894),
            .I(N__19891));
    Span4Mux_h I__3729 (
            .O(N__19891),
            .I(N__19888));
    Span4Mux_h I__3728 (
            .O(N__19888),
            .I(N__19885));
    Odrv4 I__3727 (
            .O(N__19885),
            .I(\this_sprites_ram.mem_out_bus5_1 ));
    InMux I__3726 (
            .O(N__19882),
            .I(N__19879));
    LocalMux I__3725 (
            .O(N__19879),
            .I(N__19876));
    Span4Mux_h I__3724 (
            .O(N__19876),
            .I(N__19873));
    Span4Mux_v I__3723 (
            .O(N__19873),
            .I(N__19870));
    Span4Mux_v I__3722 (
            .O(N__19870),
            .I(N__19867));
    Span4Mux_v I__3721 (
            .O(N__19867),
            .I(N__19864));
    Odrv4 I__3720 (
            .O(N__19864),
            .I(\this_sprites_ram.mem_out_bus1_1 ));
    InMux I__3719 (
            .O(N__19861),
            .I(N__19858));
    LocalMux I__3718 (
            .O(N__19858),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ));
    CascadeMux I__3717 (
            .O(N__19855),
            .I(\this_ppu.N_91_cascade_ ));
    InMux I__3716 (
            .O(N__19852),
            .I(N__19848));
    CascadeMux I__3715 (
            .O(N__19851),
            .I(N__19845));
    LocalMux I__3714 (
            .O(N__19848),
            .I(N__19842));
    InMux I__3713 (
            .O(N__19845),
            .I(N__19839));
    Odrv4 I__3712 (
            .O(N__19842),
            .I(\this_ppu.M_count_qZ1Z_1 ));
    LocalMux I__3711 (
            .O(N__19839),
            .I(\this_ppu.M_count_qZ1Z_1 ));
    CascadeMux I__3710 (
            .O(N__19834),
            .I(N__19830));
    InMux I__3709 (
            .O(N__19833),
            .I(N__19827));
    InMux I__3708 (
            .O(N__19830),
            .I(N__19824));
    LocalMux I__3707 (
            .O(N__19827),
            .I(N__19821));
    LocalMux I__3706 (
            .O(N__19824),
            .I(N__19818));
    Odrv4 I__3705 (
            .O(N__19821),
            .I(\this_ppu.M_count_qZ1Z_2 ));
    Odrv4 I__3704 (
            .O(N__19818),
            .I(\this_ppu.M_count_qZ1Z_2 ));
    InMux I__3703 (
            .O(N__19813),
            .I(N__19809));
    CascadeMux I__3702 (
            .O(N__19812),
            .I(N__19805));
    LocalMux I__3701 (
            .O(N__19809),
            .I(N__19802));
    InMux I__3700 (
            .O(N__19808),
            .I(N__19799));
    InMux I__3699 (
            .O(N__19805),
            .I(N__19796));
    Odrv4 I__3698 (
            .O(N__19802),
            .I(\this_ppu.M_count_qZ1Z_0 ));
    LocalMux I__3697 (
            .O(N__19799),
            .I(\this_ppu.M_count_qZ1Z_0 ));
    LocalMux I__3696 (
            .O(N__19796),
            .I(\this_ppu.M_count_qZ1Z_0 ));
    InMux I__3695 (
            .O(N__19789),
            .I(N__19786));
    LocalMux I__3694 (
            .O(N__19786),
            .I(N__19783));
    Span4Mux_v I__3693 (
            .O(N__19783),
            .I(N__19780));
    Span4Mux_v I__3692 (
            .O(N__19780),
            .I(N__19777));
    Sp12to4 I__3691 (
            .O(N__19777),
            .I(N__19774));
    Span12Mux_h I__3690 (
            .O(N__19774),
            .I(N__19771));
    Odrv12 I__3689 (
            .O(N__19771),
            .I(\this_sprites_ram.mem_out_bus6_0 ));
    InMux I__3688 (
            .O(N__19768),
            .I(N__19765));
    LocalMux I__3687 (
            .O(N__19765),
            .I(N__19762));
    Span4Mux_h I__3686 (
            .O(N__19762),
            .I(N__19759));
    Span4Mux_h I__3685 (
            .O(N__19759),
            .I(N__19756));
    Odrv4 I__3684 (
            .O(N__19756),
            .I(\this_sprites_ram.mem_out_bus2_0 ));
    InMux I__3683 (
            .O(N__19753),
            .I(N__19747));
    InMux I__3682 (
            .O(N__19752),
            .I(N__19742));
    InMux I__3681 (
            .O(N__19751),
            .I(N__19742));
    InMux I__3680 (
            .O(N__19750),
            .I(N__19739));
    LocalMux I__3679 (
            .O(N__19747),
            .I(N__19736));
    LocalMux I__3678 (
            .O(N__19742),
            .I(N__19733));
    LocalMux I__3677 (
            .O(N__19739),
            .I(N__19730));
    Span4Mux_h I__3676 (
            .O(N__19736),
            .I(N__19727));
    Span4Mux_v I__3675 (
            .O(N__19733),
            .I(N__19724));
    Span4Mux_h I__3674 (
            .O(N__19730),
            .I(N__19721));
    Odrv4 I__3673 (
            .O(N__19727),
            .I(\this_vga_signals.if_m8_0_a3_1_1_1 ));
    Odrv4 I__3672 (
            .O(N__19724),
            .I(\this_vga_signals.if_m8_0_a3_1_1_1 ));
    Odrv4 I__3671 (
            .O(N__19721),
            .I(\this_vga_signals.if_m8_0_a3_1_1_1 ));
    CascadeMux I__3670 (
            .O(N__19714),
            .I(N__19711));
    InMux I__3669 (
            .O(N__19711),
            .I(N__19697));
    InMux I__3668 (
            .O(N__19710),
            .I(N__19694));
    InMux I__3667 (
            .O(N__19709),
            .I(N__19687));
    InMux I__3666 (
            .O(N__19708),
            .I(N__19687));
    InMux I__3665 (
            .O(N__19707),
            .I(N__19684));
    CascadeMux I__3664 (
            .O(N__19706),
            .I(N__19681));
    CascadeMux I__3663 (
            .O(N__19705),
            .I(N__19677));
    CascadeMux I__3662 (
            .O(N__19704),
            .I(N__19672));
    InMux I__3661 (
            .O(N__19703),
            .I(N__19668));
    InMux I__3660 (
            .O(N__19702),
            .I(N__19665));
    InMux I__3659 (
            .O(N__19701),
            .I(N__19660));
    InMux I__3658 (
            .O(N__19700),
            .I(N__19657));
    LocalMux I__3657 (
            .O(N__19697),
            .I(N__19652));
    LocalMux I__3656 (
            .O(N__19694),
            .I(N__19652));
    InMux I__3655 (
            .O(N__19693),
            .I(N__19649));
    CascadeMux I__3654 (
            .O(N__19692),
            .I(N__19645));
    LocalMux I__3653 (
            .O(N__19687),
            .I(N__19638));
    LocalMux I__3652 (
            .O(N__19684),
            .I(N__19635));
    InMux I__3651 (
            .O(N__19681),
            .I(N__19630));
    InMux I__3650 (
            .O(N__19680),
            .I(N__19630));
    InMux I__3649 (
            .O(N__19677),
            .I(N__19625));
    InMux I__3648 (
            .O(N__19676),
            .I(N__19625));
    InMux I__3647 (
            .O(N__19675),
            .I(N__19618));
    InMux I__3646 (
            .O(N__19672),
            .I(N__19618));
    InMux I__3645 (
            .O(N__19671),
            .I(N__19618));
    LocalMux I__3644 (
            .O(N__19668),
            .I(N__19612));
    LocalMux I__3643 (
            .O(N__19665),
            .I(N__19609));
    InMux I__3642 (
            .O(N__19664),
            .I(N__19604));
    InMux I__3641 (
            .O(N__19663),
            .I(N__19604));
    LocalMux I__3640 (
            .O(N__19660),
            .I(N__19601));
    LocalMux I__3639 (
            .O(N__19657),
            .I(N__19594));
    Span4Mux_v I__3638 (
            .O(N__19652),
            .I(N__19594));
    LocalMux I__3637 (
            .O(N__19649),
            .I(N__19594));
    InMux I__3636 (
            .O(N__19648),
            .I(N__19587));
    InMux I__3635 (
            .O(N__19645),
            .I(N__19587));
    InMux I__3634 (
            .O(N__19644),
            .I(N__19587));
    InMux I__3633 (
            .O(N__19643),
            .I(N__19584));
    InMux I__3632 (
            .O(N__19642),
            .I(N__19579));
    InMux I__3631 (
            .O(N__19641),
            .I(N__19579));
    Span4Mux_v I__3630 (
            .O(N__19638),
            .I(N__19574));
    Span4Mux_v I__3629 (
            .O(N__19635),
            .I(N__19574));
    LocalMux I__3628 (
            .O(N__19630),
            .I(N__19567));
    LocalMux I__3627 (
            .O(N__19625),
            .I(N__19567));
    LocalMux I__3626 (
            .O(N__19618),
            .I(N__19567));
    InMux I__3625 (
            .O(N__19617),
            .I(N__19562));
    InMux I__3624 (
            .O(N__19616),
            .I(N__19562));
    InMux I__3623 (
            .O(N__19615),
            .I(N__19559));
    Span4Mux_h I__3622 (
            .O(N__19612),
            .I(N__19546));
    Span4Mux_v I__3621 (
            .O(N__19609),
            .I(N__19546));
    LocalMux I__3620 (
            .O(N__19604),
            .I(N__19546));
    Span4Mux_h I__3619 (
            .O(N__19601),
            .I(N__19546));
    Span4Mux_h I__3618 (
            .O(N__19594),
            .I(N__19546));
    LocalMux I__3617 (
            .O(N__19587),
            .I(N__19546));
    LocalMux I__3616 (
            .O(N__19584),
            .I(N__19541));
    LocalMux I__3615 (
            .O(N__19579),
            .I(N__19541));
    Odrv4 I__3614 (
            .O(N__19574),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv12 I__3613 (
            .O(N__19567),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__3612 (
            .O(N__19562),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__3611 (
            .O(N__19559),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__3610 (
            .O(N__19546),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv12 I__3609 (
            .O(N__19541),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__3608 (
            .O(N__19528),
            .I(N__19514));
    CascadeMux I__3607 (
            .O(N__19527),
            .I(N__19509));
    CascadeMux I__3606 (
            .O(N__19526),
            .I(N__19504));
    InMux I__3605 (
            .O(N__19525),
            .I(N__19501));
    InMux I__3604 (
            .O(N__19524),
            .I(N__19492));
    InMux I__3603 (
            .O(N__19523),
            .I(N__19492));
    InMux I__3602 (
            .O(N__19522),
            .I(N__19492));
    InMux I__3601 (
            .O(N__19521),
            .I(N__19492));
    InMux I__3600 (
            .O(N__19520),
            .I(N__19489));
    InMux I__3599 (
            .O(N__19519),
            .I(N__19482));
    InMux I__3598 (
            .O(N__19518),
            .I(N__19482));
    InMux I__3597 (
            .O(N__19517),
            .I(N__19482));
    LocalMux I__3596 (
            .O(N__19514),
            .I(N__19479));
    InMux I__3595 (
            .O(N__19513),
            .I(N__19476));
    CascadeMux I__3594 (
            .O(N__19512),
            .I(N__19467));
    InMux I__3593 (
            .O(N__19509),
            .I(N__19464));
    CascadeMux I__3592 (
            .O(N__19508),
            .I(N__19459));
    InMux I__3591 (
            .O(N__19507),
            .I(N__19452));
    InMux I__3590 (
            .O(N__19504),
            .I(N__19449));
    LocalMux I__3589 (
            .O(N__19501),
            .I(N__19444));
    LocalMux I__3588 (
            .O(N__19492),
            .I(N__19444));
    LocalMux I__3587 (
            .O(N__19489),
            .I(N__19439));
    LocalMux I__3586 (
            .O(N__19482),
            .I(N__19439));
    Span4Mux_v I__3585 (
            .O(N__19479),
            .I(N__19434));
    LocalMux I__3584 (
            .O(N__19476),
            .I(N__19434));
    InMux I__3583 (
            .O(N__19475),
            .I(N__19431));
    InMux I__3582 (
            .O(N__19474),
            .I(N__19428));
    InMux I__3581 (
            .O(N__19473),
            .I(N__19423));
    InMux I__3580 (
            .O(N__19472),
            .I(N__19423));
    InMux I__3579 (
            .O(N__19471),
            .I(N__19416));
    InMux I__3578 (
            .O(N__19470),
            .I(N__19416));
    InMux I__3577 (
            .O(N__19467),
            .I(N__19416));
    LocalMux I__3576 (
            .O(N__19464),
            .I(N__19413));
    InMux I__3575 (
            .O(N__19463),
            .I(N__19410));
    InMux I__3574 (
            .O(N__19462),
            .I(N__19403));
    InMux I__3573 (
            .O(N__19459),
            .I(N__19403));
    InMux I__3572 (
            .O(N__19458),
            .I(N__19403));
    InMux I__3571 (
            .O(N__19457),
            .I(N__19396));
    InMux I__3570 (
            .O(N__19456),
            .I(N__19396));
    InMux I__3569 (
            .O(N__19455),
            .I(N__19396));
    LocalMux I__3568 (
            .O(N__19452),
            .I(N__19387));
    LocalMux I__3567 (
            .O(N__19449),
            .I(N__19387));
    Span4Mux_v I__3566 (
            .O(N__19444),
            .I(N__19387));
    Span4Mux_v I__3565 (
            .O(N__19439),
            .I(N__19387));
    Span4Mux_h I__3564 (
            .O(N__19434),
            .I(N__19380));
    LocalMux I__3563 (
            .O(N__19431),
            .I(N__19380));
    LocalMux I__3562 (
            .O(N__19428),
            .I(N__19380));
    LocalMux I__3561 (
            .O(N__19423),
            .I(N__19375));
    LocalMux I__3560 (
            .O(N__19416),
            .I(N__19375));
    Odrv12 I__3559 (
            .O(N__19413),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    LocalMux I__3558 (
            .O(N__19410),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    LocalMux I__3557 (
            .O(N__19403),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    LocalMux I__3556 (
            .O(N__19396),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    Odrv4 I__3555 (
            .O(N__19387),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    Odrv4 I__3554 (
            .O(N__19380),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    Odrv4 I__3553 (
            .O(N__19375),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    CascadeMux I__3552 (
            .O(N__19360),
            .I(N__19357));
    InMux I__3551 (
            .O(N__19357),
            .I(N__19353));
    InMux I__3550 (
            .O(N__19356),
            .I(N__19350));
    LocalMux I__3549 (
            .O(N__19353),
            .I(N__19347));
    LocalMux I__3548 (
            .O(N__19350),
            .I(N__19344));
    Span4Mux_h I__3547 (
            .O(N__19347),
            .I(N__19341));
    Span4Mux_h I__3546 (
            .O(N__19344),
            .I(N__19338));
    Odrv4 I__3545 (
            .O(N__19341),
            .I(\this_vga_signals.if_N_5_0 ));
    Odrv4 I__3544 (
            .O(N__19338),
            .I(\this_vga_signals.if_N_5_0 ));
    InMux I__3543 (
            .O(N__19333),
            .I(N__19330));
    LocalMux I__3542 (
            .O(N__19330),
            .I(N__19327));
    Odrv4 I__3541 (
            .O(N__19327),
            .I(\this_reset_cond.M_stage_qZ0Z_4 ));
    InMux I__3540 (
            .O(N__19324),
            .I(N__19321));
    LocalMux I__3539 (
            .O(N__19321),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ));
    InMux I__3538 (
            .O(N__19318),
            .I(N__19315));
    LocalMux I__3537 (
            .O(N__19315),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ));
    InMux I__3536 (
            .O(N__19312),
            .I(N__19309));
    LocalMux I__3535 (
            .O(N__19309),
            .I(N__19306));
    Span4Mux_h I__3534 (
            .O(N__19306),
            .I(N__19303));
    Odrv4 I__3533 (
            .O(N__19303),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ));
    InMux I__3532 (
            .O(N__19300),
            .I(N__19297));
    LocalMux I__3531 (
            .O(N__19297),
            .I(\this_reset_cond.M_stage_qZ0Z_5 ));
    InMux I__3530 (
            .O(N__19294),
            .I(N__19291));
    LocalMux I__3529 (
            .O(N__19291),
            .I(N__19288));
    Span4Mux_v I__3528 (
            .O(N__19288),
            .I(N__19285));
    Span4Mux_h I__3527 (
            .O(N__19285),
            .I(N__19282));
    Odrv4 I__3526 (
            .O(N__19282),
            .I(\this_sprites_ram.mem_out_bus4_1 ));
    InMux I__3525 (
            .O(N__19279),
            .I(N__19276));
    LocalMux I__3524 (
            .O(N__19276),
            .I(N__19273));
    Span4Mux_v I__3523 (
            .O(N__19273),
            .I(N__19270));
    Sp12to4 I__3522 (
            .O(N__19270),
            .I(N__19267));
    Span12Mux_h I__3521 (
            .O(N__19267),
            .I(N__19264));
    Span12Mux_v I__3520 (
            .O(N__19264),
            .I(N__19261));
    Odrv12 I__3519 (
            .O(N__19261),
            .I(\this_sprites_ram.mem_out_bus0_1 ));
    CascadeMux I__3518 (
            .O(N__19258),
            .I(N__19250));
    CascadeMux I__3517 (
            .O(N__19257),
            .I(N__19243));
    InMux I__3516 (
            .O(N__19256),
            .I(N__19238));
    CascadeMux I__3515 (
            .O(N__19255),
            .I(N__19234));
    CascadeMux I__3514 (
            .O(N__19254),
            .I(N__19225));
    CascadeMux I__3513 (
            .O(N__19253),
            .I(N__19222));
    InMux I__3512 (
            .O(N__19250),
            .I(N__19218));
    CascadeMux I__3511 (
            .O(N__19249),
            .I(N__19213));
    CascadeMux I__3510 (
            .O(N__19248),
            .I(N__19210));
    CascadeMux I__3509 (
            .O(N__19247),
            .I(N__19207));
    InMux I__3508 (
            .O(N__19246),
            .I(N__19204));
    InMux I__3507 (
            .O(N__19243),
            .I(N__19198));
    InMux I__3506 (
            .O(N__19242),
            .I(N__19193));
    InMux I__3505 (
            .O(N__19241),
            .I(N__19193));
    LocalMux I__3504 (
            .O(N__19238),
            .I(N__19190));
    InMux I__3503 (
            .O(N__19237),
            .I(N__19185));
    InMux I__3502 (
            .O(N__19234),
            .I(N__19185));
    InMux I__3501 (
            .O(N__19233),
            .I(N__19182));
    CascadeMux I__3500 (
            .O(N__19232),
            .I(N__19179));
    CascadeMux I__3499 (
            .O(N__19231),
            .I(N__19176));
    InMux I__3498 (
            .O(N__19230),
            .I(N__19173));
    InMux I__3497 (
            .O(N__19229),
            .I(N__19170));
    InMux I__3496 (
            .O(N__19228),
            .I(N__19167));
    InMux I__3495 (
            .O(N__19225),
            .I(N__19164));
    InMux I__3494 (
            .O(N__19222),
            .I(N__19159));
    InMux I__3493 (
            .O(N__19221),
            .I(N__19159));
    LocalMux I__3492 (
            .O(N__19218),
            .I(N__19156));
    InMux I__3491 (
            .O(N__19217),
            .I(N__19153));
    InMux I__3490 (
            .O(N__19216),
            .I(N__19150));
    InMux I__3489 (
            .O(N__19213),
            .I(N__19147));
    InMux I__3488 (
            .O(N__19210),
            .I(N__19142));
    InMux I__3487 (
            .O(N__19207),
            .I(N__19142));
    LocalMux I__3486 (
            .O(N__19204),
            .I(N__19135));
    InMux I__3485 (
            .O(N__19203),
            .I(N__19132));
    InMux I__3484 (
            .O(N__19202),
            .I(N__19125));
    InMux I__3483 (
            .O(N__19201),
            .I(N__19125));
    LocalMux I__3482 (
            .O(N__19198),
            .I(N__19122));
    LocalMux I__3481 (
            .O(N__19193),
            .I(N__19115));
    Span4Mux_h I__3480 (
            .O(N__19190),
            .I(N__19115));
    LocalMux I__3479 (
            .O(N__19185),
            .I(N__19115));
    LocalMux I__3478 (
            .O(N__19182),
            .I(N__19112));
    InMux I__3477 (
            .O(N__19179),
            .I(N__19107));
    InMux I__3476 (
            .O(N__19176),
            .I(N__19107));
    LocalMux I__3475 (
            .O(N__19173),
            .I(N__19104));
    LocalMux I__3474 (
            .O(N__19170),
            .I(N__19099));
    LocalMux I__3473 (
            .O(N__19167),
            .I(N__19099));
    LocalMux I__3472 (
            .O(N__19164),
            .I(N__19094));
    LocalMux I__3471 (
            .O(N__19159),
            .I(N__19094));
    Span4Mux_v I__3470 (
            .O(N__19156),
            .I(N__19089));
    LocalMux I__3469 (
            .O(N__19153),
            .I(N__19089));
    LocalMux I__3468 (
            .O(N__19150),
            .I(N__19082));
    LocalMux I__3467 (
            .O(N__19147),
            .I(N__19082));
    LocalMux I__3466 (
            .O(N__19142),
            .I(N__19082));
    InMux I__3465 (
            .O(N__19141),
            .I(N__19073));
    InMux I__3464 (
            .O(N__19140),
            .I(N__19073));
    InMux I__3463 (
            .O(N__19139),
            .I(N__19073));
    InMux I__3462 (
            .O(N__19138),
            .I(N__19073));
    Span4Mux_v I__3461 (
            .O(N__19135),
            .I(N__19070));
    LocalMux I__3460 (
            .O(N__19132),
            .I(N__19067));
    InMux I__3459 (
            .O(N__19131),
            .I(N__19064));
    InMux I__3458 (
            .O(N__19130),
            .I(N__19061));
    LocalMux I__3457 (
            .O(N__19125),
            .I(N__19058));
    Span4Mux_v I__3456 (
            .O(N__19122),
            .I(N__19053));
    Span4Mux_v I__3455 (
            .O(N__19115),
            .I(N__19053));
    Span4Mux_h I__3454 (
            .O(N__19112),
            .I(N__19048));
    LocalMux I__3453 (
            .O(N__19107),
            .I(N__19048));
    Span4Mux_h I__3452 (
            .O(N__19104),
            .I(N__19035));
    Span4Mux_v I__3451 (
            .O(N__19099),
            .I(N__19035));
    Span4Mux_v I__3450 (
            .O(N__19094),
            .I(N__19035));
    Span4Mux_v I__3449 (
            .O(N__19089),
            .I(N__19035));
    Span4Mux_v I__3448 (
            .O(N__19082),
            .I(N__19035));
    LocalMux I__3447 (
            .O(N__19073),
            .I(N__19035));
    Odrv4 I__3446 (
            .O(N__19070),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__3445 (
            .O(N__19067),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__3444 (
            .O(N__19064),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__3443 (
            .O(N__19061),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv12 I__3442 (
            .O(N__19058),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__3441 (
            .O(N__19053),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__3440 (
            .O(N__19048),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__3439 (
            .O(N__19035),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    CascadeMux I__3438 (
            .O(N__19018),
            .I(N__19015));
    InMux I__3437 (
            .O(N__19015),
            .I(N__19001));
    CascadeMux I__3436 (
            .O(N__19014),
            .I(N__18997));
    CascadeMux I__3435 (
            .O(N__19013),
            .I(N__18992));
    InMux I__3434 (
            .O(N__19012),
            .I(N__18986));
    InMux I__3433 (
            .O(N__19011),
            .I(N__18986));
    InMux I__3432 (
            .O(N__19010),
            .I(N__18979));
    InMux I__3431 (
            .O(N__19009),
            .I(N__18979));
    InMux I__3430 (
            .O(N__19008),
            .I(N__18979));
    InMux I__3429 (
            .O(N__19007),
            .I(N__18973));
    CascadeMux I__3428 (
            .O(N__19006),
            .I(N__18969));
    CascadeMux I__3427 (
            .O(N__19005),
            .I(N__18966));
    CascadeMux I__3426 (
            .O(N__19004),
            .I(N__18961));
    LocalMux I__3425 (
            .O(N__19001),
            .I(N__18957));
    InMux I__3424 (
            .O(N__19000),
            .I(N__18952));
    InMux I__3423 (
            .O(N__18997),
            .I(N__18952));
    InMux I__3422 (
            .O(N__18996),
            .I(N__18945));
    InMux I__3421 (
            .O(N__18995),
            .I(N__18945));
    InMux I__3420 (
            .O(N__18992),
            .I(N__18945));
    InMux I__3419 (
            .O(N__18991),
            .I(N__18942));
    LocalMux I__3418 (
            .O(N__18986),
            .I(N__18937));
    LocalMux I__3417 (
            .O(N__18979),
            .I(N__18937));
    InMux I__3416 (
            .O(N__18978),
            .I(N__18930));
    InMux I__3415 (
            .O(N__18977),
            .I(N__18930));
    InMux I__3414 (
            .O(N__18976),
            .I(N__18930));
    LocalMux I__3413 (
            .O(N__18973),
            .I(N__18927));
    InMux I__3412 (
            .O(N__18972),
            .I(N__18924));
    InMux I__3411 (
            .O(N__18969),
            .I(N__18921));
    InMux I__3410 (
            .O(N__18966),
            .I(N__18914));
    InMux I__3409 (
            .O(N__18965),
            .I(N__18914));
    InMux I__3408 (
            .O(N__18964),
            .I(N__18914));
    InMux I__3407 (
            .O(N__18961),
            .I(N__18910));
    InMux I__3406 (
            .O(N__18960),
            .I(N__18907));
    Span4Mux_v I__3405 (
            .O(N__18957),
            .I(N__18904));
    LocalMux I__3404 (
            .O(N__18952),
            .I(N__18901));
    LocalMux I__3403 (
            .O(N__18945),
            .I(N__18898));
    LocalMux I__3402 (
            .O(N__18942),
            .I(N__18895));
    Span4Mux_v I__3401 (
            .O(N__18937),
            .I(N__18892));
    LocalMux I__3400 (
            .O(N__18930),
            .I(N__18883));
    Span4Mux_h I__3399 (
            .O(N__18927),
            .I(N__18883));
    LocalMux I__3398 (
            .O(N__18924),
            .I(N__18883));
    LocalMux I__3397 (
            .O(N__18921),
            .I(N__18883));
    LocalMux I__3396 (
            .O(N__18914),
            .I(N__18880));
    InMux I__3395 (
            .O(N__18913),
            .I(N__18877));
    LocalMux I__3394 (
            .O(N__18910),
            .I(N__18872));
    LocalMux I__3393 (
            .O(N__18907),
            .I(N__18872));
    Span4Mux_h I__3392 (
            .O(N__18904),
            .I(N__18865));
    Span4Mux_h I__3391 (
            .O(N__18901),
            .I(N__18865));
    Span4Mux_v I__3390 (
            .O(N__18898),
            .I(N__18865));
    Span4Mux_v I__3389 (
            .O(N__18895),
            .I(N__18858));
    Span4Mux_h I__3388 (
            .O(N__18892),
            .I(N__18858));
    Span4Mux_v I__3387 (
            .O(N__18883),
            .I(N__18858));
    Span4Mux_h I__3386 (
            .O(N__18880),
            .I(N__18855));
    LocalMux I__3385 (
            .O(N__18877),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv12 I__3384 (
            .O(N__18872),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__3383 (
            .O(N__18865),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__3382 (
            .O(N__18858),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__3381 (
            .O(N__18855),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    InMux I__3380 (
            .O(N__18844),
            .I(N__18839));
    CascadeMux I__3379 (
            .O(N__18843),
            .I(N__18836));
    CascadeMux I__3378 (
            .O(N__18842),
            .I(N__18831));
    LocalMux I__3377 (
            .O(N__18839),
            .I(N__18827));
    InMux I__3376 (
            .O(N__18836),
            .I(N__18822));
    InMux I__3375 (
            .O(N__18835),
            .I(N__18822));
    InMux I__3374 (
            .O(N__18834),
            .I(N__18817));
    InMux I__3373 (
            .O(N__18831),
            .I(N__18817));
    InMux I__3372 (
            .O(N__18830),
            .I(N__18814));
    Odrv4 I__3371 (
            .O(N__18827),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__3370 (
            .O(N__18822),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__3369 (
            .O(N__18817),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__3368 (
            .O(N__18814),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    InMux I__3367 (
            .O(N__18805),
            .I(N__18802));
    LocalMux I__3366 (
            .O(N__18802),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0 ));
    InMux I__3365 (
            .O(N__18799),
            .I(N__18796));
    LocalMux I__3364 (
            .O(N__18796),
            .I(N__18793));
    Span4Mux_h I__3363 (
            .O(N__18793),
            .I(N__18790));
    Span4Mux_v I__3362 (
            .O(N__18790),
            .I(N__18787));
    Span4Mux_h I__3361 (
            .O(N__18787),
            .I(N__18784));
    Odrv4 I__3360 (
            .O(N__18784),
            .I(\this_sprites_ram.mem_out_bus4_2 ));
    InMux I__3359 (
            .O(N__18781),
            .I(N__18778));
    LocalMux I__3358 (
            .O(N__18778),
            .I(N__18775));
    Span4Mux_h I__3357 (
            .O(N__18775),
            .I(N__18772));
    Span4Mux_h I__3356 (
            .O(N__18772),
            .I(N__18769));
    Span4Mux_v I__3355 (
            .O(N__18769),
            .I(N__18766));
    Span4Mux_v I__3354 (
            .O(N__18766),
            .I(N__18763));
    Odrv4 I__3353 (
            .O(N__18763),
            .I(\this_sprites_ram.mem_out_bus0_2 ));
    CascadeMux I__3352 (
            .O(N__18760),
            .I(\this_ppu.un1_M_count_q_1_axb_0_cascade_ ));
    InMux I__3351 (
            .O(N__18757),
            .I(N__18754));
    LocalMux I__3350 (
            .O(N__18754),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_6 ));
    InMux I__3349 (
            .O(N__18751),
            .I(N__18747));
    InMux I__3348 (
            .O(N__18750),
            .I(N__18744));
    LocalMux I__3347 (
            .O(N__18747),
            .I(N__18741));
    LocalMux I__3346 (
            .O(N__18744),
            .I(N__18738));
    Span4Mux_v I__3345 (
            .O(N__18741),
            .I(N__18735));
    Odrv12 I__3344 (
            .O(N__18738),
            .I(\this_ppu.line_clk.M_last_qZ0 ));
    Odrv4 I__3343 (
            .O(N__18735),
            .I(\this_ppu.line_clk.M_last_qZ0 ));
    InMux I__3342 (
            .O(N__18730),
            .I(N__18727));
    LocalMux I__3341 (
            .O(N__18727),
            .I(M_this_vga_signals_line_clk_0));
    CascadeMux I__3340 (
            .O(N__18724),
            .I(\this_ppu.N_82_i_cascade_ ));
    InMux I__3339 (
            .O(N__18721),
            .I(N__18718));
    LocalMux I__3338 (
            .O(N__18718),
            .I(\this_ppu.M_last_q_RNIMRAD5_3 ));
    InMux I__3337 (
            .O(N__18715),
            .I(N__18712));
    LocalMux I__3336 (
            .O(N__18712),
            .I(\this_reset_cond.M_stage_qZ0Z_3 ));
    InMux I__3335 (
            .O(N__18709),
            .I(N__18706));
    LocalMux I__3334 (
            .O(N__18706),
            .I(N__18703));
    Span4Mux_h I__3333 (
            .O(N__18703),
            .I(N__18700));
    Span4Mux_v I__3332 (
            .O(N__18700),
            .I(N__18697));
    Span4Mux_h I__3331 (
            .O(N__18697),
            .I(N__18694));
    Odrv4 I__3330 (
            .O(N__18694),
            .I(\this_sprites_ram.mem_out_bus4_0 ));
    InMux I__3329 (
            .O(N__18691),
            .I(N__18688));
    LocalMux I__3328 (
            .O(N__18688),
            .I(N__18685));
    Span4Mux_h I__3327 (
            .O(N__18685),
            .I(N__18682));
    Span4Mux_h I__3326 (
            .O(N__18682),
            .I(N__18679));
    Span4Mux_v I__3325 (
            .O(N__18679),
            .I(N__18676));
    Span4Mux_v I__3324 (
            .O(N__18676),
            .I(N__18673));
    Odrv4 I__3323 (
            .O(N__18673),
            .I(\this_sprites_ram.mem_out_bus0_0 ));
    InMux I__3322 (
            .O(N__18670),
            .I(\this_ppu.un1_M_count_q_1_cry_2 ));
    InMux I__3321 (
            .O(N__18667),
            .I(N__18664));
    LocalMux I__3320 (
            .O(N__18664),
            .I(\this_ppu.M_last_q_RNIMRAD5_4 ));
    InMux I__3319 (
            .O(N__18661),
            .I(\this_ppu.un1_M_count_q_1_cry_3 ));
    InMux I__3318 (
            .O(N__18658),
            .I(\this_ppu.un1_M_count_q_1_cry_4 ));
    InMux I__3317 (
            .O(N__18655),
            .I(N__18652));
    LocalMux I__3316 (
            .O(N__18652),
            .I(\this_ppu.M_last_q_RNIMRAD5_5 ));
    InMux I__3315 (
            .O(N__18649),
            .I(\this_ppu.un1_M_count_q_1_cry_5 ));
    InMux I__3314 (
            .O(N__18646),
            .I(\this_ppu.un1_M_count_q_1_cry_6 ));
    InMux I__3313 (
            .O(N__18643),
            .I(N__18640));
    LocalMux I__3312 (
            .O(N__18640),
            .I(\this_ppu.M_last_q_RNIMRAD5_1 ));
    InMux I__3311 (
            .O(N__18637),
            .I(N__18634));
    LocalMux I__3310 (
            .O(N__18634),
            .I(\this_ppu.M_last_q_RNIMRAD5_0 ));
    InMux I__3309 (
            .O(N__18631),
            .I(N__18628));
    LocalMux I__3308 (
            .O(N__18628),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_4 ));
    InMux I__3307 (
            .O(N__18625),
            .I(N__18622));
    LocalMux I__3306 (
            .O(N__18622),
            .I(\this_vga_signals.i13_mux_0_i ));
    InMux I__3305 (
            .O(N__18619),
            .I(N__18616));
    LocalMux I__3304 (
            .O(N__18616),
            .I(N__18613));
    Odrv4 I__3303 (
            .O(N__18613),
            .I(\this_vga_signals.if_i1_mux ));
    CascadeMux I__3302 (
            .O(N__18610),
            .I(\this_vga_signals.g1_0_0_cascade_ ));
    CascadeMux I__3301 (
            .O(N__18607),
            .I(N__18604));
    InMux I__3300 (
            .O(N__18604),
            .I(N__18601));
    LocalMux I__3299 (
            .O(N__18601),
            .I(N__18598));
    Span4Mux_h I__3298 (
            .O(N__18598),
            .I(N__18595));
    Span4Mux_h I__3297 (
            .O(N__18595),
            .I(N__18592));
    Span4Mux_h I__3296 (
            .O(N__18592),
            .I(N__18589));
    Odrv4 I__3295 (
            .O(N__18589),
            .I(M_this_vga_signals_address_7));
    InMux I__3294 (
            .O(N__18586),
            .I(N__18583));
    LocalMux I__3293 (
            .O(N__18583),
            .I(N__18580));
    Span4Mux_h I__3292 (
            .O(N__18580),
            .I(N__18576));
    InMux I__3291 (
            .O(N__18579),
            .I(N__18573));
    Span4Mux_v I__3290 (
            .O(N__18576),
            .I(N__18567));
    LocalMux I__3289 (
            .O(N__18573),
            .I(N__18567));
    InMux I__3288 (
            .O(N__18572),
            .I(N__18564));
    Span4Mux_h I__3287 (
            .O(N__18567),
            .I(N__18561));
    LocalMux I__3286 (
            .O(N__18564),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__3285 (
            .O(N__18561),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    InMux I__3284 (
            .O(N__18556),
            .I(N__18553));
    LocalMux I__3283 (
            .O(N__18553),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_N_4L5_1 ));
    InMux I__3282 (
            .O(N__18550),
            .I(N__18545));
    CascadeMux I__3281 (
            .O(N__18549),
            .I(N__18541));
    CascadeMux I__3280 (
            .O(N__18548),
            .I(N__18538));
    LocalMux I__3279 (
            .O(N__18545),
            .I(N__18535));
    InMux I__3278 (
            .O(N__18544),
            .I(N__18528));
    InMux I__3277 (
            .O(N__18541),
            .I(N__18528));
    InMux I__3276 (
            .O(N__18538),
            .I(N__18528));
    Span4Mux_h I__3275 (
            .O(N__18535),
            .I(N__18523));
    LocalMux I__3274 (
            .O(N__18528),
            .I(N__18520));
    InMux I__3273 (
            .O(N__18527),
            .I(N__18517));
    InMux I__3272 (
            .O(N__18526),
            .I(N__18514));
    Span4Mux_v I__3271 (
            .O(N__18523),
            .I(N__18506));
    Span4Mux_v I__3270 (
            .O(N__18520),
            .I(N__18506));
    LocalMux I__3269 (
            .O(N__18517),
            .I(N__18506));
    LocalMux I__3268 (
            .O(N__18514),
            .I(N__18503));
    InMux I__3267 (
            .O(N__18513),
            .I(N__18500));
    Span4Mux_h I__3266 (
            .O(N__18506),
            .I(N__18497));
    Odrv12 I__3265 (
            .O(N__18503),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__3264 (
            .O(N__18500),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__3263 (
            .O(N__18497),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    CascadeMux I__3262 (
            .O(N__18490),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_N_4L5_cascade_ ));
    InMux I__3261 (
            .O(N__18487),
            .I(N__18484));
    LocalMux I__3260 (
            .O(N__18484),
            .I(\this_vga_signals.N_5_i ));
    InMux I__3259 (
            .O(N__18481),
            .I(N__18478));
    LocalMux I__3258 (
            .O(N__18478),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_0 ));
    InMux I__3257 (
            .O(N__18475),
            .I(N__18472));
    LocalMux I__3256 (
            .O(N__18472),
            .I(N__18469));
    Span12Mux_h I__3255 (
            .O(N__18469),
            .I(N__18466));
    Odrv12 I__3254 (
            .O(N__18466),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    InMux I__3253 (
            .O(N__18463),
            .I(N__18460));
    LocalMux I__3252 (
            .O(N__18460),
            .I(\this_ppu.un1_M_count_q_1_cry_0_0_c_RNOZ0 ));
    InMux I__3251 (
            .O(N__18457),
            .I(N__18454));
    LocalMux I__3250 (
            .O(N__18454),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_1 ));
    InMux I__3249 (
            .O(N__18451),
            .I(\this_ppu.un1_M_count_q_1_cry_0 ));
    InMux I__3248 (
            .O(N__18448),
            .I(N__18445));
    LocalMux I__3247 (
            .O(N__18445),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_2 ));
    InMux I__3246 (
            .O(N__18442),
            .I(\this_ppu.un1_M_count_q_1_cry_1 ));
    InMux I__3245 (
            .O(N__18439),
            .I(N__18436));
    LocalMux I__3244 (
            .O(N__18436),
            .I(N__18433));
    Span4Mux_h I__3243 (
            .O(N__18433),
            .I(N__18430));
    Odrv4 I__3242 (
            .O(N__18430),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2_0 ));
    InMux I__3241 (
            .O(N__18427),
            .I(N__18424));
    LocalMux I__3240 (
            .O(N__18424),
            .I(\this_vga_signals.g0_1_1_0 ));
    InMux I__3239 (
            .O(N__18421),
            .I(N__18417));
    InMux I__3238 (
            .O(N__18420),
            .I(N__18414));
    LocalMux I__3237 (
            .O(N__18417),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    LocalMux I__3236 (
            .O(N__18414),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    CascadeMux I__3235 (
            .O(N__18409),
            .I(\this_vga_signals.g0_1_2_0_cascade_ ));
    InMux I__3234 (
            .O(N__18406),
            .I(N__18403));
    LocalMux I__3233 (
            .O(N__18403),
            .I(\this_vga_signals.g1_3 ));
    CascadeMux I__3232 (
            .O(N__18400),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_2_cascade_ ));
    InMux I__3231 (
            .O(N__18397),
            .I(N__18386));
    InMux I__3230 (
            .O(N__18396),
            .I(N__18381));
    InMux I__3229 (
            .O(N__18395),
            .I(N__18381));
    InMux I__3228 (
            .O(N__18394),
            .I(N__18378));
    InMux I__3227 (
            .O(N__18393),
            .I(N__18373));
    InMux I__3226 (
            .O(N__18392),
            .I(N__18373));
    InMux I__3225 (
            .O(N__18391),
            .I(N__18363));
    InMux I__3224 (
            .O(N__18390),
            .I(N__18363));
    CascadeMux I__3223 (
            .O(N__18389),
            .I(N__18357));
    LocalMux I__3222 (
            .O(N__18386),
            .I(N__18349));
    LocalMux I__3221 (
            .O(N__18381),
            .I(N__18349));
    LocalMux I__3220 (
            .O(N__18378),
            .I(N__18346));
    LocalMux I__3219 (
            .O(N__18373),
            .I(N__18343));
    InMux I__3218 (
            .O(N__18372),
            .I(N__18340));
    InMux I__3217 (
            .O(N__18371),
            .I(N__18331));
    InMux I__3216 (
            .O(N__18370),
            .I(N__18331));
    InMux I__3215 (
            .O(N__18369),
            .I(N__18331));
    InMux I__3214 (
            .O(N__18368),
            .I(N__18331));
    LocalMux I__3213 (
            .O(N__18363),
            .I(N__18324));
    InMux I__3212 (
            .O(N__18362),
            .I(N__18321));
    InMux I__3211 (
            .O(N__18361),
            .I(N__18316));
    InMux I__3210 (
            .O(N__18360),
            .I(N__18316));
    InMux I__3209 (
            .O(N__18357),
            .I(N__18311));
    InMux I__3208 (
            .O(N__18356),
            .I(N__18311));
    InMux I__3207 (
            .O(N__18355),
            .I(N__18306));
    InMux I__3206 (
            .O(N__18354),
            .I(N__18306));
    Span4Mux_v I__3205 (
            .O(N__18349),
            .I(N__18295));
    Span4Mux_h I__3204 (
            .O(N__18346),
            .I(N__18295));
    Span4Mux_v I__3203 (
            .O(N__18343),
            .I(N__18295));
    LocalMux I__3202 (
            .O(N__18340),
            .I(N__18295));
    LocalMux I__3201 (
            .O(N__18331),
            .I(N__18295));
    InMux I__3200 (
            .O(N__18330),
            .I(N__18288));
    InMux I__3199 (
            .O(N__18329),
            .I(N__18288));
    InMux I__3198 (
            .O(N__18328),
            .I(N__18288));
    InMux I__3197 (
            .O(N__18327),
            .I(N__18285));
    Odrv4 I__3196 (
            .O(N__18324),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__3195 (
            .O(N__18321),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__3194 (
            .O(N__18316),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__3193 (
            .O(N__18311),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__3192 (
            .O(N__18306),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    Odrv4 I__3191 (
            .O(N__18295),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__3190 (
            .O(N__18288),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__3189 (
            .O(N__18285),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    InMux I__3188 (
            .O(N__18268),
            .I(N__18259));
    InMux I__3187 (
            .O(N__18267),
            .I(N__18256));
    InMux I__3186 (
            .O(N__18266),
            .I(N__18251));
    InMux I__3185 (
            .O(N__18265),
            .I(N__18251));
    InMux I__3184 (
            .O(N__18264),
            .I(N__18248));
    InMux I__3183 (
            .O(N__18263),
            .I(N__18243));
    InMux I__3182 (
            .O(N__18262),
            .I(N__18243));
    LocalMux I__3181 (
            .O(N__18259),
            .I(if_generate_plus_mult1_un68_sum_axb1_520));
    LocalMux I__3180 (
            .O(N__18256),
            .I(if_generate_plus_mult1_un68_sum_axb1_520));
    LocalMux I__3179 (
            .O(N__18251),
            .I(if_generate_plus_mult1_un68_sum_axb1_520));
    LocalMux I__3178 (
            .O(N__18248),
            .I(if_generate_plus_mult1_un68_sum_axb1_520));
    LocalMux I__3177 (
            .O(N__18243),
            .I(if_generate_plus_mult1_un68_sum_axb1_520));
    InMux I__3176 (
            .O(N__18232),
            .I(N__18225));
    InMux I__3175 (
            .O(N__18231),
            .I(N__18222));
    InMux I__3174 (
            .O(N__18230),
            .I(N__18214));
    InMux I__3173 (
            .O(N__18229),
            .I(N__18209));
    InMux I__3172 (
            .O(N__18228),
            .I(N__18209));
    LocalMux I__3171 (
            .O(N__18225),
            .I(N__18204));
    LocalMux I__3170 (
            .O(N__18222),
            .I(N__18204));
    InMux I__3169 (
            .O(N__18221),
            .I(N__18197));
    InMux I__3168 (
            .O(N__18220),
            .I(N__18197));
    InMux I__3167 (
            .O(N__18219),
            .I(N__18197));
    InMux I__3166 (
            .O(N__18218),
            .I(N__18194));
    InMux I__3165 (
            .O(N__18217),
            .I(N__18191));
    LocalMux I__3164 (
            .O(N__18214),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__3163 (
            .O(N__18209),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    Odrv4 I__3162 (
            .O(N__18204),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__3161 (
            .O(N__18197),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__3160 (
            .O(N__18194),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__3159 (
            .O(N__18191),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    CascadeMux I__3158 (
            .O(N__18178),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ));
    InMux I__3157 (
            .O(N__18175),
            .I(N__18172));
    LocalMux I__3156 (
            .O(N__18172),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ));
    InMux I__3155 (
            .O(N__18169),
            .I(N__18166));
    LocalMux I__3154 (
            .O(N__18166),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_i ));
    InMux I__3153 (
            .O(N__18163),
            .I(N__18160));
    LocalMux I__3152 (
            .O(N__18160),
            .I(N__18157));
    Span4Mux_h I__3151 (
            .O(N__18157),
            .I(N__18153));
    InMux I__3150 (
            .O(N__18156),
            .I(N__18150));
    Odrv4 I__3149 (
            .O(N__18153),
            .I(\this_vga_signals.g2_0_0_0 ));
    LocalMux I__3148 (
            .O(N__18150),
            .I(\this_vga_signals.g2_0_0_0 ));
    InMux I__3147 (
            .O(N__18145),
            .I(N__18142));
    LocalMux I__3146 (
            .O(N__18142),
            .I(N__18138));
    InMux I__3145 (
            .O(N__18141),
            .I(N__18135));
    Odrv12 I__3144 (
            .O(N__18138),
            .I(\this_vga_signals.g1_1 ));
    LocalMux I__3143 (
            .O(N__18135),
            .I(\this_vga_signals.g1_1 ));
    CascadeMux I__3142 (
            .O(N__18130),
            .I(N__18124));
    CascadeMux I__3141 (
            .O(N__18129),
            .I(N__18120));
    CascadeMux I__3140 (
            .O(N__18128),
            .I(N__18117));
    CascadeMux I__3139 (
            .O(N__18127),
            .I(N__18112));
    InMux I__3138 (
            .O(N__18124),
            .I(N__18109));
    CascadeMux I__3137 (
            .O(N__18123),
            .I(N__18106));
    InMux I__3136 (
            .O(N__18120),
            .I(N__18097));
    InMux I__3135 (
            .O(N__18117),
            .I(N__18094));
    InMux I__3134 (
            .O(N__18116),
            .I(N__18091));
    CascadeMux I__3133 (
            .O(N__18115),
            .I(N__18085));
    InMux I__3132 (
            .O(N__18112),
            .I(N__18080));
    LocalMux I__3131 (
            .O(N__18109),
            .I(N__18077));
    InMux I__3130 (
            .O(N__18106),
            .I(N__18074));
    InMux I__3129 (
            .O(N__18105),
            .I(N__18071));
    InMux I__3128 (
            .O(N__18104),
            .I(N__18068));
    InMux I__3127 (
            .O(N__18103),
            .I(N__18065));
    InMux I__3126 (
            .O(N__18102),
            .I(N__18060));
    InMux I__3125 (
            .O(N__18101),
            .I(N__18060));
    CascadeMux I__3124 (
            .O(N__18100),
            .I(N__18057));
    LocalMux I__3123 (
            .O(N__18097),
            .I(N__18054));
    LocalMux I__3122 (
            .O(N__18094),
            .I(N__18051));
    LocalMux I__3121 (
            .O(N__18091),
            .I(N__18048));
    InMux I__3120 (
            .O(N__18090),
            .I(N__18043));
    InMux I__3119 (
            .O(N__18089),
            .I(N__18043));
    CascadeMux I__3118 (
            .O(N__18088),
            .I(N__18039));
    InMux I__3117 (
            .O(N__18085),
            .I(N__18035));
    InMux I__3116 (
            .O(N__18084),
            .I(N__18032));
    CascadeMux I__3115 (
            .O(N__18083),
            .I(N__18028));
    LocalMux I__3114 (
            .O(N__18080),
            .I(N__18019));
    Span4Mux_v I__3113 (
            .O(N__18077),
            .I(N__18019));
    LocalMux I__3112 (
            .O(N__18074),
            .I(N__18019));
    LocalMux I__3111 (
            .O(N__18071),
            .I(N__18014));
    LocalMux I__3110 (
            .O(N__18068),
            .I(N__18014));
    LocalMux I__3109 (
            .O(N__18065),
            .I(N__18009));
    LocalMux I__3108 (
            .O(N__18060),
            .I(N__18009));
    InMux I__3107 (
            .O(N__18057),
            .I(N__18006));
    Span4Mux_v I__3106 (
            .O(N__18054),
            .I(N__17997));
    Span4Mux_v I__3105 (
            .O(N__18051),
            .I(N__17997));
    Span4Mux_v I__3104 (
            .O(N__18048),
            .I(N__17997));
    LocalMux I__3103 (
            .O(N__18043),
            .I(N__17997));
    InMux I__3102 (
            .O(N__18042),
            .I(N__17994));
    InMux I__3101 (
            .O(N__18039),
            .I(N__17989));
    InMux I__3100 (
            .O(N__18038),
            .I(N__17989));
    LocalMux I__3099 (
            .O(N__18035),
            .I(N__17984));
    LocalMux I__3098 (
            .O(N__18032),
            .I(N__17984));
    InMux I__3097 (
            .O(N__18031),
            .I(N__17981));
    InMux I__3096 (
            .O(N__18028),
            .I(N__17978));
    InMux I__3095 (
            .O(N__18027),
            .I(N__17973));
    InMux I__3094 (
            .O(N__18026),
            .I(N__17973));
    Span4Mux_h I__3093 (
            .O(N__18019),
            .I(N__17968));
    Span4Mux_h I__3092 (
            .O(N__18014),
            .I(N__17968));
    Span4Mux_v I__3091 (
            .O(N__18009),
            .I(N__17963));
    LocalMux I__3090 (
            .O(N__18006),
            .I(N__17963));
    Odrv4 I__3089 (
            .O(N__17997),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__3088 (
            .O(N__17994),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__3087 (
            .O(N__17989),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__3086 (
            .O(N__17984),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__3085 (
            .O(N__17981),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__3084 (
            .O(N__17978),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__3083 (
            .O(N__17973),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__3082 (
            .O(N__17968),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__3081 (
            .O(N__17963),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    InMux I__3080 (
            .O(N__17944),
            .I(N__17936));
    InMux I__3079 (
            .O(N__17943),
            .I(N__17933));
    InMux I__3078 (
            .O(N__17942),
            .I(N__17930));
    InMux I__3077 (
            .O(N__17941),
            .I(N__17922));
    InMux I__3076 (
            .O(N__17940),
            .I(N__17922));
    InMux I__3075 (
            .O(N__17939),
            .I(N__17922));
    LocalMux I__3074 (
            .O(N__17936),
            .I(N__17912));
    LocalMux I__3073 (
            .O(N__17933),
            .I(N__17907));
    LocalMux I__3072 (
            .O(N__17930),
            .I(N__17907));
    InMux I__3071 (
            .O(N__17929),
            .I(N__17904));
    LocalMux I__3070 (
            .O(N__17922),
            .I(N__17898));
    InMux I__3069 (
            .O(N__17921),
            .I(N__17891));
    InMux I__3068 (
            .O(N__17920),
            .I(N__17891));
    InMux I__3067 (
            .O(N__17919),
            .I(N__17891));
    InMux I__3066 (
            .O(N__17918),
            .I(N__17888));
    CascadeMux I__3065 (
            .O(N__17917),
            .I(N__17884));
    InMux I__3064 (
            .O(N__17916),
            .I(N__17880));
    InMux I__3063 (
            .O(N__17915),
            .I(N__17877));
    Span4Mux_v I__3062 (
            .O(N__17912),
            .I(N__17870));
    Span4Mux_v I__3061 (
            .O(N__17907),
            .I(N__17870));
    LocalMux I__3060 (
            .O(N__17904),
            .I(N__17870));
    InMux I__3059 (
            .O(N__17903),
            .I(N__17863));
    InMux I__3058 (
            .O(N__17902),
            .I(N__17863));
    InMux I__3057 (
            .O(N__17901),
            .I(N__17863));
    Span4Mux_h I__3056 (
            .O(N__17898),
            .I(N__17856));
    LocalMux I__3055 (
            .O(N__17891),
            .I(N__17856));
    LocalMux I__3054 (
            .O(N__17888),
            .I(N__17856));
    InMux I__3053 (
            .O(N__17887),
            .I(N__17849));
    InMux I__3052 (
            .O(N__17884),
            .I(N__17849));
    InMux I__3051 (
            .O(N__17883),
            .I(N__17849));
    LocalMux I__3050 (
            .O(N__17880),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__3049 (
            .O(N__17877),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__3048 (
            .O(N__17870),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__3047 (
            .O(N__17863),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__3046 (
            .O(N__17856),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__3045 (
            .O(N__17849),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    InMux I__3044 (
            .O(N__17836),
            .I(N__17833));
    LocalMux I__3043 (
            .O(N__17833),
            .I(N__17830));
    Span4Mux_h I__3042 (
            .O(N__17830),
            .I(N__17827));
    Odrv4 I__3041 (
            .O(N__17827),
            .I(\this_vga_signals.g1_0_2 ));
    InMux I__3040 (
            .O(N__17824),
            .I(N__17821));
    LocalMux I__3039 (
            .O(N__17821),
            .I(\this_vga_signals.g0_0_0 ));
    InMux I__3038 (
            .O(N__17818),
            .I(N__17814));
    InMux I__3037 (
            .O(N__17817),
            .I(N__17808));
    LocalMux I__3036 (
            .O(N__17814),
            .I(N__17798));
    InMux I__3035 (
            .O(N__17813),
            .I(N__17795));
    InMux I__3034 (
            .O(N__17812),
            .I(N__17790));
    InMux I__3033 (
            .O(N__17811),
            .I(N__17790));
    LocalMux I__3032 (
            .O(N__17808),
            .I(N__17786));
    InMux I__3031 (
            .O(N__17807),
            .I(N__17781));
    InMux I__3030 (
            .O(N__17806),
            .I(N__17781));
    InMux I__3029 (
            .O(N__17805),
            .I(N__17778));
    InMux I__3028 (
            .O(N__17804),
            .I(N__17775));
    InMux I__3027 (
            .O(N__17803),
            .I(N__17772));
    InMux I__3026 (
            .O(N__17802),
            .I(N__17769));
    InMux I__3025 (
            .O(N__17801),
            .I(N__17766));
    Span4Mux_v I__3024 (
            .O(N__17798),
            .I(N__17763));
    LocalMux I__3023 (
            .O(N__17795),
            .I(N__17758));
    LocalMux I__3022 (
            .O(N__17790),
            .I(N__17758));
    InMux I__3021 (
            .O(N__17789),
            .I(N__17755));
    Span4Mux_v I__3020 (
            .O(N__17786),
            .I(N__17748));
    LocalMux I__3019 (
            .O(N__17781),
            .I(N__17748));
    LocalMux I__3018 (
            .O(N__17778),
            .I(N__17748));
    LocalMux I__3017 (
            .O(N__17775),
            .I(N__17739));
    LocalMux I__3016 (
            .O(N__17772),
            .I(N__17739));
    LocalMux I__3015 (
            .O(N__17769),
            .I(N__17739));
    LocalMux I__3014 (
            .O(N__17766),
            .I(N__17739));
    Span4Mux_h I__3013 (
            .O(N__17763),
            .I(N__17734));
    Span4Mux_v I__3012 (
            .O(N__17758),
            .I(N__17734));
    LocalMux I__3011 (
            .O(N__17755),
            .I(N__17727));
    Span4Mux_v I__3010 (
            .O(N__17748),
            .I(N__17727));
    Span4Mux_v I__3009 (
            .O(N__17739),
            .I(N__17727));
    Odrv4 I__3008 (
            .O(N__17734),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__3007 (
            .O(N__17727),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    InMux I__3006 (
            .O(N__17722),
            .I(N__17719));
    LocalMux I__3005 (
            .O(N__17719),
            .I(N__17716));
    Odrv12 I__3004 (
            .O(N__17716),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_0_0_0 ));
    InMux I__3003 (
            .O(N__17713),
            .I(N__17710));
    LocalMux I__3002 (
            .O(N__17710),
            .I(\this_vga_signals.m21_0_1 ));
    InMux I__3001 (
            .O(N__17707),
            .I(N__17704));
    LocalMux I__3000 (
            .O(N__17704),
            .I(N__17701));
    Span4Mux_h I__2999 (
            .O(N__17701),
            .I(N__17698));
    Odrv4 I__2998 (
            .O(N__17698),
            .I(\this_vga_signals.i14_mux_i ));
    CascadeMux I__2997 (
            .O(N__17695),
            .I(\this_vga_signals.N_25_0_0_cascade_ ));
    CascadeMux I__2996 (
            .O(N__17692),
            .I(\this_vga_signals.M_vcounter_q_RNITP439_0Z0Z_2_cascade_ ));
    CascadeMux I__2995 (
            .O(N__17689),
            .I(N__17686));
    InMux I__2994 (
            .O(N__17686),
            .I(N__17683));
    LocalMux I__2993 (
            .O(N__17683),
            .I(\this_vga_signals.m16_0_1 ));
    InMux I__2992 (
            .O(N__17680),
            .I(N__17669));
    InMux I__2991 (
            .O(N__17679),
            .I(N__17666));
    InMux I__2990 (
            .O(N__17678),
            .I(N__17659));
    InMux I__2989 (
            .O(N__17677),
            .I(N__17659));
    InMux I__2988 (
            .O(N__17676),
            .I(N__17659));
    InMux I__2987 (
            .O(N__17675),
            .I(N__17654));
    InMux I__2986 (
            .O(N__17674),
            .I(N__17651));
    InMux I__2985 (
            .O(N__17673),
            .I(N__17641));
    InMux I__2984 (
            .O(N__17672),
            .I(N__17641));
    LocalMux I__2983 (
            .O(N__17669),
            .I(N__17634));
    LocalMux I__2982 (
            .O(N__17666),
            .I(N__17634));
    LocalMux I__2981 (
            .O(N__17659),
            .I(N__17634));
    InMux I__2980 (
            .O(N__17658),
            .I(N__17629));
    InMux I__2979 (
            .O(N__17657),
            .I(N__17629));
    LocalMux I__2978 (
            .O(N__17654),
            .I(N__17624));
    LocalMux I__2977 (
            .O(N__17651),
            .I(N__17624));
    InMux I__2976 (
            .O(N__17650),
            .I(N__17621));
    InMux I__2975 (
            .O(N__17649),
            .I(N__17612));
    InMux I__2974 (
            .O(N__17648),
            .I(N__17612));
    InMux I__2973 (
            .O(N__17647),
            .I(N__17612));
    InMux I__2972 (
            .O(N__17646),
            .I(N__17612));
    LocalMux I__2971 (
            .O(N__17641),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i));
    Odrv4 I__2970 (
            .O(N__17634),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i));
    LocalMux I__2969 (
            .O(N__17629),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i));
    Odrv12 I__2968 (
            .O(N__17624),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i));
    LocalMux I__2967 (
            .O(N__17621),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i));
    LocalMux I__2966 (
            .O(N__17612),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i));
    InMux I__2965 (
            .O(N__17599),
            .I(N__17596));
    LocalMux I__2964 (
            .O(N__17596),
            .I(N__17590));
    InMux I__2963 (
            .O(N__17595),
            .I(N__17586));
    InMux I__2962 (
            .O(N__17594),
            .I(N__17581));
    InMux I__2961 (
            .O(N__17593),
            .I(N__17581));
    Span4Mux_h I__2960 (
            .O(N__17590),
            .I(N__17578));
    InMux I__2959 (
            .O(N__17589),
            .I(N__17575));
    LocalMux I__2958 (
            .O(N__17586),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0));
    LocalMux I__2957 (
            .O(N__17581),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0));
    Odrv4 I__2956 (
            .O(N__17578),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0));
    LocalMux I__2955 (
            .O(N__17575),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0));
    CascadeMux I__2954 (
            .O(N__17566),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_cascade_ ));
    InMux I__2953 (
            .O(N__17563),
            .I(N__17560));
    LocalMux I__2952 (
            .O(N__17560),
            .I(N__17557));
    Span4Mux_h I__2951 (
            .O(N__17557),
            .I(N__17554));
    Odrv4 I__2950 (
            .O(N__17554),
            .I(\this_vga_signals.g0_12 ));
    InMux I__2949 (
            .O(N__17551),
            .I(N__17548));
    LocalMux I__2948 (
            .O(N__17548),
            .I(\this_vga_signals.M_vcounter_q_RNITP439Z0Z_2 ));
    InMux I__2947 (
            .O(N__17545),
            .I(N__17542));
    LocalMux I__2946 (
            .O(N__17542),
            .I(N__17539));
    Odrv4 I__2945 (
            .O(N__17539),
            .I(\this_vga_signals.g2_1_1 ));
    InMux I__2944 (
            .O(N__17536),
            .I(N__17533));
    LocalMux I__2943 (
            .O(N__17533),
            .I(\this_vga_signals.g1_1_1_0 ));
    CascadeMux I__2942 (
            .O(N__17530),
            .I(N__17527));
    InMux I__2941 (
            .O(N__17527),
            .I(N__17524));
    LocalMux I__2940 (
            .O(N__17524),
            .I(N__17521));
    Odrv4 I__2939 (
            .O(N__17521),
            .I(\this_vga_signals.if_N_5_1 ));
    InMux I__2938 (
            .O(N__17518),
            .I(N__17515));
    LocalMux I__2937 (
            .O(N__17515),
            .I(\this_vga_signals.g0_5_0 ));
    CascadeMux I__2936 (
            .O(N__17512),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_cascade_ ));
    InMux I__2935 (
            .O(N__17509),
            .I(N__17505));
    CascadeMux I__2934 (
            .O(N__17508),
            .I(N__17502));
    LocalMux I__2933 (
            .O(N__17505),
            .I(N__17499));
    InMux I__2932 (
            .O(N__17502),
            .I(N__17496));
    Span4Mux_v I__2931 (
            .O(N__17499),
            .I(N__17491));
    LocalMux I__2930 (
            .O(N__17496),
            .I(N__17491));
    Span4Mux_h I__2929 (
            .O(N__17491),
            .I(N__17488));
    Span4Mux_h I__2928 (
            .O(N__17488),
            .I(N__17485));
    Odrv4 I__2927 (
            .O(N__17485),
            .I(\this_vga_signals.vaddress_2_5 ));
    CascadeMux I__2926 (
            .O(N__17482),
            .I(\this_vga_signals.g1_1_0_0_cascade_ ));
    InMux I__2925 (
            .O(N__17479),
            .I(N__17476));
    LocalMux I__2924 (
            .O(N__17476),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_0_0 ));
    InMux I__2923 (
            .O(N__17473),
            .I(N__17470));
    LocalMux I__2922 (
            .O(N__17470),
            .I(\this_vga_signals.g1_2_0_0 ));
    InMux I__2921 (
            .O(N__17467),
            .I(N__17462));
    InMux I__2920 (
            .O(N__17466),
            .I(N__17458));
    InMux I__2919 (
            .O(N__17465),
            .I(N__17455));
    LocalMux I__2918 (
            .O(N__17462),
            .I(N__17452));
    InMux I__2917 (
            .O(N__17461),
            .I(N__17449));
    LocalMux I__2916 (
            .O(N__17458),
            .I(\this_vga_signals.if_i2_mux ));
    LocalMux I__2915 (
            .O(N__17455),
            .I(\this_vga_signals.if_i2_mux ));
    Odrv4 I__2914 (
            .O(N__17452),
            .I(\this_vga_signals.if_i2_mux ));
    LocalMux I__2913 (
            .O(N__17449),
            .I(\this_vga_signals.if_i2_mux ));
    InMux I__2912 (
            .O(N__17440),
            .I(N__17437));
    LocalMux I__2911 (
            .O(N__17437),
            .I(\this_vga_signals.M_vcounter_d7lt3 ));
    InMux I__2910 (
            .O(N__17434),
            .I(N__17430));
    InMux I__2909 (
            .O(N__17433),
            .I(N__17427));
    LocalMux I__2908 (
            .O(N__17430),
            .I(N__17424));
    LocalMux I__2907 (
            .O(N__17427),
            .I(N__17421));
    Span4Mux_v I__2906 (
            .O(N__17424),
            .I(N__17416));
    Span4Mux_v I__2905 (
            .O(N__17421),
            .I(N__17416));
    Span4Mux_h I__2904 (
            .O(N__17416),
            .I(N__17413));
    Span4Mux_h I__2903 (
            .O(N__17413),
            .I(N__17410));
    Odrv4 I__2902 (
            .O(N__17410),
            .I(\this_vga_signals.M_vcounter_d7lt9_1 ));
    CascadeMux I__2901 (
            .O(N__17407),
            .I(\this_vga_signals.M_vcounter_d7lt9_1_cascade_ ));
    InMux I__2900 (
            .O(N__17404),
            .I(N__17400));
    InMux I__2899 (
            .O(N__17403),
            .I(N__17397));
    LocalMux I__2898 (
            .O(N__17400),
            .I(N__17394));
    LocalMux I__2897 (
            .O(N__17397),
            .I(N__17389));
    Span4Mux_v I__2896 (
            .O(N__17394),
            .I(N__17389));
    Odrv4 I__2895 (
            .O(N__17389),
            .I(\this_vga_signals.un4_lvisibility_1 ));
    InMux I__2894 (
            .O(N__17386),
            .I(N__17383));
    LocalMux I__2893 (
            .O(N__17383),
            .I(N__17379));
    InMux I__2892 (
            .O(N__17382),
            .I(N__17376));
    Span4Mux_v I__2891 (
            .O(N__17379),
            .I(N__17371));
    LocalMux I__2890 (
            .O(N__17376),
            .I(N__17371));
    Span4Mux_h I__2889 (
            .O(N__17371),
            .I(N__17368));
    Odrv4 I__2888 (
            .O(N__17368),
            .I(\this_vga_signals.if_m8_0_a3_1_1_0 ));
    InMux I__2887 (
            .O(N__17365),
            .I(N__17362));
    LocalMux I__2886 (
            .O(N__17362),
            .I(N__17359));
    Span4Mux_v I__2885 (
            .O(N__17359),
            .I(N__17356));
    Odrv4 I__2884 (
            .O(N__17356),
            .I(\this_vga_signals.g0_0 ));
    CascadeMux I__2883 (
            .O(N__17353),
            .I(\this_vga_signals.vaddress_1_5_cascade_ ));
    InMux I__2882 (
            .O(N__17350),
            .I(N__17347));
    LocalMux I__2881 (
            .O(N__17347),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_0_1 ));
    InMux I__2880 (
            .O(N__17344),
            .I(N__17332));
    InMux I__2879 (
            .O(N__17343),
            .I(N__17327));
    InMux I__2878 (
            .O(N__17342),
            .I(N__17324));
    InMux I__2877 (
            .O(N__17341),
            .I(N__17319));
    InMux I__2876 (
            .O(N__17340),
            .I(N__17319));
    InMux I__2875 (
            .O(N__17339),
            .I(N__17314));
    InMux I__2874 (
            .O(N__17338),
            .I(N__17314));
    InMux I__2873 (
            .O(N__17337),
            .I(N__17307));
    InMux I__2872 (
            .O(N__17336),
            .I(N__17307));
    InMux I__2871 (
            .O(N__17335),
            .I(N__17307));
    LocalMux I__2870 (
            .O(N__17332),
            .I(N__17300));
    InMux I__2869 (
            .O(N__17331),
            .I(N__17297));
    InMux I__2868 (
            .O(N__17330),
            .I(N__17294));
    LocalMux I__2867 (
            .O(N__17327),
            .I(N__17289));
    LocalMux I__2866 (
            .O(N__17324),
            .I(N__17289));
    LocalMux I__2865 (
            .O(N__17319),
            .I(N__17286));
    LocalMux I__2864 (
            .O(N__17314),
            .I(N__17283));
    LocalMux I__2863 (
            .O(N__17307),
            .I(N__17280));
    InMux I__2862 (
            .O(N__17306),
            .I(N__17275));
    InMux I__2861 (
            .O(N__17305),
            .I(N__17275));
    InMux I__2860 (
            .O(N__17304),
            .I(N__17270));
    InMux I__2859 (
            .O(N__17303),
            .I(N__17270));
    Span4Mux_h I__2858 (
            .O(N__17300),
            .I(N__17267));
    LocalMux I__2857 (
            .O(N__17297),
            .I(N__17260));
    LocalMux I__2856 (
            .O(N__17294),
            .I(N__17260));
    Span4Mux_h I__2855 (
            .O(N__17289),
            .I(N__17260));
    Span4Mux_h I__2854 (
            .O(N__17286),
            .I(N__17257));
    Odrv12 I__2853 (
            .O(N__17283),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__2852 (
            .O(N__17280),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__2851 (
            .O(N__17275),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__2850 (
            .O(N__17270),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__2849 (
            .O(N__17267),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__2848 (
            .O(N__17260),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__2847 (
            .O(N__17257),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    InMux I__2846 (
            .O(N__17242),
            .I(N__17239));
    LocalMux I__2845 (
            .O(N__17239),
            .I(\this_vga_signals.vaddress_1_5 ));
    InMux I__2844 (
            .O(N__17236),
            .I(N__17229));
    InMux I__2843 (
            .O(N__17235),
            .I(N__17226));
    InMux I__2842 (
            .O(N__17234),
            .I(N__17221));
    InMux I__2841 (
            .O(N__17233),
            .I(N__17212));
    InMux I__2840 (
            .O(N__17232),
            .I(N__17212));
    LocalMux I__2839 (
            .O(N__17229),
            .I(N__17208));
    LocalMux I__2838 (
            .O(N__17226),
            .I(N__17205));
    InMux I__2837 (
            .O(N__17225),
            .I(N__17201));
    InMux I__2836 (
            .O(N__17224),
            .I(N__17196));
    LocalMux I__2835 (
            .O(N__17221),
            .I(N__17193));
    InMux I__2834 (
            .O(N__17220),
            .I(N__17190));
    InMux I__2833 (
            .O(N__17219),
            .I(N__17183));
    InMux I__2832 (
            .O(N__17218),
            .I(N__17183));
    InMux I__2831 (
            .O(N__17217),
            .I(N__17183));
    LocalMux I__2830 (
            .O(N__17212),
            .I(N__17180));
    InMux I__2829 (
            .O(N__17211),
            .I(N__17167));
    Span4Mux_v I__2828 (
            .O(N__17208),
            .I(N__17162));
    Span4Mux_v I__2827 (
            .O(N__17205),
            .I(N__17162));
    InMux I__2826 (
            .O(N__17204),
            .I(N__17159));
    LocalMux I__2825 (
            .O(N__17201),
            .I(N__17156));
    InMux I__2824 (
            .O(N__17200),
            .I(N__17151));
    InMux I__2823 (
            .O(N__17199),
            .I(N__17151));
    LocalMux I__2822 (
            .O(N__17196),
            .I(N__17140));
    Span4Mux_h I__2821 (
            .O(N__17193),
            .I(N__17140));
    LocalMux I__2820 (
            .O(N__17190),
            .I(N__17140));
    LocalMux I__2819 (
            .O(N__17183),
            .I(N__17140));
    Span4Mux_h I__2818 (
            .O(N__17180),
            .I(N__17140));
    InMux I__2817 (
            .O(N__17179),
            .I(N__17137));
    InMux I__2816 (
            .O(N__17178),
            .I(N__17132));
    InMux I__2815 (
            .O(N__17177),
            .I(N__17132));
    InMux I__2814 (
            .O(N__17176),
            .I(N__17127));
    InMux I__2813 (
            .O(N__17175),
            .I(N__17127));
    InMux I__2812 (
            .O(N__17174),
            .I(N__17116));
    InMux I__2811 (
            .O(N__17173),
            .I(N__17116));
    InMux I__2810 (
            .O(N__17172),
            .I(N__17116));
    InMux I__2809 (
            .O(N__17171),
            .I(N__17116));
    InMux I__2808 (
            .O(N__17170),
            .I(N__17116));
    LocalMux I__2807 (
            .O(N__17167),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__2806 (
            .O(N__17162),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2805 (
            .O(N__17159),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__2804 (
            .O(N__17156),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2803 (
            .O(N__17151),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__2802 (
            .O(N__17140),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2801 (
            .O(N__17137),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2800 (
            .O(N__17132),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2799 (
            .O(N__17127),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2798 (
            .O(N__17116),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    CascadeMux I__2797 (
            .O(N__17095),
            .I(\this_vga_signals.vaddress_2_6_cascade_ ));
    InMux I__2796 (
            .O(N__17092),
            .I(N__17089));
    LocalMux I__2795 (
            .O(N__17089),
            .I(\this_vga_signals.g1_2_0 ));
    CascadeMux I__2794 (
            .O(N__17086),
            .I(M_this_vga_signals_line_clk_0_cascade_));
    CascadeMux I__2793 (
            .O(N__17083),
            .I(\this_ppu.M_state_d_0_sqmuxa_cascade_ ));
    InMux I__2792 (
            .O(N__17080),
            .I(N__17077));
    LocalMux I__2791 (
            .O(N__17077),
            .I(N__17074));
    Span4Mux_h I__2790 (
            .O(N__17074),
            .I(N__17071));
    Span4Mux_v I__2789 (
            .O(N__17071),
            .I(N__17068));
    Odrv4 I__2788 (
            .O(N__17068),
            .I(\this_sprites_ram.mem_out_bus5_2 ));
    InMux I__2787 (
            .O(N__17065),
            .I(N__17062));
    LocalMux I__2786 (
            .O(N__17062),
            .I(N__17059));
    Span12Mux_v I__2785 (
            .O(N__17059),
            .I(N__17056));
    Odrv12 I__2784 (
            .O(N__17056),
            .I(\this_sprites_ram.mem_out_bus1_2 ));
    InMux I__2783 (
            .O(N__17053),
            .I(N__17050));
    LocalMux I__2782 (
            .O(N__17050),
            .I(N__17047));
    Span12Mux_v I__2781 (
            .O(N__17047),
            .I(N__17044));
    Odrv12 I__2780 (
            .O(N__17044),
            .I(\this_sprites_ram.mem_out_bus7_1 ));
    InMux I__2779 (
            .O(N__17041),
            .I(N__17038));
    LocalMux I__2778 (
            .O(N__17038),
            .I(N__17035));
    Span12Mux_v I__2777 (
            .O(N__17035),
            .I(N__17032));
    Odrv12 I__2776 (
            .O(N__17032),
            .I(\this_sprites_ram.mem_out_bus3_1 ));
    InMux I__2775 (
            .O(N__17029),
            .I(N__17025));
    CascadeMux I__2774 (
            .O(N__17028),
            .I(N__17022));
    LocalMux I__2773 (
            .O(N__17025),
            .I(N__17019));
    InMux I__2772 (
            .O(N__17022),
            .I(N__17015));
    Span4Mux_h I__2771 (
            .O(N__17019),
            .I(N__17012));
    CascadeMux I__2770 (
            .O(N__17018),
            .I(N__17009));
    LocalMux I__2769 (
            .O(N__17015),
            .I(N__17005));
    Span4Mux_v I__2768 (
            .O(N__17012),
            .I(N__17002));
    InMux I__2767 (
            .O(N__17009),
            .I(N__16999));
    InMux I__2766 (
            .O(N__17008),
            .I(N__16996));
    Span4Mux_v I__2765 (
            .O(N__17005),
            .I(N__16993));
    Span4Mux_v I__2764 (
            .O(N__17002),
            .I(N__16988));
    LocalMux I__2763 (
            .O(N__16999),
            .I(N__16988));
    LocalMux I__2762 (
            .O(N__16996),
            .I(N__16985));
    Span4Mux_h I__2761 (
            .O(N__16993),
            .I(N__16982));
    Span4Mux_v I__2760 (
            .O(N__16988),
            .I(N__16979));
    Odrv12 I__2759 (
            .O(N__16985),
            .I(this_vga_signals_vvisibility));
    Odrv4 I__2758 (
            .O(N__16982),
            .I(this_vga_signals_vvisibility));
    Odrv4 I__2757 (
            .O(N__16979),
            .I(this_vga_signals_vvisibility));
    InMux I__2756 (
            .O(N__16972),
            .I(N__16968));
    InMux I__2755 (
            .O(N__16971),
            .I(N__16965));
    LocalMux I__2754 (
            .O(N__16968),
            .I(N__16962));
    LocalMux I__2753 (
            .O(N__16965),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0 ));
    Odrv4 I__2752 (
            .O(N__16962),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0 ));
    InMux I__2751 (
            .O(N__16957),
            .I(N__16954));
    LocalMux I__2750 (
            .O(N__16954),
            .I(N__16951));
    Span4Mux_h I__2749 (
            .O(N__16951),
            .I(N__16947));
    InMux I__2748 (
            .O(N__16950),
            .I(N__16944));
    Odrv4 I__2747 (
            .O(N__16947),
            .I(this_vga_signals_un5_vaddress_g1_1_0));
    LocalMux I__2746 (
            .O(N__16944),
            .I(this_vga_signals_un5_vaddress_g1_1_0));
    CascadeMux I__2745 (
            .O(N__16939),
            .I(N__16936));
    InMux I__2744 (
            .O(N__16936),
            .I(N__16933));
    LocalMux I__2743 (
            .O(N__16933),
            .I(N__16930));
    Span4Mux_h I__2742 (
            .O(N__16930),
            .I(N__16927));
    Odrv4 I__2741 (
            .O(N__16927),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_0 ));
    InMux I__2740 (
            .O(N__16924),
            .I(N__16921));
    LocalMux I__2739 (
            .O(N__16921),
            .I(\this_vga_signals.g1_2 ));
    InMux I__2738 (
            .O(N__16918),
            .I(N__16915));
    LocalMux I__2737 (
            .O(N__16915),
            .I(\this_vga_signals.m21_0_1_1 ));
    InMux I__2736 (
            .O(N__16912),
            .I(N__16909));
    LocalMux I__2735 (
            .O(N__16909),
            .I(N__16906));
    Span4Mux_h I__2734 (
            .O(N__16906),
            .I(N__16903));
    Odrv4 I__2733 (
            .O(N__16903),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ));
    InMux I__2732 (
            .O(N__16900),
            .I(N__16897));
    LocalMux I__2731 (
            .O(N__16897),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ));
    InMux I__2730 (
            .O(N__16894),
            .I(N__16891));
    LocalMux I__2729 (
            .O(N__16891),
            .I(N__16888));
    Span4Mux_v I__2728 (
            .O(N__16888),
            .I(N__16885));
    Sp12to4 I__2727 (
            .O(N__16885),
            .I(N__16882));
    Odrv12 I__2726 (
            .O(N__16882),
            .I(M_this_ppu_vram_data_0));
    InMux I__2725 (
            .O(N__16879),
            .I(N__16876));
    LocalMux I__2724 (
            .O(N__16876),
            .I(\this_vga_ramdac.m16 ));
    InMux I__2723 (
            .O(N__16873),
            .I(N__16870));
    LocalMux I__2722 (
            .O(N__16870),
            .I(N__16865));
    InMux I__2721 (
            .O(N__16869),
            .I(N__16862));
    InMux I__2720 (
            .O(N__16868),
            .I(N__16859));
    Span4Mux_v I__2719 (
            .O(N__16865),
            .I(N__16856));
    LocalMux I__2718 (
            .O(N__16862),
            .I(N__16851));
    LocalMux I__2717 (
            .O(N__16859),
            .I(N__16848));
    Sp12to4 I__2716 (
            .O(N__16856),
            .I(N__16845));
    InMux I__2715 (
            .O(N__16855),
            .I(N__16840));
    InMux I__2714 (
            .O(N__16854),
            .I(N__16840));
    Sp12to4 I__2713 (
            .O(N__16851),
            .I(N__16837));
    Span12Mux_v I__2712 (
            .O(N__16848),
            .I(N__16832));
    Span12Mux_s3_h I__2711 (
            .O(N__16845),
            .I(N__16832));
    LocalMux I__2710 (
            .O(N__16840),
            .I(N__16827));
    Span12Mux_v I__2709 (
            .O(N__16837),
            .I(N__16827));
    Span12Mux_h I__2708 (
            .O(N__16832),
            .I(N__16824));
    Span12Mux_h I__2707 (
            .O(N__16827),
            .I(N__16821));
    Odrv12 I__2706 (
            .O(N__16824),
            .I(M_this_vram_read_data_2));
    Odrv12 I__2705 (
            .O(N__16821),
            .I(M_this_vram_read_data_2));
    InMux I__2704 (
            .O(N__16816),
            .I(N__16811));
    InMux I__2703 (
            .O(N__16815),
            .I(N__16808));
    InMux I__2702 (
            .O(N__16814),
            .I(N__16805));
    LocalMux I__2701 (
            .O(N__16811),
            .I(N__16800));
    LocalMux I__2700 (
            .O(N__16808),
            .I(N__16795));
    LocalMux I__2699 (
            .O(N__16805),
            .I(N__16795));
    CascadeMux I__2698 (
            .O(N__16804),
            .I(N__16792));
    InMux I__2697 (
            .O(N__16803),
            .I(N__16788));
    Span4Mux_v I__2696 (
            .O(N__16800),
            .I(N__16785));
    Span4Mux_v I__2695 (
            .O(N__16795),
            .I(N__16782));
    InMux I__2694 (
            .O(N__16792),
            .I(N__16777));
    InMux I__2693 (
            .O(N__16791),
            .I(N__16777));
    LocalMux I__2692 (
            .O(N__16788),
            .I(N__16774));
    Sp12to4 I__2691 (
            .O(N__16785),
            .I(N__16769));
    Sp12to4 I__2690 (
            .O(N__16782),
            .I(N__16769));
    LocalMux I__2689 (
            .O(N__16777),
            .I(N__16764));
    Span12Mux_v I__2688 (
            .O(N__16774),
            .I(N__16764));
    Span12Mux_h I__2687 (
            .O(N__16769),
            .I(N__16761));
    Span12Mux_h I__2686 (
            .O(N__16764),
            .I(N__16758));
    Odrv12 I__2685 (
            .O(N__16761),
            .I(M_this_vram_read_data_1));
    Odrv12 I__2684 (
            .O(N__16758),
            .I(M_this_vram_read_data_1));
    InMux I__2683 (
            .O(N__16753),
            .I(N__16748));
    CascadeMux I__2682 (
            .O(N__16752),
            .I(N__16744));
    InMux I__2681 (
            .O(N__16751),
            .I(N__16740));
    LocalMux I__2680 (
            .O(N__16748),
            .I(N__16736));
    InMux I__2679 (
            .O(N__16747),
            .I(N__16733));
    InMux I__2678 (
            .O(N__16744),
            .I(N__16728));
    InMux I__2677 (
            .O(N__16743),
            .I(N__16728));
    LocalMux I__2676 (
            .O(N__16740),
            .I(N__16725));
    InMux I__2675 (
            .O(N__16739),
            .I(N__16722));
    Span4Mux_h I__2674 (
            .O(N__16736),
            .I(N__16717));
    LocalMux I__2673 (
            .O(N__16733),
            .I(N__16717));
    LocalMux I__2672 (
            .O(N__16728),
            .I(N__16714));
    Span4Mux_h I__2671 (
            .O(N__16725),
            .I(N__16711));
    LocalMux I__2670 (
            .O(N__16722),
            .I(N__16706));
    Span4Mux_h I__2669 (
            .O(N__16717),
            .I(N__16706));
    Span4Mux_v I__2668 (
            .O(N__16714),
            .I(N__16701));
    Span4Mux_h I__2667 (
            .O(N__16711),
            .I(N__16701));
    Span4Mux_h I__2666 (
            .O(N__16706),
            .I(N__16698));
    Span4Mux_h I__2665 (
            .O(N__16701),
            .I(N__16695));
    Sp12to4 I__2664 (
            .O(N__16698),
            .I(N__16692));
    Span4Mux_h I__2663 (
            .O(N__16695),
            .I(N__16689));
    Span12Mux_v I__2662 (
            .O(N__16692),
            .I(N__16686));
    Span4Mux_h I__2661 (
            .O(N__16689),
            .I(N__16683));
    Odrv12 I__2660 (
            .O(N__16686),
            .I(M_this_vram_read_data_0));
    Odrv4 I__2659 (
            .O(N__16683),
            .I(M_this_vram_read_data_0));
    CascadeMux I__2658 (
            .O(N__16678),
            .I(N__16675));
    InMux I__2657 (
            .O(N__16675),
            .I(N__16670));
    CascadeMux I__2656 (
            .O(N__16674),
            .I(N__16667));
    CascadeMux I__2655 (
            .O(N__16673),
            .I(N__16663));
    LocalMux I__2654 (
            .O(N__16670),
            .I(N__16660));
    InMux I__2653 (
            .O(N__16667),
            .I(N__16657));
    InMux I__2652 (
            .O(N__16666),
            .I(N__16654));
    InMux I__2651 (
            .O(N__16663),
            .I(N__16651));
    Span4Mux_h I__2650 (
            .O(N__16660),
            .I(N__16646));
    LocalMux I__2649 (
            .O(N__16657),
            .I(N__16646));
    LocalMux I__2648 (
            .O(N__16654),
            .I(N__16641));
    LocalMux I__2647 (
            .O(N__16651),
            .I(N__16636));
    Span4Mux_h I__2646 (
            .O(N__16646),
            .I(N__16636));
    InMux I__2645 (
            .O(N__16645),
            .I(N__16631));
    InMux I__2644 (
            .O(N__16644),
            .I(N__16631));
    Span4Mux_v I__2643 (
            .O(N__16641),
            .I(N__16628));
    Span4Mux_h I__2642 (
            .O(N__16636),
            .I(N__16625));
    LocalMux I__2641 (
            .O(N__16631),
            .I(N__16622));
    Sp12to4 I__2640 (
            .O(N__16628),
            .I(N__16619));
    Span4Mux_h I__2639 (
            .O(N__16625),
            .I(N__16616));
    Span4Mux_h I__2638 (
            .O(N__16622),
            .I(N__16613));
    Span12Mux_s4_h I__2637 (
            .O(N__16619),
            .I(N__16610));
    Span4Mux_h I__2636 (
            .O(N__16616),
            .I(N__16607));
    Sp12to4 I__2635 (
            .O(N__16613),
            .I(N__16602));
    Span12Mux_h I__2634 (
            .O(N__16610),
            .I(N__16602));
    Span4Mux_h I__2633 (
            .O(N__16607),
            .I(N__16599));
    Odrv12 I__2632 (
            .O(N__16602),
            .I(M_this_vram_read_data_3));
    Odrv4 I__2631 (
            .O(N__16599),
            .I(M_this_vram_read_data_3));
    InMux I__2630 (
            .O(N__16594),
            .I(N__16591));
    LocalMux I__2629 (
            .O(N__16591),
            .I(\this_vga_ramdac.i2_mux ));
    InMux I__2628 (
            .O(N__16588),
            .I(N__16579));
    InMux I__2627 (
            .O(N__16587),
            .I(N__16579));
    InMux I__2626 (
            .O(N__16586),
            .I(N__16575));
    InMux I__2625 (
            .O(N__16585),
            .I(N__16572));
    InMux I__2624 (
            .O(N__16584),
            .I(N__16567));
    LocalMux I__2623 (
            .O(N__16579),
            .I(N__16564));
    InMux I__2622 (
            .O(N__16578),
            .I(N__16561));
    LocalMux I__2621 (
            .O(N__16575),
            .I(N__16557));
    LocalMux I__2620 (
            .O(N__16572),
            .I(N__16554));
    InMux I__2619 (
            .O(N__16571),
            .I(N__16551));
    InMux I__2618 (
            .O(N__16570),
            .I(N__16548));
    LocalMux I__2617 (
            .O(N__16567),
            .I(N__16545));
    Span4Mux_v I__2616 (
            .O(N__16564),
            .I(N__16540));
    LocalMux I__2615 (
            .O(N__16561),
            .I(N__16540));
    InMux I__2614 (
            .O(N__16560),
            .I(N__16535));
    Span4Mux_v I__2613 (
            .O(N__16557),
            .I(N__16530));
    Span4Mux_v I__2612 (
            .O(N__16554),
            .I(N__16530));
    LocalMux I__2611 (
            .O(N__16551),
            .I(N__16525));
    LocalMux I__2610 (
            .O(N__16548),
            .I(N__16525));
    Span4Mux_v I__2609 (
            .O(N__16545),
            .I(N__16520));
    Span4Mux_h I__2608 (
            .O(N__16540),
            .I(N__16520));
    InMux I__2607 (
            .O(N__16539),
            .I(N__16515));
    InMux I__2606 (
            .O(N__16538),
            .I(N__16515));
    LocalMux I__2605 (
            .O(N__16535),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2604 (
            .O(N__16530),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv12 I__2603 (
            .O(N__16525),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2602 (
            .O(N__16520),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2601 (
            .O(N__16515),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    CascadeMux I__2600 (
            .O(N__16504),
            .I(N__16495));
    CascadeMux I__2599 (
            .O(N__16503),
            .I(N__16491));
    InMux I__2598 (
            .O(N__16502),
            .I(N__16488));
    InMux I__2597 (
            .O(N__16501),
            .I(N__16485));
    InMux I__2596 (
            .O(N__16500),
            .I(N__16482));
    InMux I__2595 (
            .O(N__16499),
            .I(N__16479));
    InMux I__2594 (
            .O(N__16498),
            .I(N__16476));
    InMux I__2593 (
            .O(N__16495),
            .I(N__16473));
    InMux I__2592 (
            .O(N__16494),
            .I(N__16470));
    InMux I__2591 (
            .O(N__16491),
            .I(N__16464));
    LocalMux I__2590 (
            .O(N__16488),
            .I(N__16461));
    LocalMux I__2589 (
            .O(N__16485),
            .I(N__16456));
    LocalMux I__2588 (
            .O(N__16482),
            .I(N__16456));
    LocalMux I__2587 (
            .O(N__16479),
            .I(N__16449));
    LocalMux I__2586 (
            .O(N__16476),
            .I(N__16449));
    LocalMux I__2585 (
            .O(N__16473),
            .I(N__16449));
    LocalMux I__2584 (
            .O(N__16470),
            .I(N__16446));
    InMux I__2583 (
            .O(N__16469),
            .I(N__16443));
    CascadeMux I__2582 (
            .O(N__16468),
            .I(N__16439));
    InMux I__2581 (
            .O(N__16467),
            .I(N__16436));
    LocalMux I__2580 (
            .O(N__16464),
            .I(N__16433));
    Span4Mux_h I__2579 (
            .O(N__16461),
            .I(N__16430));
    Span4Mux_h I__2578 (
            .O(N__16456),
            .I(N__16425));
    Span4Mux_v I__2577 (
            .O(N__16449),
            .I(N__16425));
    Span4Mux_v I__2576 (
            .O(N__16446),
            .I(N__16420));
    LocalMux I__2575 (
            .O(N__16443),
            .I(N__16420));
    InMux I__2574 (
            .O(N__16442),
            .I(N__16415));
    InMux I__2573 (
            .O(N__16439),
            .I(N__16415));
    LocalMux I__2572 (
            .O(N__16436),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2571 (
            .O(N__16433),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2570 (
            .O(N__16430),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2569 (
            .O(N__16425),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2568 (
            .O(N__16420),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2567 (
            .O(N__16415),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    CascadeMux I__2566 (
            .O(N__16402),
            .I(N__16399));
    InMux I__2565 (
            .O(N__16399),
            .I(N__16396));
    LocalMux I__2564 (
            .O(N__16396),
            .I(N__16392));
    InMux I__2563 (
            .O(N__16395),
            .I(N__16389));
    Odrv4 I__2562 (
            .O(N__16392),
            .I(\this_vga_signals.line_clk_1 ));
    LocalMux I__2561 (
            .O(N__16389),
            .I(\this_vga_signals.line_clk_1 ));
    InMux I__2560 (
            .O(N__16384),
            .I(N__16381));
    LocalMux I__2559 (
            .O(N__16381),
            .I(N__16378));
    Odrv4 I__2558 (
            .O(N__16378),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    InMux I__2557 (
            .O(N__16375),
            .I(N__16372));
    LocalMux I__2556 (
            .O(N__16372),
            .I(N__16369));
    Odrv4 I__2555 (
            .O(N__16369),
            .I(\this_vga_signals.g0_2_0_2 ));
    InMux I__2554 (
            .O(N__16366),
            .I(N__16363));
    LocalMux I__2553 (
            .O(N__16363),
            .I(\this_vga_signals.g1_0_0_0_1 ));
    InMux I__2552 (
            .O(N__16360),
            .I(N__16357));
    LocalMux I__2551 (
            .O(N__16357),
            .I(\this_vga_signals.N_51 ));
    InMux I__2550 (
            .O(N__16354),
            .I(N__16351));
    LocalMux I__2549 (
            .O(N__16351),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_0 ));
    InMux I__2548 (
            .O(N__16348),
            .I(N__16344));
    InMux I__2547 (
            .O(N__16347),
            .I(N__16341));
    LocalMux I__2546 (
            .O(N__16344),
            .I(N__16338));
    LocalMux I__2545 (
            .O(N__16341),
            .I(N__16335));
    Span4Mux_h I__2544 (
            .O(N__16338),
            .I(N__16332));
    Odrv4 I__2543 (
            .O(N__16335),
            .I(\this_vga_signals.g2_1 ));
    Odrv4 I__2542 (
            .O(N__16332),
            .I(\this_vga_signals.g2_1 ));
    InMux I__2541 (
            .O(N__16327),
            .I(N__16324));
    LocalMux I__2540 (
            .O(N__16324),
            .I(N__16321));
    Odrv4 I__2539 (
            .O(N__16321),
            .I(\this_vga_signals.g1_0 ));
    CascadeMux I__2538 (
            .O(N__16318),
            .I(\this_vga_signals.g1_N_4L5_1_cascade_ ));
    CascadeMux I__2537 (
            .O(N__16315),
            .I(\this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5EZ0Z1_cascade_ ));
    InMux I__2536 (
            .O(N__16312),
            .I(N__16303));
    InMux I__2535 (
            .O(N__16311),
            .I(N__16303));
    InMux I__2534 (
            .O(N__16310),
            .I(N__16298));
    InMux I__2533 (
            .O(N__16309),
            .I(N__16298));
    InMux I__2532 (
            .O(N__16308),
            .I(N__16295));
    LocalMux I__2531 (
            .O(N__16303),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    LocalMux I__2530 (
            .O(N__16298),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    LocalMux I__2529 (
            .O(N__16295),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    InMux I__2528 (
            .O(N__16288),
            .I(N__16285));
    LocalMux I__2527 (
            .O(N__16285),
            .I(\this_vga_signals.g0_1_1 ));
    CascadeMux I__2526 (
            .O(N__16282),
            .I(N__16277));
    InMux I__2525 (
            .O(N__16281),
            .I(N__16274));
    InMux I__2524 (
            .O(N__16280),
            .I(N__16271));
    InMux I__2523 (
            .O(N__16277),
            .I(N__16268));
    LocalMux I__2522 (
            .O(N__16274),
            .I(\this_vga_signals.d_N_3_0_i ));
    LocalMux I__2521 (
            .O(N__16271),
            .I(\this_vga_signals.d_N_3_0_i ));
    LocalMux I__2520 (
            .O(N__16268),
            .I(\this_vga_signals.d_N_3_0_i ));
    InMux I__2519 (
            .O(N__16261),
            .I(N__16258));
    LocalMux I__2518 (
            .O(N__16258),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_x0 ));
    CascadeMux I__2517 (
            .O(N__16255),
            .I(\this_vga_signals.mult1_un61_sum_c3_cascade_ ));
    InMux I__2516 (
            .O(N__16252),
            .I(N__16249));
    LocalMux I__2515 (
            .O(N__16249),
            .I(\this_vga_signals.g0_7 ));
    InMux I__2514 (
            .O(N__16246),
            .I(N__16243));
    LocalMux I__2513 (
            .O(N__16243),
            .I(\this_vga_signals.g2_2 ));
    InMux I__2512 (
            .O(N__16240),
            .I(N__16237));
    LocalMux I__2511 (
            .O(N__16237),
            .I(m18x_N_3LZ0Z3));
    InMux I__2510 (
            .O(N__16234),
            .I(N__16231));
    LocalMux I__2509 (
            .O(N__16231),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI5BS7NZ0Z_5 ));
    CascadeMux I__2508 (
            .O(N__16228),
            .I(N__16225));
    InMux I__2507 (
            .O(N__16225),
            .I(N__16221));
    InMux I__2506 (
            .O(N__16224),
            .I(N__16218));
    LocalMux I__2505 (
            .O(N__16221),
            .I(N__16213));
    LocalMux I__2504 (
            .O(N__16218),
            .I(N__16213));
    Odrv4 I__2503 (
            .O(N__16213),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_0_0 ));
    CascadeMux I__2502 (
            .O(N__16210),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0_x0_cascade_ ));
    CascadeMux I__2501 (
            .O(N__16207),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0_cascade_ ));
    InMux I__2500 (
            .O(N__16204),
            .I(N__16201));
    LocalMux I__2499 (
            .O(N__16201),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0_x1 ));
    InMux I__2498 (
            .O(N__16198),
            .I(N__16195));
    LocalMux I__2497 (
            .O(N__16195),
            .I(N__16192));
    Span4Mux_h I__2496 (
            .O(N__16192),
            .I(N__16189));
    Span4Mux_v I__2495 (
            .O(N__16189),
            .I(N__16186));
    Odrv4 I__2494 (
            .O(N__16186),
            .I(\this_vga_signals.vaddress_4_5 ));
    InMux I__2493 (
            .O(N__16183),
            .I(N__16180));
    LocalMux I__2492 (
            .O(N__16180),
            .I(N__16175));
    CascadeMux I__2491 (
            .O(N__16179),
            .I(N__16172));
    CascadeMux I__2490 (
            .O(N__16178),
            .I(N__16169));
    Span4Mux_h I__2489 (
            .O(N__16175),
            .I(N__16163));
    InMux I__2488 (
            .O(N__16172),
            .I(N__16158));
    InMux I__2487 (
            .O(N__16169),
            .I(N__16158));
    InMux I__2486 (
            .O(N__16168),
            .I(N__16155));
    InMux I__2485 (
            .O(N__16167),
            .I(N__16150));
    InMux I__2484 (
            .O(N__16166),
            .I(N__16150));
    Odrv4 I__2483 (
            .O(N__16163),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__2482 (
            .O(N__16158),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__2481 (
            .O(N__16155),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__2480 (
            .O(N__16150),
            .I(\this_vga_signals.vaddress_5 ));
    CascadeMux I__2479 (
            .O(N__16141),
            .I(N__16131));
    InMux I__2478 (
            .O(N__16140),
            .I(N__16128));
    InMux I__2477 (
            .O(N__16139),
            .I(N__16123));
    InMux I__2476 (
            .O(N__16138),
            .I(N__16123));
    InMux I__2475 (
            .O(N__16137),
            .I(N__16118));
    InMux I__2474 (
            .O(N__16136),
            .I(N__16118));
    InMux I__2473 (
            .O(N__16135),
            .I(N__16113));
    InMux I__2472 (
            .O(N__16134),
            .I(N__16113));
    InMux I__2471 (
            .O(N__16131),
            .I(N__16110));
    LocalMux I__2470 (
            .O(N__16128),
            .I(N__16107));
    LocalMux I__2469 (
            .O(N__16123),
            .I(N__16104));
    LocalMux I__2468 (
            .O(N__16118),
            .I(N__16099));
    LocalMux I__2467 (
            .O(N__16113),
            .I(N__16099));
    LocalMux I__2466 (
            .O(N__16110),
            .I(N__16092));
    Span4Mux_h I__2465 (
            .O(N__16107),
            .I(N__16092));
    Span4Mux_v I__2464 (
            .O(N__16104),
            .I(N__16092));
    Odrv4 I__2463 (
            .O(N__16099),
            .I(\this_vga_signals.vaddress_6 ));
    Odrv4 I__2462 (
            .O(N__16092),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__2461 (
            .O(N__16087),
            .I(N__16084));
    LocalMux I__2460 (
            .O(N__16084),
            .I(N__16081));
    Odrv4 I__2459 (
            .O(N__16081),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_0 ));
    CascadeMux I__2458 (
            .O(N__16078),
            .I(\this_vga_signals.mult1_un47_sum_c3_cascade_ ));
    InMux I__2457 (
            .O(N__16075),
            .I(N__16072));
    LocalMux I__2456 (
            .O(N__16072),
            .I(\this_vga_signals.N_5_i_0_0 ));
    CascadeMux I__2455 (
            .O(N__16069),
            .I(N__16066));
    InMux I__2454 (
            .O(N__16066),
            .I(N__16063));
    LocalMux I__2453 (
            .O(N__16063),
            .I(\this_vga_signals.i2_mux ));
    CascadeMux I__2452 (
            .O(N__16060),
            .I(\this_vga_signals.i2_mux_cascade_ ));
    CascadeMux I__2451 (
            .O(N__16057),
            .I(\this_vga_signals.if_i2_mux_cascade_ ));
    InMux I__2450 (
            .O(N__16054),
            .I(N__16051));
    LocalMux I__2449 (
            .O(N__16051),
            .I(N__16047));
    InMux I__2448 (
            .O(N__16050),
            .I(N__16044));
    Span4Mux_v I__2447 (
            .O(N__16047),
            .I(N__16041));
    LocalMux I__2446 (
            .O(N__16044),
            .I(N__16036));
    Span4Mux_h I__2445 (
            .O(N__16041),
            .I(N__16036));
    Odrv4 I__2444 (
            .O(N__16036),
            .I(\this_vga_signals.vaddress_0_6 ));
    InMux I__2443 (
            .O(N__16033),
            .I(N__16026));
    InMux I__2442 (
            .O(N__16032),
            .I(N__16026));
    InMux I__2441 (
            .O(N__16031),
            .I(N__16023));
    LocalMux I__2440 (
            .O(N__16026),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    LocalMux I__2439 (
            .O(N__16023),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    InMux I__2438 (
            .O(N__16018),
            .I(N__16013));
    InMux I__2437 (
            .O(N__16017),
            .I(N__16010));
    InMux I__2436 (
            .O(N__16016),
            .I(N__16007));
    LocalMux I__2435 (
            .O(N__16013),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    LocalMux I__2434 (
            .O(N__16010),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    LocalMux I__2433 (
            .O(N__16007),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    InMux I__2432 (
            .O(N__16000),
            .I(N__15991));
    InMux I__2431 (
            .O(N__15999),
            .I(N__15987));
    InMux I__2430 (
            .O(N__15998),
            .I(N__15984));
    InMux I__2429 (
            .O(N__15997),
            .I(N__15981));
    InMux I__2428 (
            .O(N__15996),
            .I(N__15976));
    InMux I__2427 (
            .O(N__15995),
            .I(N__15976));
    InMux I__2426 (
            .O(N__15994),
            .I(N__15972));
    LocalMux I__2425 (
            .O(N__15991),
            .I(N__15969));
    InMux I__2424 (
            .O(N__15990),
            .I(N__15966));
    LocalMux I__2423 (
            .O(N__15987),
            .I(N__15961));
    LocalMux I__2422 (
            .O(N__15984),
            .I(N__15955));
    LocalMux I__2421 (
            .O(N__15981),
            .I(N__15955));
    LocalMux I__2420 (
            .O(N__15976),
            .I(N__15952));
    InMux I__2419 (
            .O(N__15975),
            .I(N__15949));
    LocalMux I__2418 (
            .O(N__15972),
            .I(N__15942));
    Span4Mux_h I__2417 (
            .O(N__15969),
            .I(N__15942));
    LocalMux I__2416 (
            .O(N__15966),
            .I(N__15942));
    InMux I__2415 (
            .O(N__15965),
            .I(N__15939));
    InMux I__2414 (
            .O(N__15964),
            .I(N__15932));
    Span12Mux_v I__2413 (
            .O(N__15961),
            .I(N__15929));
    InMux I__2412 (
            .O(N__15960),
            .I(N__15926));
    Span4Mux_v I__2411 (
            .O(N__15955),
            .I(N__15921));
    Span4Mux_v I__2410 (
            .O(N__15952),
            .I(N__15921));
    LocalMux I__2409 (
            .O(N__15949),
            .I(N__15914));
    Span4Mux_v I__2408 (
            .O(N__15942),
            .I(N__15914));
    LocalMux I__2407 (
            .O(N__15939),
            .I(N__15914));
    InMux I__2406 (
            .O(N__15938),
            .I(N__15911));
    InMux I__2405 (
            .O(N__15937),
            .I(N__15908));
    InMux I__2404 (
            .O(N__15936),
            .I(N__15903));
    InMux I__2403 (
            .O(N__15935),
            .I(N__15903));
    LocalMux I__2402 (
            .O(N__15932),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv12 I__2401 (
            .O(N__15929),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2400 (
            .O(N__15926),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__2399 (
            .O(N__15921),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__2398 (
            .O(N__15914),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2397 (
            .O(N__15911),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2396 (
            .O(N__15908),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2395 (
            .O(N__15903),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    InMux I__2394 (
            .O(N__15886),
            .I(N__15882));
    InMux I__2393 (
            .O(N__15885),
            .I(N__15879));
    LocalMux I__2392 (
            .O(N__15882),
            .I(N__15876));
    LocalMux I__2391 (
            .O(N__15879),
            .I(N__15871));
    Span4Mux_v I__2390 (
            .O(N__15876),
            .I(N__15868));
    InMux I__2389 (
            .O(N__15875),
            .I(N__15863));
    InMux I__2388 (
            .O(N__15874),
            .I(N__15863));
    Span12Mux_s5_h I__2387 (
            .O(N__15871),
            .I(N__15858));
    Span4Mux_h I__2386 (
            .O(N__15868),
            .I(N__15853));
    LocalMux I__2385 (
            .O(N__15863),
            .I(N__15853));
    InMux I__2384 (
            .O(N__15862),
            .I(N__15848));
    InMux I__2383 (
            .O(N__15861),
            .I(N__15848));
    Odrv12 I__2382 (
            .O(N__15858),
            .I(G_384));
    Odrv4 I__2381 (
            .O(N__15853),
            .I(G_384));
    LocalMux I__2380 (
            .O(N__15848),
            .I(G_384));
    InMux I__2379 (
            .O(N__15841),
            .I(N__15838));
    LocalMux I__2378 (
            .O(N__15838),
            .I(N__15835));
    Span4Mux_v I__2377 (
            .O(N__15835),
            .I(N__15831));
    CascadeMux I__2376 (
            .O(N__15834),
            .I(N__15828));
    Span4Mux_h I__2375 (
            .O(N__15831),
            .I(N__15825));
    InMux I__2374 (
            .O(N__15828),
            .I(N__15822));
    Odrv4 I__2373 (
            .O(N__15825),
            .I(\this_vga_ramdac.N_2873_reto ));
    LocalMux I__2372 (
            .O(N__15822),
            .I(\this_vga_ramdac.N_2873_reto ));
    InMux I__2371 (
            .O(N__15817),
            .I(N__15811));
    InMux I__2370 (
            .O(N__15816),
            .I(N__15811));
    LocalMux I__2369 (
            .O(N__15811),
            .I(N_3_0));
    InMux I__2368 (
            .O(N__15808),
            .I(N__15802));
    InMux I__2367 (
            .O(N__15807),
            .I(N__15802));
    LocalMux I__2366 (
            .O(N__15802),
            .I(N_2_0));
    InMux I__2365 (
            .O(N__15799),
            .I(N__15796));
    LocalMux I__2364 (
            .O(N__15796),
            .I(M_this_vga_signals_pixel_clk_0_0));
    CEMux I__2363 (
            .O(N__15793),
            .I(N__15789));
    CEMux I__2362 (
            .O(N__15792),
            .I(N__15786));
    LocalMux I__2361 (
            .O(N__15789),
            .I(N__15783));
    LocalMux I__2360 (
            .O(N__15786),
            .I(N__15780));
    Span4Mux_v I__2359 (
            .O(N__15783),
            .I(N__15777));
    Span4Mux_h I__2358 (
            .O(N__15780),
            .I(N__15774));
    Span4Mux_v I__2357 (
            .O(N__15777),
            .I(N__15771));
    Span4Mux_v I__2356 (
            .O(N__15774),
            .I(N__15768));
    Odrv4 I__2355 (
            .O(N__15771),
            .I(\this_sprites_ram.mem_WE_2 ));
    Odrv4 I__2354 (
            .O(N__15768),
            .I(\this_sprites_ram.mem_WE_2 ));
    CascadeMux I__2353 (
            .O(N__15763),
            .I(N__15760));
    CascadeBuf I__2352 (
            .O(N__15760),
            .I(N__15757));
    CascadeMux I__2351 (
            .O(N__15757),
            .I(N__15754));
    CascadeBuf I__2350 (
            .O(N__15754),
            .I(N__15751));
    CascadeMux I__2349 (
            .O(N__15751),
            .I(N__15748));
    CascadeBuf I__2348 (
            .O(N__15748),
            .I(N__15745));
    CascadeMux I__2347 (
            .O(N__15745),
            .I(N__15742));
    CascadeBuf I__2346 (
            .O(N__15742),
            .I(N__15739));
    CascadeMux I__2345 (
            .O(N__15739),
            .I(N__15736));
    CascadeBuf I__2344 (
            .O(N__15736),
            .I(N__15733));
    CascadeMux I__2343 (
            .O(N__15733),
            .I(N__15730));
    CascadeBuf I__2342 (
            .O(N__15730),
            .I(N__15727));
    CascadeMux I__2341 (
            .O(N__15727),
            .I(N__15724));
    CascadeBuf I__2340 (
            .O(N__15724),
            .I(N__15721));
    CascadeMux I__2339 (
            .O(N__15721),
            .I(N__15718));
    CascadeBuf I__2338 (
            .O(N__15718),
            .I(N__15715));
    CascadeMux I__2337 (
            .O(N__15715),
            .I(N__15712));
    CascadeBuf I__2336 (
            .O(N__15712),
            .I(N__15709));
    CascadeMux I__2335 (
            .O(N__15709),
            .I(N__15706));
    CascadeBuf I__2334 (
            .O(N__15706),
            .I(N__15703));
    CascadeMux I__2333 (
            .O(N__15703),
            .I(N__15700));
    CascadeBuf I__2332 (
            .O(N__15700),
            .I(N__15697));
    CascadeMux I__2331 (
            .O(N__15697),
            .I(N__15694));
    CascadeBuf I__2330 (
            .O(N__15694),
            .I(N__15691));
    CascadeMux I__2329 (
            .O(N__15691),
            .I(N__15688));
    CascadeBuf I__2328 (
            .O(N__15688),
            .I(N__15685));
    CascadeMux I__2327 (
            .O(N__15685),
            .I(N__15682));
    CascadeBuf I__2326 (
            .O(N__15682),
            .I(N__15678));
    CascadeMux I__2325 (
            .O(N__15681),
            .I(N__15675));
    CascadeMux I__2324 (
            .O(N__15678),
            .I(N__15672));
    InMux I__2323 (
            .O(N__15675),
            .I(N__15669));
    CascadeBuf I__2322 (
            .O(N__15672),
            .I(N__15666));
    LocalMux I__2321 (
            .O(N__15669),
            .I(N__15663));
    CascadeMux I__2320 (
            .O(N__15666),
            .I(N__15660));
    Span4Mux_v I__2319 (
            .O(N__15663),
            .I(N__15656));
    InMux I__2318 (
            .O(N__15660),
            .I(N__15652));
    InMux I__2317 (
            .O(N__15659),
            .I(N__15649));
    Sp12to4 I__2316 (
            .O(N__15656),
            .I(N__15644));
    InMux I__2315 (
            .O(N__15655),
            .I(N__15641));
    LocalMux I__2314 (
            .O(N__15652),
            .I(N__15638));
    LocalMux I__2313 (
            .O(N__15649),
            .I(N__15635));
    InMux I__2312 (
            .O(N__15648),
            .I(N__15630));
    InMux I__2311 (
            .O(N__15647),
            .I(N__15630));
    Span12Mux_h I__2310 (
            .O(N__15644),
            .I(N__15627));
    LocalMux I__2309 (
            .O(N__15641),
            .I(N__15622));
    Span12Mux_s10_h I__2308 (
            .O(N__15638),
            .I(N__15622));
    Odrv4 I__2307 (
            .O(N__15635),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__2306 (
            .O(N__15630),
            .I(M_this_ppu_vram_addr_7));
    Odrv12 I__2305 (
            .O(N__15627),
            .I(M_this_ppu_vram_addr_7));
    Odrv12 I__2304 (
            .O(N__15622),
            .I(M_this_ppu_vram_addr_7));
    CascadeMux I__2303 (
            .O(N__15613),
            .I(N__15610));
    CascadeBuf I__2302 (
            .O(N__15610),
            .I(N__15607));
    CascadeMux I__2301 (
            .O(N__15607),
            .I(N__15604));
    CascadeBuf I__2300 (
            .O(N__15604),
            .I(N__15601));
    CascadeMux I__2299 (
            .O(N__15601),
            .I(N__15598));
    CascadeBuf I__2298 (
            .O(N__15598),
            .I(N__15595));
    CascadeMux I__2297 (
            .O(N__15595),
            .I(N__15592));
    CascadeBuf I__2296 (
            .O(N__15592),
            .I(N__15589));
    CascadeMux I__2295 (
            .O(N__15589),
            .I(N__15586));
    CascadeBuf I__2294 (
            .O(N__15586),
            .I(N__15583));
    CascadeMux I__2293 (
            .O(N__15583),
            .I(N__15580));
    CascadeBuf I__2292 (
            .O(N__15580),
            .I(N__15577));
    CascadeMux I__2291 (
            .O(N__15577),
            .I(N__15574));
    CascadeBuf I__2290 (
            .O(N__15574),
            .I(N__15571));
    CascadeMux I__2289 (
            .O(N__15571),
            .I(N__15568));
    CascadeBuf I__2288 (
            .O(N__15568),
            .I(N__15565));
    CascadeMux I__2287 (
            .O(N__15565),
            .I(N__15562));
    CascadeBuf I__2286 (
            .O(N__15562),
            .I(N__15559));
    CascadeMux I__2285 (
            .O(N__15559),
            .I(N__15556));
    CascadeBuf I__2284 (
            .O(N__15556),
            .I(N__15553));
    CascadeMux I__2283 (
            .O(N__15553),
            .I(N__15550));
    CascadeBuf I__2282 (
            .O(N__15550),
            .I(N__15547));
    CascadeMux I__2281 (
            .O(N__15547),
            .I(N__15544));
    CascadeBuf I__2280 (
            .O(N__15544),
            .I(N__15541));
    CascadeMux I__2279 (
            .O(N__15541),
            .I(N__15538));
    CascadeBuf I__2278 (
            .O(N__15538),
            .I(N__15535));
    CascadeMux I__2277 (
            .O(N__15535),
            .I(N__15532));
    CascadeBuf I__2276 (
            .O(N__15532),
            .I(N__15529));
    CascadeMux I__2275 (
            .O(N__15529),
            .I(N__15526));
    CascadeBuf I__2274 (
            .O(N__15526),
            .I(N__15523));
    CascadeMux I__2273 (
            .O(N__15523),
            .I(N__15520));
    InMux I__2272 (
            .O(N__15520),
            .I(N__15517));
    LocalMux I__2271 (
            .O(N__15517),
            .I(N__15514));
    Span4Mux_h I__2270 (
            .O(N__15514),
            .I(N__15509));
    InMux I__2269 (
            .O(N__15513),
            .I(N__15506));
    InMux I__2268 (
            .O(N__15512),
            .I(N__15502));
    Span4Mux_v I__2267 (
            .O(N__15509),
            .I(N__15499));
    LocalMux I__2266 (
            .O(N__15506),
            .I(N__15496));
    InMux I__2265 (
            .O(N__15505),
            .I(N__15493));
    LocalMux I__2264 (
            .O(N__15502),
            .I(N__15488));
    Span4Mux_v I__2263 (
            .O(N__15499),
            .I(N__15488));
    Odrv4 I__2262 (
            .O(N__15496),
            .I(M_this_ppu_sprites_addr_4));
    LocalMux I__2261 (
            .O(N__15493),
            .I(M_this_ppu_sprites_addr_4));
    Odrv4 I__2260 (
            .O(N__15488),
            .I(M_this_ppu_sprites_addr_4));
    InMux I__2259 (
            .O(N__15481),
            .I(N__15478));
    LocalMux I__2258 (
            .O(N__15478),
            .I(\this_vga_signals.g0_2_0_2_x1 ));
    CascadeMux I__2257 (
            .O(N__15475),
            .I(\this_vga_signals.g0_2_0_2_x0_cascade_ ));
    CascadeMux I__2256 (
            .O(N__15472),
            .I(\this_vga_signals.g0_2_0_2_cascade_ ));
    InMux I__2255 (
            .O(N__15469),
            .I(N__15466));
    LocalMux I__2254 (
            .O(N__15466),
            .I(N__15463));
    Span4Mux_v I__2253 (
            .O(N__15463),
            .I(N__15460));
    Sp12to4 I__2252 (
            .O(N__15460),
            .I(N__15457));
    Span12Mux_v I__2251 (
            .O(N__15457),
            .I(N__15454));
    Odrv12 I__2250 (
            .O(N__15454),
            .I(\this_sprites_ram.mem_out_bus7_2 ));
    InMux I__2249 (
            .O(N__15451),
            .I(N__15448));
    LocalMux I__2248 (
            .O(N__15448),
            .I(N__15445));
    Span4Mux_v I__2247 (
            .O(N__15445),
            .I(N__15442));
    Span4Mux_h I__2246 (
            .O(N__15442),
            .I(N__15439));
    Odrv4 I__2245 (
            .O(N__15439),
            .I(\this_sprites_ram.mem_out_bus3_2 ));
    InMux I__2244 (
            .O(N__15436),
            .I(N__15433));
    LocalMux I__2243 (
            .O(N__15433),
            .I(N__15430));
    Span4Mux_h I__2242 (
            .O(N__15430),
            .I(N__15427));
    Span4Mux_v I__2241 (
            .O(N__15427),
            .I(N__15424));
    Odrv4 I__2240 (
            .O(N__15424),
            .I(\this_sprites_ram.mem_out_bus5_0 ));
    InMux I__2239 (
            .O(N__15421),
            .I(N__15418));
    LocalMux I__2238 (
            .O(N__15418),
            .I(N__15415));
    Span4Mux_h I__2237 (
            .O(N__15415),
            .I(N__15412));
    Span4Mux_v I__2236 (
            .O(N__15412),
            .I(N__15409));
    Span4Mux_v I__2235 (
            .O(N__15409),
            .I(N__15406));
    Odrv4 I__2234 (
            .O(N__15406),
            .I(\this_sprites_ram.mem_out_bus1_0 ));
    CEMux I__2233 (
            .O(N__15403),
            .I(N__15399));
    CEMux I__2232 (
            .O(N__15402),
            .I(N__15396));
    LocalMux I__2231 (
            .O(N__15399),
            .I(N__15393));
    LocalMux I__2230 (
            .O(N__15396),
            .I(N__15390));
    Span4Mux_v I__2229 (
            .O(N__15393),
            .I(N__15387));
    Span4Mux_h I__2228 (
            .O(N__15390),
            .I(N__15384));
    Odrv4 I__2227 (
            .O(N__15387),
            .I(\this_sprites_ram.mem_WE_8 ));
    Odrv4 I__2226 (
            .O(N__15384),
            .I(\this_sprites_ram.mem_WE_8 ));
    InMux I__2225 (
            .O(N__15379),
            .I(N__15376));
    LocalMux I__2224 (
            .O(N__15376),
            .I(\this_vga_ramdac.m6 ));
    InMux I__2223 (
            .O(N__15373),
            .I(N__15370));
    LocalMux I__2222 (
            .O(N__15370),
            .I(N__15366));
    CascadeMux I__2221 (
            .O(N__15369),
            .I(N__15363));
    Span12Mux_s6_h I__2220 (
            .O(N__15366),
            .I(N__15360));
    InMux I__2219 (
            .O(N__15363),
            .I(N__15357));
    Odrv12 I__2218 (
            .O(N__15360),
            .I(\this_vga_ramdac.N_2871_reto ));
    LocalMux I__2217 (
            .O(N__15357),
            .I(\this_vga_ramdac.N_2871_reto ));
    CascadeMux I__2216 (
            .O(N__15352),
            .I(G_384_cascade_));
    InMux I__2215 (
            .O(N__15349),
            .I(N__15346));
    LocalMux I__2214 (
            .O(N__15346),
            .I(N__15343));
    Span4Mux_h I__2213 (
            .O(N__15343),
            .I(N__15340));
    Span4Mux_h I__2212 (
            .O(N__15340),
            .I(N__15336));
    InMux I__2211 (
            .O(N__15339),
            .I(N__15333));
    Odrv4 I__2210 (
            .O(N__15336),
            .I(\this_vga_ramdac.N_2872_reto ));
    LocalMux I__2209 (
            .O(N__15333),
            .I(\this_vga_ramdac.N_2872_reto ));
    CascadeMux I__2208 (
            .O(N__15328),
            .I(\this_vga_signals.if_N_5_cascade_ ));
    InMux I__2207 (
            .O(N__15325),
            .I(N__15319));
    InMux I__2206 (
            .O(N__15324),
            .I(N__15314));
    InMux I__2205 (
            .O(N__15323),
            .I(N__15314));
    InMux I__2204 (
            .O(N__15322),
            .I(N__15311));
    LocalMux I__2203 (
            .O(N__15319),
            .I(N__15305));
    LocalMux I__2202 (
            .O(N__15314),
            .I(N__15300));
    LocalMux I__2201 (
            .O(N__15311),
            .I(N__15300));
    InMux I__2200 (
            .O(N__15310),
            .I(N__15297));
    InMux I__2199 (
            .O(N__15309),
            .I(N__15292));
    InMux I__2198 (
            .O(N__15308),
            .I(N__15292));
    Span4Mux_h I__2197 (
            .O(N__15305),
            .I(N__15285));
    Span4Mux_v I__2196 (
            .O(N__15300),
            .I(N__15285));
    LocalMux I__2195 (
            .O(N__15297),
            .I(N__15280));
    LocalMux I__2194 (
            .O(N__15292),
            .I(N__15280));
    InMux I__2193 (
            .O(N__15291),
            .I(N__15275));
    InMux I__2192 (
            .O(N__15290),
            .I(N__15275));
    Odrv4 I__2191 (
            .O(N__15285),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__2190 (
            .O(N__15280),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__2189 (
            .O(N__15275),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    CascadeMux I__2188 (
            .O(N__15268),
            .I(\this_vga_signals.vaddress_5_cascade_ ));
    InMux I__2187 (
            .O(N__15265),
            .I(N__15261));
    InMux I__2186 (
            .O(N__15264),
            .I(N__15258));
    LocalMux I__2185 (
            .O(N__15261),
            .I(\this_vga_signals.g1_0_0_0 ));
    LocalMux I__2184 (
            .O(N__15258),
            .I(\this_vga_signals.g1_0_0_0 ));
    InMux I__2183 (
            .O(N__15253),
            .I(N__15250));
    LocalMux I__2182 (
            .O(N__15250),
            .I(\this_vga_signals.g0_1_2_0_1 ));
    CascadeMux I__2181 (
            .O(N__15247),
            .I(\this_vga_signals.g0_1_2_cascade_ ));
    InMux I__2180 (
            .O(N__15244),
            .I(N__15241));
    LocalMux I__2179 (
            .O(N__15241),
            .I(\this_vga_signals.g1_0_1_0_0 ));
    InMux I__2178 (
            .O(N__15238),
            .I(N__15235));
    LocalMux I__2177 (
            .O(N__15235),
            .I(N__15232));
    Odrv4 I__2176 (
            .O(N__15232),
            .I(\this_vga_signals.g2_0 ));
    InMux I__2175 (
            .O(N__15229),
            .I(N__15226));
    LocalMux I__2174 (
            .O(N__15226),
            .I(N__15223));
    Span4Mux_v I__2173 (
            .O(N__15223),
            .I(N__15220));
    Span4Mux_h I__2172 (
            .O(N__15220),
            .I(N__15217));
    Odrv4 I__2171 (
            .O(N__15217),
            .I(\this_vga_signals.g1_1_1 ));
    InMux I__2170 (
            .O(N__15214),
            .I(N__15211));
    LocalMux I__2169 (
            .O(N__15211),
            .I(\this_vga_signals.N_5_i_0 ));
    InMux I__2168 (
            .O(N__15208),
            .I(N__15205));
    LocalMux I__2167 (
            .O(N__15205),
            .I(\this_vga_signals.N_50 ));
    CascadeMux I__2166 (
            .O(N__15202),
            .I(\this_vga_signals.vaddress_1_6_cascade_ ));
    InMux I__2165 (
            .O(N__15199),
            .I(N__15196));
    LocalMux I__2164 (
            .O(N__15196),
            .I(N__15193));
    Span4Mux_v I__2163 (
            .O(N__15193),
            .I(N__15190));
    Odrv4 I__2162 (
            .O(N__15190),
            .I(\this_vga_signals.if_m8_0_a3_1_1_3 ));
    InMux I__2161 (
            .O(N__15187),
            .I(N__15184));
    LocalMux I__2160 (
            .O(N__15184),
            .I(N__15179));
    InMux I__2159 (
            .O(N__15183),
            .I(N__15174));
    InMux I__2158 (
            .O(N__15182),
            .I(N__15174));
    Span4Mux_v I__2157 (
            .O(N__15179),
            .I(N__15169));
    LocalMux I__2156 (
            .O(N__15174),
            .I(N__15169));
    Odrv4 I__2155 (
            .O(N__15169),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    InMux I__2154 (
            .O(N__15166),
            .I(N__15163));
    LocalMux I__2153 (
            .O(N__15163),
            .I(N__15160));
    Span4Mux_v I__2152 (
            .O(N__15160),
            .I(N__15155));
    InMux I__2151 (
            .O(N__15159),
            .I(N__15150));
    InMux I__2150 (
            .O(N__15158),
            .I(N__15150));
    Odrv4 I__2149 (
            .O(N__15155),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__2148 (
            .O(N__15150),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    CEMux I__2147 (
            .O(N__15145),
            .I(N__15121));
    CEMux I__2146 (
            .O(N__15144),
            .I(N__15121));
    CEMux I__2145 (
            .O(N__15143),
            .I(N__15121));
    CEMux I__2144 (
            .O(N__15142),
            .I(N__15121));
    CEMux I__2143 (
            .O(N__15141),
            .I(N__15121));
    CEMux I__2142 (
            .O(N__15140),
            .I(N__15121));
    CEMux I__2141 (
            .O(N__15139),
            .I(N__15121));
    CEMux I__2140 (
            .O(N__15138),
            .I(N__15121));
    GlobalMux I__2139 (
            .O(N__15121),
            .I(N__15118));
    gio2CtrlBuf I__2138 (
            .O(N__15118),
            .I(\this_vga_signals.N_614_1_g ));
    SRMux I__2137 (
            .O(N__15115),
            .I(N__15088));
    SRMux I__2136 (
            .O(N__15114),
            .I(N__15088));
    SRMux I__2135 (
            .O(N__15113),
            .I(N__15088));
    SRMux I__2134 (
            .O(N__15112),
            .I(N__15088));
    SRMux I__2133 (
            .O(N__15111),
            .I(N__15088));
    SRMux I__2132 (
            .O(N__15110),
            .I(N__15088));
    SRMux I__2131 (
            .O(N__15109),
            .I(N__15088));
    SRMux I__2130 (
            .O(N__15108),
            .I(N__15088));
    SRMux I__2129 (
            .O(N__15107),
            .I(N__15088));
    GlobalMux I__2128 (
            .O(N__15088),
            .I(N__15085));
    gio2CtrlBuf I__2127 (
            .O(N__15085),
            .I(\this_vga_signals.N_931_g ));
    CascadeMux I__2126 (
            .O(N__15082),
            .I(N__15078));
    InMux I__2125 (
            .O(N__15081),
            .I(N__15073));
    InMux I__2124 (
            .O(N__15078),
            .I(N__15067));
    InMux I__2123 (
            .O(N__15077),
            .I(N__15067));
    CascadeMux I__2122 (
            .O(N__15076),
            .I(N__15061));
    LocalMux I__2121 (
            .O(N__15073),
            .I(N__15057));
    InMux I__2120 (
            .O(N__15072),
            .I(N__15054));
    LocalMux I__2119 (
            .O(N__15067),
            .I(N__15051));
    InMux I__2118 (
            .O(N__15066),
            .I(N__15048));
    InMux I__2117 (
            .O(N__15065),
            .I(N__15045));
    InMux I__2116 (
            .O(N__15064),
            .I(N__15040));
    InMux I__2115 (
            .O(N__15061),
            .I(N__15040));
    CascadeMux I__2114 (
            .O(N__15060),
            .I(N__15036));
    Span4Mux_v I__2113 (
            .O(N__15057),
            .I(N__15031));
    LocalMux I__2112 (
            .O(N__15054),
            .I(N__15031));
    Span4Mux_v I__2111 (
            .O(N__15051),
            .I(N__15022));
    LocalMux I__2110 (
            .O(N__15048),
            .I(N__15022));
    LocalMux I__2109 (
            .O(N__15045),
            .I(N__15022));
    LocalMux I__2108 (
            .O(N__15040),
            .I(N__15022));
    InMux I__2107 (
            .O(N__15039),
            .I(N__15017));
    InMux I__2106 (
            .O(N__15036),
            .I(N__15017));
    Odrv4 I__2105 (
            .O(N__15031),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv4 I__2104 (
            .O(N__15022),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__2103 (
            .O(N__15017),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    CascadeMux I__2102 (
            .O(N__15010),
            .I(\this_vga_signals.if_m8_0_a3_1_1_1_cascade_ ));
    InMux I__2101 (
            .O(N__15007),
            .I(N__15004));
    LocalMux I__2100 (
            .O(N__15004),
            .I(\this_vga_signals.mult1_un40_sum_axb1_0 ));
    CascadeMux I__2099 (
            .O(N__15001),
            .I(\this_vga_signals.SUM_2_i_1_2_3_cascade_ ));
    InMux I__2098 (
            .O(N__14998),
            .I(N__14995));
    LocalMux I__2097 (
            .O(N__14995),
            .I(N__14988));
    InMux I__2096 (
            .O(N__14994),
            .I(N__14983));
    InMux I__2095 (
            .O(N__14993),
            .I(N__14983));
    InMux I__2094 (
            .O(N__14992),
            .I(N__14978));
    InMux I__2093 (
            .O(N__14991),
            .I(N__14978));
    Odrv4 I__2092 (
            .O(N__14988),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__2091 (
            .O(N__14983),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__2090 (
            .O(N__14978),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    CascadeMux I__2089 (
            .O(N__14971),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_ ));
    InMux I__2088 (
            .O(N__14968),
            .I(N__14962));
    InMux I__2087 (
            .O(N__14967),
            .I(N__14959));
    InMux I__2086 (
            .O(N__14966),
            .I(N__14954));
    InMux I__2085 (
            .O(N__14965),
            .I(N__14954));
    LocalMux I__2084 (
            .O(N__14962),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__2083 (
            .O(N__14959),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__2082 (
            .O(N__14954),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    InMux I__2081 (
            .O(N__14947),
            .I(N__14944));
    LocalMux I__2080 (
            .O(N__14944),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ));
    CascadeMux I__2079 (
            .O(N__14941),
            .I(N__14934));
    InMux I__2078 (
            .O(N__14940),
            .I(N__14931));
    InMux I__2077 (
            .O(N__14939),
            .I(N__14928));
    InMux I__2076 (
            .O(N__14938),
            .I(N__14923));
    InMux I__2075 (
            .O(N__14937),
            .I(N__14923));
    InMux I__2074 (
            .O(N__14934),
            .I(N__14920));
    LocalMux I__2073 (
            .O(N__14931),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__2072 (
            .O(N__14928),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__2071 (
            .O(N__14923),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__2070 (
            .O(N__14920),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    InMux I__2069 (
            .O(N__14911),
            .I(N__14904));
    InMux I__2068 (
            .O(N__14910),
            .I(N__14904));
    InMux I__2067 (
            .O(N__14909),
            .I(N__14901));
    LocalMux I__2066 (
            .O(N__14904),
            .I(N__14898));
    LocalMux I__2065 (
            .O(N__14901),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    Odrv4 I__2064 (
            .O(N__14898),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    CascadeMux I__2063 (
            .O(N__14893),
            .I(N__14887));
    InMux I__2062 (
            .O(N__14892),
            .I(N__14883));
    InMux I__2061 (
            .O(N__14891),
            .I(N__14880));
    InMux I__2060 (
            .O(N__14890),
            .I(N__14877));
    InMux I__2059 (
            .O(N__14887),
            .I(N__14872));
    InMux I__2058 (
            .O(N__14886),
            .I(N__14872));
    LocalMux I__2057 (
            .O(N__14883),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__2056 (
            .O(N__14880),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__2055 (
            .O(N__14877),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__2054 (
            .O(N__14872),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    InMux I__2053 (
            .O(N__14863),
            .I(N__14860));
    LocalMux I__2052 (
            .O(N__14860),
            .I(\this_vga_signals.SUM_2_i_1_0_3 ));
    CascadeMux I__2051 (
            .O(N__14857),
            .I(N__14854));
    InMux I__2050 (
            .O(N__14854),
            .I(N__14851));
    LocalMux I__2049 (
            .O(N__14851),
            .I(\this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5Z0Z_0 ));
    InMux I__2048 (
            .O(N__14848),
            .I(N__14845));
    LocalMux I__2047 (
            .O(N__14845),
            .I(\this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJHZ0Z5 ));
    CascadeMux I__2046 (
            .O(N__14842),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i_cascade_));
    InMux I__2045 (
            .O(N__14839),
            .I(N__14836));
    LocalMux I__2044 (
            .O(N__14836),
            .I(N__14830));
    InMux I__2043 (
            .O(N__14835),
            .I(N__14825));
    InMux I__2042 (
            .O(N__14834),
            .I(N__14825));
    InMux I__2041 (
            .O(N__14833),
            .I(N__14822));
    Span4Mux_v I__2040 (
            .O(N__14830),
            .I(N__14817));
    LocalMux I__2039 (
            .O(N__14825),
            .I(N__14817));
    LocalMux I__2038 (
            .O(N__14822),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    Odrv4 I__2037 (
            .O(N__14817),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    InMux I__2036 (
            .O(N__14812),
            .I(N__14809));
    LocalMux I__2035 (
            .O(N__14809),
            .I(N__14806));
    Span4Mux_v I__2034 (
            .O(N__14806),
            .I(N__14801));
    InMux I__2033 (
            .O(N__14805),
            .I(N__14798));
    InMux I__2032 (
            .O(N__14804),
            .I(N__14795));
    Odrv4 I__2031 (
            .O(N__14801),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    LocalMux I__2030 (
            .O(N__14798),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    LocalMux I__2029 (
            .O(N__14795),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    InMux I__2028 (
            .O(N__14788),
            .I(N__14782));
    InMux I__2027 (
            .O(N__14787),
            .I(N__14782));
    LocalMux I__2026 (
            .O(N__14782),
            .I(N__14779));
    Span4Mux_h I__2025 (
            .O(N__14779),
            .I(N__14775));
    InMux I__2024 (
            .O(N__14778),
            .I(N__14772));
    Odrv4 I__2023 (
            .O(N__14775),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    LocalMux I__2022 (
            .O(N__14772),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    CascadeMux I__2021 (
            .O(N__14767),
            .I(N__14764));
    InMux I__2020 (
            .O(N__14764),
            .I(N__14761));
    LocalMux I__2019 (
            .O(N__14761),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    CascadeMux I__2018 (
            .O(N__14758),
            .I(N__14755));
    InMux I__2017 (
            .O(N__14755),
            .I(N__14752));
    LocalMux I__2016 (
            .O(N__14752),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1 ));
    InMux I__2015 (
            .O(N__14749),
            .I(N__14746));
    LocalMux I__2014 (
            .O(N__14746),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    CascadeMux I__2013 (
            .O(N__14743),
            .I(\this_vga_signals.N_1_4_1_cascade_ ));
    CascadeMux I__2012 (
            .O(N__14740),
            .I(N_2_0_cascade_));
    InMux I__2011 (
            .O(N__14737),
            .I(N__14732));
    InMux I__2010 (
            .O(N__14736),
            .I(N__14729));
    InMux I__2009 (
            .O(N__14735),
            .I(N__14726));
    LocalMux I__2008 (
            .O(N__14732),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__2007 (
            .O(N__14729),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__2006 (
            .O(N__14726),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    CascadeMux I__2005 (
            .O(N__14719),
            .I(N__14711));
    CascadeMux I__2004 (
            .O(N__14718),
            .I(N__14707));
    CEMux I__2003 (
            .O(N__14717),
            .I(N__14703));
    InMux I__2002 (
            .O(N__14716),
            .I(N__14700));
    InMux I__2001 (
            .O(N__14715),
            .I(N__14695));
    InMux I__2000 (
            .O(N__14714),
            .I(N__14695));
    InMux I__1999 (
            .O(N__14711),
            .I(N__14684));
    InMux I__1998 (
            .O(N__14710),
            .I(N__14684));
    InMux I__1997 (
            .O(N__14707),
            .I(N__14679));
    InMux I__1996 (
            .O(N__14706),
            .I(N__14679));
    LocalMux I__1995 (
            .O(N__14703),
            .I(N__14676));
    LocalMux I__1994 (
            .O(N__14700),
            .I(N__14673));
    LocalMux I__1993 (
            .O(N__14695),
            .I(N__14670));
    InMux I__1992 (
            .O(N__14694),
            .I(N__14665));
    InMux I__1991 (
            .O(N__14693),
            .I(N__14665));
    InMux I__1990 (
            .O(N__14692),
            .I(N__14659));
    InMux I__1989 (
            .O(N__14691),
            .I(N__14659));
    InMux I__1988 (
            .O(N__14690),
            .I(N__14654));
    InMux I__1987 (
            .O(N__14689),
            .I(N__14654));
    LocalMux I__1986 (
            .O(N__14684),
            .I(N__14651));
    LocalMux I__1985 (
            .O(N__14679),
            .I(N__14645));
    Span4Mux_h I__1984 (
            .O(N__14676),
            .I(N__14645));
    Span4Mux_h I__1983 (
            .O(N__14673),
            .I(N__14642));
    Sp12to4 I__1982 (
            .O(N__14670),
            .I(N__14637));
    LocalMux I__1981 (
            .O(N__14665),
            .I(N__14637));
    InMux I__1980 (
            .O(N__14664),
            .I(N__14633));
    LocalMux I__1979 (
            .O(N__14659),
            .I(N__14626));
    LocalMux I__1978 (
            .O(N__14654),
            .I(N__14626));
    Span4Mux_h I__1977 (
            .O(N__14651),
            .I(N__14626));
    InMux I__1976 (
            .O(N__14650),
            .I(N__14623));
    Span4Mux_h I__1975 (
            .O(N__14645),
            .I(N__14620));
    Span4Mux_h I__1974 (
            .O(N__14642),
            .I(N__14617));
    Span12Mux_h I__1973 (
            .O(N__14637),
            .I(N__14614));
    InMux I__1972 (
            .O(N__14636),
            .I(N__14611));
    LocalMux I__1971 (
            .O(N__14633),
            .I(N__14604));
    Span4Mux_h I__1970 (
            .O(N__14626),
            .I(N__14604));
    LocalMux I__1969 (
            .O(N__14623),
            .I(N__14604));
    Odrv4 I__1968 (
            .O(N__14620),
            .I(M_counter_q_RNILQS8_1));
    Odrv4 I__1967 (
            .O(N__14617),
            .I(M_counter_q_RNILQS8_1));
    Odrv12 I__1966 (
            .O(N__14614),
            .I(M_counter_q_RNILQS8_1));
    LocalMux I__1965 (
            .O(N__14611),
            .I(M_counter_q_RNILQS8_1));
    Odrv4 I__1964 (
            .O(N__14604),
            .I(M_counter_q_RNILQS8_1));
    CascadeMux I__1963 (
            .O(N__14593),
            .I(\this_vga_signals.M_pcounter_q_3_1_cascade_ ));
    CascadeMux I__1962 (
            .O(N__14590),
            .I(N__14586));
    CascadeMux I__1961 (
            .O(N__14589),
            .I(N__14582));
    InMux I__1960 (
            .O(N__14586),
            .I(N__14579));
    InMux I__1959 (
            .O(N__14585),
            .I(N__14574));
    InMux I__1958 (
            .O(N__14582),
            .I(N__14574));
    LocalMux I__1957 (
            .O(N__14579),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    LocalMux I__1956 (
            .O(N__14574),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    CascadeMux I__1955 (
            .O(N__14569),
            .I(N_3_0_cascade_));
    InMux I__1954 (
            .O(N__14566),
            .I(N__14558));
    InMux I__1953 (
            .O(N__14565),
            .I(N__14558));
    InMux I__1952 (
            .O(N__14564),
            .I(N__14553));
    InMux I__1951 (
            .O(N__14563),
            .I(N__14553));
    LocalMux I__1950 (
            .O(N__14558),
            .I(\this_vga_signals.M_pcounter_q_i_5_1 ));
    LocalMux I__1949 (
            .O(N__14553),
            .I(\this_vga_signals.M_pcounter_q_i_5_1 ));
    InMux I__1948 (
            .O(N__14548),
            .I(N__14544));
    InMux I__1947 (
            .O(N__14547),
            .I(N__14541));
    LocalMux I__1946 (
            .O(N__14544),
            .I(\this_vga_signals.M_pcounter_q_i_5_0 ));
    LocalMux I__1945 (
            .O(N__14541),
            .I(\this_vga_signals.M_pcounter_q_i_5_0 ));
    CascadeMux I__1944 (
            .O(N__14536),
            .I(N__14532));
    InMux I__1943 (
            .O(N__14535),
            .I(N__14525));
    InMux I__1942 (
            .O(N__14532),
            .I(N__14522));
    InMux I__1941 (
            .O(N__14531),
            .I(N__14519));
    InMux I__1940 (
            .O(N__14530),
            .I(N__14512));
    InMux I__1939 (
            .O(N__14529),
            .I(N__14512));
    InMux I__1938 (
            .O(N__14528),
            .I(N__14512));
    LocalMux I__1937 (
            .O(N__14525),
            .I(N__14509));
    LocalMux I__1936 (
            .O(N__14522),
            .I(N__14506));
    LocalMux I__1935 (
            .O(N__14519),
            .I(N__14501));
    LocalMux I__1934 (
            .O(N__14512),
            .I(N__14498));
    Span4Mux_h I__1933 (
            .O(N__14509),
            .I(N__14493));
    Span4Mux_h I__1932 (
            .O(N__14506),
            .I(N__14493));
    InMux I__1931 (
            .O(N__14505),
            .I(N__14488));
    InMux I__1930 (
            .O(N__14504),
            .I(N__14488));
    Span4Mux_h I__1929 (
            .O(N__14501),
            .I(N__14485));
    Span4Mux_h I__1928 (
            .O(N__14498),
            .I(N__14482));
    Span4Mux_v I__1927 (
            .O(N__14493),
            .I(N__14479));
    LocalMux I__1926 (
            .O(N__14488),
            .I(N__14476));
    Span4Mux_h I__1925 (
            .O(N__14485),
            .I(N__14472));
    Span4Mux_h I__1924 (
            .O(N__14482),
            .I(N__14469));
    Span4Mux_v I__1923 (
            .O(N__14479),
            .I(N__14464));
    Span4Mux_h I__1922 (
            .O(N__14476),
            .I(N__14464));
    InMux I__1921 (
            .O(N__14475),
            .I(N__14461));
    Odrv4 I__1920 (
            .O(N__14472),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__1919 (
            .O(N__14469),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__1918 (
            .O(N__14464),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    LocalMux I__1917 (
            .O(N__14461),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    InMux I__1916 (
            .O(N__14452),
            .I(N__14449));
    LocalMux I__1915 (
            .O(N__14449),
            .I(\this_vga_signals.M_pcounter_q_3_0 ));
    CEMux I__1914 (
            .O(N__14446),
            .I(N__14442));
    CEMux I__1913 (
            .O(N__14445),
            .I(N__14439));
    LocalMux I__1912 (
            .O(N__14442),
            .I(N__14436));
    LocalMux I__1911 (
            .O(N__14439),
            .I(N__14433));
    Span4Mux_v I__1910 (
            .O(N__14436),
            .I(N__14430));
    Span4Mux_h I__1909 (
            .O(N__14433),
            .I(N__14427));
    Odrv4 I__1908 (
            .O(N__14430),
            .I(\this_sprites_ram.mem_WE_4 ));
    Odrv4 I__1907 (
            .O(N__14427),
            .I(\this_sprites_ram.mem_WE_4 ));
    InMux I__1906 (
            .O(N__14422),
            .I(N__14419));
    LocalMux I__1905 (
            .O(N__14419),
            .I(N__14416));
    Span4Mux_v I__1904 (
            .O(N__14416),
            .I(N__14412));
    InMux I__1903 (
            .O(N__14415),
            .I(N__14409));
    Odrv4 I__1902 (
            .O(N__14412),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    LocalMux I__1901 (
            .O(N__14409),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    InMux I__1900 (
            .O(N__14404),
            .I(N__14401));
    LocalMux I__1899 (
            .O(N__14401),
            .I(N__14397));
    CascadeMux I__1898 (
            .O(N__14400),
            .I(N__14393));
    Span4Mux_h I__1897 (
            .O(N__14397),
            .I(N__14389));
    InMux I__1896 (
            .O(N__14396),
            .I(N__14386));
    InMux I__1895 (
            .O(N__14393),
            .I(N__14381));
    InMux I__1894 (
            .O(N__14392),
            .I(N__14381));
    Odrv4 I__1893 (
            .O(N__14389),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__1892 (
            .O(N__14386),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__1891 (
            .O(N__14381),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    InMux I__1890 (
            .O(N__14374),
            .I(N__14371));
    LocalMux I__1889 (
            .O(N__14371),
            .I(N__14368));
    Span4Mux_v I__1888 (
            .O(N__14368),
            .I(N__14363));
    InMux I__1887 (
            .O(N__14367),
            .I(N__14358));
    InMux I__1886 (
            .O(N__14366),
            .I(N__14358));
    Odrv4 I__1885 (
            .O(N__14363),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_2 ));
    LocalMux I__1884 (
            .O(N__14358),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_2 ));
    CascadeMux I__1883 (
            .O(N__14353),
            .I(N__14350));
    InMux I__1882 (
            .O(N__14350),
            .I(N__14347));
    LocalMux I__1881 (
            .O(N__14347),
            .I(N__14344));
    Span12Mux_h I__1880 (
            .O(N__14344),
            .I(N__14341));
    Odrv12 I__1879 (
            .O(N__14341),
            .I(M_this_vga_signals_address_3));
    CEMux I__1878 (
            .O(N__14338),
            .I(N__14335));
    LocalMux I__1877 (
            .O(N__14335),
            .I(N__14331));
    CEMux I__1876 (
            .O(N__14334),
            .I(N__14328));
    Span4Mux_h I__1875 (
            .O(N__14331),
            .I(N__14325));
    LocalMux I__1874 (
            .O(N__14328),
            .I(N__14322));
    Span4Mux_h I__1873 (
            .O(N__14325),
            .I(N__14319));
    Span4Mux_h I__1872 (
            .O(N__14322),
            .I(N__14316));
    Odrv4 I__1871 (
            .O(N__14319),
            .I(\this_sprites_ram.mem_WE_6 ));
    Odrv4 I__1870 (
            .O(N__14316),
            .I(\this_sprites_ram.mem_WE_6 ));
    InMux I__1869 (
            .O(N__14311),
            .I(N__14308));
    LocalMux I__1868 (
            .O(N__14308),
            .I(N__14305));
    Span4Mux_v I__1867 (
            .O(N__14305),
            .I(N__14298));
    InMux I__1866 (
            .O(N__14304),
            .I(N__14295));
    InMux I__1865 (
            .O(N__14303),
            .I(N__14290));
    InMux I__1864 (
            .O(N__14302),
            .I(N__14290));
    InMux I__1863 (
            .O(N__14301),
            .I(N__14287));
    Odrv4 I__1862 (
            .O(N__14298),
            .I(\this_vga_signals.N_3_2_1 ));
    LocalMux I__1861 (
            .O(N__14295),
            .I(\this_vga_signals.N_3_2_1 ));
    LocalMux I__1860 (
            .O(N__14290),
            .I(\this_vga_signals.N_3_2_1 ));
    LocalMux I__1859 (
            .O(N__14287),
            .I(\this_vga_signals.N_3_2_1 ));
    CascadeMux I__1858 (
            .O(N__14278),
            .I(N__14275));
    InMux I__1857 (
            .O(N__14275),
            .I(N__14272));
    LocalMux I__1856 (
            .O(N__14272),
            .I(N__14269));
    Span12Mux_h I__1855 (
            .O(N__14269),
            .I(N__14266));
    Odrv12 I__1854 (
            .O(N__14266),
            .I(M_this_vga_signals_address_6));
    CascadeMux I__1853 (
            .O(N__14263),
            .I(N__14260));
    InMux I__1852 (
            .O(N__14260),
            .I(N__14256));
    InMux I__1851 (
            .O(N__14259),
            .I(N__14253));
    LocalMux I__1850 (
            .O(N__14256),
            .I(N__14250));
    LocalMux I__1849 (
            .O(N__14253),
            .I(N__14247));
    Span4Mux_v I__1848 (
            .O(N__14250),
            .I(N__14242));
    Span4Mux_v I__1847 (
            .O(N__14247),
            .I(N__14242));
    Odrv4 I__1846 (
            .O(N__14242),
            .I(\this_vga_signals.M_vcounter_d7lto8_1 ));
    CascadeMux I__1845 (
            .O(N__14239),
            .I(N__14236));
    InMux I__1844 (
            .O(N__14236),
            .I(N__14233));
    LocalMux I__1843 (
            .O(N__14233),
            .I(\this_vga_signals.M_lcounter_d_0_sqmuxa ));
    CascadeMux I__1842 (
            .O(N__14230),
            .I(\this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_ ));
    InMux I__1841 (
            .O(N__14227),
            .I(N__14224));
    LocalMux I__1840 (
            .O(N__14224),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_1_0 ));
    CascadeMux I__1839 (
            .O(N__14221),
            .I(\this_vga_signals.g1_0_0_1_cascade_ ));
    CascadeMux I__1838 (
            .O(N__14218),
            .I(\this_vga_signals.g2_0_1_cascade_ ));
    InMux I__1837 (
            .O(N__14215),
            .I(N__14212));
    LocalMux I__1836 (
            .O(N__14212),
            .I(\this_vga_signals.vaddress_6_6 ));
    InMux I__1835 (
            .O(N__14209),
            .I(N__14206));
    LocalMux I__1834 (
            .O(N__14206),
            .I(\this_vga_signals.N_4_1_0 ));
    CascadeMux I__1833 (
            .O(N__14203),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_ ));
    InMux I__1832 (
            .O(N__14200),
            .I(N__14197));
    LocalMux I__1831 (
            .O(N__14197),
            .I(\this_vga_signals.g0_i_x4_0_0 ));
    CascadeMux I__1830 (
            .O(N__14194),
            .I(\this_vga_signals.g1_4_cascade_ ));
    InMux I__1829 (
            .O(N__14191),
            .I(N__14188));
    LocalMux I__1828 (
            .O(N__14188),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_1_0_0_1 ));
    CascadeMux I__1827 (
            .O(N__14185),
            .I(\this_vga_signals.g0_2_0_0_1_cascade_ ));
    InMux I__1826 (
            .O(N__14182),
            .I(N__14179));
    LocalMux I__1825 (
            .O(N__14179),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_0_0_0 ));
    CascadeMux I__1824 (
            .O(N__14176),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ));
    InMux I__1823 (
            .O(N__14173),
            .I(N__14170));
    LocalMux I__1822 (
            .O(N__14170),
            .I(N__14167));
    Odrv4 I__1821 (
            .O(N__14167),
            .I(\this_vga_signals.g1_0_1 ));
    InMux I__1820 (
            .O(N__14164),
            .I(N__14161));
    LocalMux I__1819 (
            .O(N__14161),
            .I(\this_vga_signals.g0_31_N_5L8 ));
    CascadeMux I__1818 (
            .O(N__14158),
            .I(N__14155));
    InMux I__1817 (
            .O(N__14155),
            .I(N__14152));
    LocalMux I__1816 (
            .O(N__14152),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_0 ));
    CascadeMux I__1815 (
            .O(N__14149),
            .I(\this_vga_signals.m9_1_cascade_ ));
    InMux I__1814 (
            .O(N__14146),
            .I(N__14143));
    LocalMux I__1813 (
            .O(N__14143),
            .I(\this_vga_signals.g2_1_0 ));
    InMux I__1812 (
            .O(N__14140),
            .I(N__14137));
    LocalMux I__1811 (
            .O(N__14137),
            .I(N__14133));
    InMux I__1810 (
            .O(N__14136),
            .I(N__14130));
    Span4Mux_h I__1809 (
            .O(N__14133),
            .I(N__14125));
    LocalMux I__1808 (
            .O(N__14130),
            .I(N__14125));
    Odrv4 I__1807 (
            .O(N__14125),
            .I(\this_vga_signals.vaddress_c2 ));
    CascadeMux I__1806 (
            .O(N__14122),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_ ));
    InMux I__1805 (
            .O(N__14119),
            .I(N__14116));
    LocalMux I__1804 (
            .O(N__14116),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    InMux I__1803 (
            .O(N__14113),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__1802 (
            .O(N__14110),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__1801 (
            .O(N__14107),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__1800 (
            .O(N__14104),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__1799 (
            .O(N__14101),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__1798 (
            .O(N__14098),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__1797 (
            .O(N__14095),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__1796 (
            .O(N__14092),
            .I(bfn_10_12_0_));
    InMux I__1795 (
            .O(N__14089),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    InMux I__1794 (
            .O(N__14086),
            .I(N__14083));
    LocalMux I__1793 (
            .O(N__14083),
            .I(N__14080));
    Odrv4 I__1792 (
            .O(N__14080),
            .I(\this_sprites_ram.mem_out_bus4_3 ));
    InMux I__1791 (
            .O(N__14077),
            .I(N__14074));
    LocalMux I__1790 (
            .O(N__14074),
            .I(N__14071));
    Span4Mux_v I__1789 (
            .O(N__14071),
            .I(N__14068));
    Span4Mux_v I__1788 (
            .O(N__14068),
            .I(N__14065));
    Span4Mux_v I__1787 (
            .O(N__14065),
            .I(N__14062));
    Odrv4 I__1786 (
            .O(N__14062),
            .I(\this_sprites_ram.mem_out_bus0_3 ));
    CascadeMux I__1785 (
            .O(N__14059),
            .I(N__14056));
    InMux I__1784 (
            .O(N__14056),
            .I(N__14053));
    LocalMux I__1783 (
            .O(N__14053),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ));
    InMux I__1782 (
            .O(N__14050),
            .I(N__14047));
    LocalMux I__1781 (
            .O(N__14047),
            .I(N__14044));
    Span4Mux_v I__1780 (
            .O(N__14044),
            .I(N__14041));
    Odrv4 I__1779 (
            .O(N__14041),
            .I(\this_sprites_ram.mem_out_bus5_3 ));
    InMux I__1778 (
            .O(N__14038),
            .I(N__14035));
    LocalMux I__1777 (
            .O(N__14035),
            .I(N__14032));
    Span4Mux_v I__1776 (
            .O(N__14032),
            .I(N__14029));
    Span4Mux_v I__1775 (
            .O(N__14029),
            .I(N__14026));
    Odrv4 I__1774 (
            .O(N__14026),
            .I(\this_sprites_ram.mem_out_bus1_3 ));
    InMux I__1773 (
            .O(N__14023),
            .I(N__14020));
    LocalMux I__1772 (
            .O(N__14020),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ));
    InMux I__1771 (
            .O(N__14017),
            .I(N__14014));
    LocalMux I__1770 (
            .O(N__14014),
            .I(N__14007));
    InMux I__1769 (
            .O(N__14013),
            .I(N__14004));
    InMux I__1768 (
            .O(N__14012),
            .I(N__14001));
    InMux I__1767 (
            .O(N__14011),
            .I(N__13998));
    InMux I__1766 (
            .O(N__14010),
            .I(N__13995));
    Span4Mux_h I__1765 (
            .O(N__14007),
            .I(N__13990));
    LocalMux I__1764 (
            .O(N__14004),
            .I(N__13985));
    LocalMux I__1763 (
            .O(N__14001),
            .I(N__13985));
    LocalMux I__1762 (
            .O(N__13998),
            .I(N__13980));
    LocalMux I__1761 (
            .O(N__13995),
            .I(N__13980));
    InMux I__1760 (
            .O(N__13994),
            .I(N__13977));
    InMux I__1759 (
            .O(N__13993),
            .I(N__13974));
    Odrv4 I__1758 (
            .O(N__13990),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    Odrv4 I__1757 (
            .O(N__13985),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    Odrv4 I__1756 (
            .O(N__13980),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1755 (
            .O(N__13977),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1754 (
            .O(N__13974),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    CascadeMux I__1753 (
            .O(N__13963),
            .I(N__13960));
    InMux I__1752 (
            .O(N__13960),
            .I(N__13957));
    LocalMux I__1751 (
            .O(N__13957),
            .I(N__13954));
    Span12Mux_h I__1750 (
            .O(N__13954),
            .I(N__13951));
    Odrv12 I__1749 (
            .O(N__13951),
            .I(M_this_vga_signals_address_4));
    InMux I__1748 (
            .O(N__13948),
            .I(N__13945));
    LocalMux I__1747 (
            .O(N__13945),
            .I(N__13942));
    Span4Mux_v I__1746 (
            .O(N__13942),
            .I(N__13939));
    Span4Mux_v I__1745 (
            .O(N__13939),
            .I(N__13936));
    Span4Mux_v I__1744 (
            .O(N__13936),
            .I(N__13933));
    Odrv4 I__1743 (
            .O(N__13933),
            .I(\this_sprites_ram.mem_out_bus7_0 ));
    InMux I__1742 (
            .O(N__13930),
            .I(N__13927));
    LocalMux I__1741 (
            .O(N__13927),
            .I(N__13924));
    Span4Mux_h I__1740 (
            .O(N__13924),
            .I(N__13921));
    Odrv4 I__1739 (
            .O(N__13921),
            .I(\this_sprites_ram.mem_out_bus3_0 ));
    InMux I__1738 (
            .O(N__13918),
            .I(N__13915));
    LocalMux I__1737 (
            .O(N__13915),
            .I(N__13910));
    InMux I__1736 (
            .O(N__13914),
            .I(N__13905));
    InMux I__1735 (
            .O(N__13913),
            .I(N__13905));
    Odrv4 I__1734 (
            .O(N__13910),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__1733 (
            .O(N__13905),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    CascadeMux I__1732 (
            .O(N__13900),
            .I(N__13897));
    InMux I__1731 (
            .O(N__13897),
            .I(N__13894));
    LocalMux I__1730 (
            .O(N__13894),
            .I(N__13891));
    Span12Mux_h I__1729 (
            .O(N__13891),
            .I(N__13888));
    Odrv12 I__1728 (
            .O(N__13888),
            .I(M_this_vga_signals_address_2));
    InMux I__1727 (
            .O(N__13885),
            .I(N__13882));
    LocalMux I__1726 (
            .O(N__13882),
            .I(N__13879));
    Span4Mux_h I__1725 (
            .O(N__13879),
            .I(N__13876));
    Odrv4 I__1724 (
            .O(N__13876),
            .I(\this_vga_ramdac.m19 ));
    InMux I__1723 (
            .O(N__13873),
            .I(N__13870));
    LocalMux I__1722 (
            .O(N__13870),
            .I(N__13867));
    Span4Mux_v I__1721 (
            .O(N__13867),
            .I(N__13863));
    CascadeMux I__1720 (
            .O(N__13866),
            .I(N__13860));
    Span4Mux_h I__1719 (
            .O(N__13863),
            .I(N__13857));
    InMux I__1718 (
            .O(N__13860),
            .I(N__13854));
    Odrv4 I__1717 (
            .O(N__13857),
            .I(\this_vga_ramdac.N_2874_reto ));
    LocalMux I__1716 (
            .O(N__13854),
            .I(\this_vga_ramdac.N_2874_reto ));
    InMux I__1715 (
            .O(N__13849),
            .I(N__13841));
    InMux I__1714 (
            .O(N__13848),
            .I(N__13841));
    InMux I__1713 (
            .O(N__13847),
            .I(N__13838));
    InMux I__1712 (
            .O(N__13846),
            .I(N__13835));
    LocalMux I__1711 (
            .O(N__13841),
            .I(N__13831));
    LocalMux I__1710 (
            .O(N__13838),
            .I(N__13826));
    LocalMux I__1709 (
            .O(N__13835),
            .I(N__13826));
    InMux I__1708 (
            .O(N__13834),
            .I(N__13822));
    Span4Mux_v I__1707 (
            .O(N__13831),
            .I(N__13817));
    Span4Mux_v I__1706 (
            .O(N__13826),
            .I(N__13817));
    InMux I__1705 (
            .O(N__13825),
            .I(N__13814));
    LocalMux I__1704 (
            .O(N__13822),
            .I(N__13806));
    Sp12to4 I__1703 (
            .O(N__13817),
            .I(N__13806));
    LocalMux I__1702 (
            .O(N__13814),
            .I(N__13806));
    InMux I__1701 (
            .O(N__13813),
            .I(N__13803));
    Odrv12 I__1700 (
            .O(N__13806),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    LocalMux I__1699 (
            .O(N__13803),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    InMux I__1698 (
            .O(N__13798),
            .I(N__13795));
    LocalMux I__1697 (
            .O(N__13795),
            .I(N__13792));
    Span4Mux_v I__1696 (
            .O(N__13792),
            .I(N__13789));
    Span4Mux_v I__1695 (
            .O(N__13789),
            .I(N__13786));
    Span4Mux_v I__1694 (
            .O(N__13786),
            .I(N__13783));
    Odrv4 I__1693 (
            .O(N__13783),
            .I(\this_sprites_ram.mem_out_bus7_3 ));
    InMux I__1692 (
            .O(N__13780),
            .I(N__13777));
    LocalMux I__1691 (
            .O(N__13777),
            .I(N__13774));
    Odrv4 I__1690 (
            .O(N__13774),
            .I(\this_sprites_ram.mem_out_bus3_3 ));
    InMux I__1689 (
            .O(N__13771),
            .I(N__13768));
    LocalMux I__1688 (
            .O(N__13768),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ));
    InMux I__1687 (
            .O(N__13765),
            .I(N__13762));
    LocalMux I__1686 (
            .O(N__13762),
            .I(N__13758));
    InMux I__1685 (
            .O(N__13761),
            .I(N__13755));
    Odrv4 I__1684 (
            .O(N__13758),
            .I(\this_vga_signals.vaddress_6_5 ));
    LocalMux I__1683 (
            .O(N__13755),
            .I(\this_vga_signals.vaddress_6_5 ));
    InMux I__1682 (
            .O(N__13750),
            .I(N__13747));
    LocalMux I__1681 (
            .O(N__13747),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_1_0_0 ));
    CascadeMux I__1680 (
            .O(N__13744),
            .I(N__13740));
    InMux I__1679 (
            .O(N__13743),
            .I(N__13735));
    InMux I__1678 (
            .O(N__13740),
            .I(N__13735));
    LocalMux I__1677 (
            .O(N__13735),
            .I(N__13732));
    Odrv4 I__1676 (
            .O(N__13732),
            .I(\this_vga_signals.vaddress_3_0_6 ));
    CascadeMux I__1675 (
            .O(N__13729),
            .I(\this_vga_signals.vaddress_3_5_cascade_ ));
    CascadeMux I__1674 (
            .O(N__13726),
            .I(\this_vga_signals.vaddress_3_6_cascade_ ));
    CascadeMux I__1673 (
            .O(N__13723),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ));
    InMux I__1672 (
            .O(N__13720),
            .I(N__13717));
    LocalMux I__1671 (
            .O(N__13717),
            .I(N__13714));
    Span4Mux_v I__1670 (
            .O(N__13714),
            .I(N__13711));
    Sp12to4 I__1669 (
            .O(N__13711),
            .I(N__13708));
    Span12Mux_h I__1668 (
            .O(N__13708),
            .I(N__13705));
    Odrv12 I__1667 (
            .O(N__13705),
            .I(M_this_ppu_vram_data_3));
    InMux I__1666 (
            .O(N__13702),
            .I(N__13699));
    LocalMux I__1665 (
            .O(N__13699),
            .I(N__13696));
    Span4Mux_v I__1664 (
            .O(N__13696),
            .I(N__13693));
    Span4Mux_v I__1663 (
            .O(N__13693),
            .I(N__13690));
    Odrv4 I__1662 (
            .O(N__13690),
            .I(\this_sprites_ram.mem_out_bus6_3 ));
    InMux I__1661 (
            .O(N__13687),
            .I(N__13684));
    LocalMux I__1660 (
            .O(N__13684),
            .I(N__13681));
    Span4Mux_v I__1659 (
            .O(N__13681),
            .I(N__13678));
    Odrv4 I__1658 (
            .O(N__13678),
            .I(\this_sprites_ram.mem_out_bus2_3 ));
    InMux I__1657 (
            .O(N__13675),
            .I(N__13672));
    LocalMux I__1656 (
            .O(N__13672),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ));
    CascadeMux I__1655 (
            .O(N__13669),
            .I(\this_vga_signals.vaddress_3_0_6_cascade_ ));
    CascadeMux I__1654 (
            .O(N__13666),
            .I(\this_vga_signals.g2_3_cascade_ ));
    CascadeMux I__1653 (
            .O(N__13663),
            .I(\this_vga_signals.g1_1_1_cascade_ ));
    CascadeMux I__1652 (
            .O(N__13660),
            .I(\this_vga_signals.g0_i_x4_0_2_cascade_ ));
    InMux I__1651 (
            .O(N__13657),
            .I(N__13654));
    LocalMux I__1650 (
            .O(N__13654),
            .I(\this_vga_signals.g0_31_N_4L6 ));
    CascadeMux I__1649 (
            .O(N__13651),
            .I(\this_vga_signals.if_m8_0_a3_1_1_4_cascade_ ));
    InMux I__1648 (
            .O(N__13648),
            .I(N__13645));
    LocalMux I__1647 (
            .O(N__13645),
            .I(\this_vga_signals.g0_31_N_3L3 ));
    InMux I__1646 (
            .O(N__13642),
            .I(N__13639));
    LocalMux I__1645 (
            .O(N__13639),
            .I(\this_vga_signals.g3_3_0 ));
    CascadeMux I__1644 (
            .O(N__13636),
            .I(\this_vga_signals.if_m8_0_a3_1_1_2_cascade_ ));
    CascadeMux I__1643 (
            .O(N__13633),
            .I(\this_vga_signals.g0_8_0_cascade_ ));
    CascadeMux I__1642 (
            .O(N__13630),
            .I(\this_vga_signals.vaddress_2_5_cascade_ ));
    InMux I__1641 (
            .O(N__13627),
            .I(N__13622));
    CascadeMux I__1640 (
            .O(N__13626),
            .I(N__13619));
    CascadeMux I__1639 (
            .O(N__13625),
            .I(N__13615));
    LocalMux I__1638 (
            .O(N__13622),
            .I(N__13609));
    InMux I__1637 (
            .O(N__13619),
            .I(N__13605));
    InMux I__1636 (
            .O(N__13618),
            .I(N__13600));
    InMux I__1635 (
            .O(N__13615),
            .I(N__13600));
    InMux I__1634 (
            .O(N__13614),
            .I(N__13595));
    InMux I__1633 (
            .O(N__13613),
            .I(N__13595));
    InMux I__1632 (
            .O(N__13612),
            .I(N__13592));
    Span4Mux_v I__1631 (
            .O(N__13609),
            .I(N__13589));
    InMux I__1630 (
            .O(N__13608),
            .I(N__13586));
    LocalMux I__1629 (
            .O(N__13605),
            .I(N__13581));
    LocalMux I__1628 (
            .O(N__13600),
            .I(N__13581));
    LocalMux I__1627 (
            .O(N__13595),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1626 (
            .O(N__13592),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__1625 (
            .O(N__13589),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1624 (
            .O(N__13586),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__1623 (
            .O(N__13581),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    InMux I__1622 (
            .O(N__13570),
            .I(N__13567));
    LocalMux I__1621 (
            .O(N__13567),
            .I(N__13564));
    Span4Mux_h I__1620 (
            .O(N__13564),
            .I(N__13560));
    InMux I__1619 (
            .O(N__13563),
            .I(N__13557));
    Odrv4 I__1618 (
            .O(N__13560),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0 ));
    LocalMux I__1617 (
            .O(N__13557),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0 ));
    InMux I__1616 (
            .O(N__13552),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__1615 (
            .O(N__13549),
            .I(bfn_7_20_0_));
    InMux I__1614 (
            .O(N__13546),
            .I(N__13542));
    InMux I__1613 (
            .O(N__13545),
            .I(N__13539));
    LocalMux I__1612 (
            .O(N__13542),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0 ));
    LocalMux I__1611 (
            .O(N__13539),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0 ));
    InMux I__1610 (
            .O(N__13534),
            .I(N__13529));
    InMux I__1609 (
            .O(N__13533),
            .I(N__13526));
    InMux I__1608 (
            .O(N__13532),
            .I(N__13522));
    LocalMux I__1607 (
            .O(N__13529),
            .I(N__13519));
    LocalMux I__1606 (
            .O(N__13526),
            .I(N__13516));
    InMux I__1605 (
            .O(N__13525),
            .I(N__13513));
    LocalMux I__1604 (
            .O(N__13522),
            .I(N__13510));
    Span4Mux_v I__1603 (
            .O(N__13519),
            .I(N__13503));
    Span4Mux_h I__1602 (
            .O(N__13516),
            .I(N__13496));
    LocalMux I__1601 (
            .O(N__13513),
            .I(N__13496));
    Span4Mux_v I__1600 (
            .O(N__13510),
            .I(N__13496));
    InMux I__1599 (
            .O(N__13509),
            .I(N__13493));
    InMux I__1598 (
            .O(N__13508),
            .I(N__13486));
    InMux I__1597 (
            .O(N__13507),
            .I(N__13486));
    InMux I__1596 (
            .O(N__13506),
            .I(N__13486));
    Odrv4 I__1595 (
            .O(N__13503),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__1594 (
            .O(N__13496),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1593 (
            .O(N__13493),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1592 (
            .O(N__13486),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    CEMux I__1591 (
            .O(N__13477),
            .I(N__13473));
    CEMux I__1590 (
            .O(N__13476),
            .I(N__13469));
    LocalMux I__1589 (
            .O(N__13473),
            .I(N__13466));
    CEMux I__1588 (
            .O(N__13472),
            .I(N__13463));
    LocalMux I__1587 (
            .O(N__13469),
            .I(N__13460));
    Span4Mux_h I__1586 (
            .O(N__13466),
            .I(N__13455));
    LocalMux I__1585 (
            .O(N__13463),
            .I(N__13455));
    Span4Mux_v I__1584 (
            .O(N__13460),
            .I(N__13452));
    Span4Mux_h I__1583 (
            .O(N__13455),
            .I(N__13449));
    Odrv4 I__1582 (
            .O(N__13452),
            .I(\this_vga_signals.N_614_0 ));
    Odrv4 I__1581 (
            .O(N__13449),
            .I(\this_vga_signals.N_614_0 ));
    SRMux I__1580 (
            .O(N__13444),
            .I(N__13440));
    SRMux I__1579 (
            .O(N__13443),
            .I(N__13437));
    LocalMux I__1578 (
            .O(N__13440),
            .I(N__13433));
    LocalMux I__1577 (
            .O(N__13437),
            .I(N__13428));
    SRMux I__1576 (
            .O(N__13436),
            .I(N__13425));
    Span4Mux_v I__1575 (
            .O(N__13433),
            .I(N__13422));
    SRMux I__1574 (
            .O(N__13432),
            .I(N__13419));
    SRMux I__1573 (
            .O(N__13431),
            .I(N__13416));
    Span4Mux_h I__1572 (
            .O(N__13428),
            .I(N__13412));
    LocalMux I__1571 (
            .O(N__13425),
            .I(N__13409));
    Span4Mux_h I__1570 (
            .O(N__13422),
            .I(N__13404));
    LocalMux I__1569 (
            .O(N__13419),
            .I(N__13404));
    LocalMux I__1568 (
            .O(N__13416),
            .I(N__13401));
    InMux I__1567 (
            .O(N__13415),
            .I(N__13398));
    Odrv4 I__1566 (
            .O(N__13412),
            .I(\this_vga_signals.N_931_1 ));
    Odrv4 I__1565 (
            .O(N__13409),
            .I(\this_vga_signals.N_931_1 ));
    Odrv4 I__1564 (
            .O(N__13404),
            .I(\this_vga_signals.N_931_1 ));
    Odrv4 I__1563 (
            .O(N__13401),
            .I(\this_vga_signals.N_931_1 ));
    LocalMux I__1562 (
            .O(N__13398),
            .I(\this_vga_signals.N_931_1 ));
    CascadeMux I__1561 (
            .O(N__13387),
            .I(\this_vga_signals.vaddress_0_5_cascade_ ));
    InMux I__1560 (
            .O(N__13384),
            .I(N__13381));
    LocalMux I__1559 (
            .O(N__13381),
            .I(N__13375));
    InMux I__1558 (
            .O(N__13380),
            .I(N__13370));
    InMux I__1557 (
            .O(N__13379),
            .I(N__13370));
    InMux I__1556 (
            .O(N__13378),
            .I(N__13367));
    Odrv12 I__1555 (
            .O(N__13375),
            .I(\this_vga_signals.mult1_un75_sum_axb2 ));
    LocalMux I__1554 (
            .O(N__13370),
            .I(\this_vga_signals.mult1_un75_sum_axb2 ));
    LocalMux I__1553 (
            .O(N__13367),
            .I(\this_vga_signals.mult1_un75_sum_axb2 ));
    InMux I__1552 (
            .O(N__13360),
            .I(N__13356));
    InMux I__1551 (
            .O(N__13359),
            .I(N__13353));
    LocalMux I__1550 (
            .O(N__13356),
            .I(\this_vga_signals.mult1_un75_sum_axb1 ));
    LocalMux I__1549 (
            .O(N__13353),
            .I(\this_vga_signals.mult1_un75_sum_axb1 ));
    InMux I__1548 (
            .O(N__13348),
            .I(N__13345));
    LocalMux I__1547 (
            .O(N__13345),
            .I(N__13342));
    Span4Mux_h I__1546 (
            .O(N__13342),
            .I(N__13338));
    InMux I__1545 (
            .O(N__13341),
            .I(N__13335));
    Odrv4 I__1544 (
            .O(N__13338),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_d ));
    LocalMux I__1543 (
            .O(N__13335),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_d ));
    InMux I__1542 (
            .O(N__13330),
            .I(N__13325));
    InMux I__1541 (
            .O(N__13329),
            .I(N__13320));
    InMux I__1540 (
            .O(N__13328),
            .I(N__13320));
    LocalMux I__1539 (
            .O(N__13325),
            .I(N__13311));
    LocalMux I__1538 (
            .O(N__13320),
            .I(N__13307));
    InMux I__1537 (
            .O(N__13319),
            .I(N__13304));
    InMux I__1536 (
            .O(N__13318),
            .I(N__13299));
    InMux I__1535 (
            .O(N__13317),
            .I(N__13299));
    InMux I__1534 (
            .O(N__13316),
            .I(N__13292));
    InMux I__1533 (
            .O(N__13315),
            .I(N__13292));
    InMux I__1532 (
            .O(N__13314),
            .I(N__13292));
    Span4Mux_h I__1531 (
            .O(N__13311),
            .I(N__13289));
    InMux I__1530 (
            .O(N__13310),
            .I(N__13286));
    Odrv4 I__1529 (
            .O(N__13307),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__1528 (
            .O(N__13304),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__1527 (
            .O(N__13299),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__1526 (
            .O(N__13292),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__1525 (
            .O(N__13289),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__1524 (
            .O(N__13286),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    CascadeMux I__1523 (
            .O(N__13273),
            .I(N__13270));
    InMux I__1522 (
            .O(N__13270),
            .I(N__13266));
    CascadeMux I__1521 (
            .O(N__13269),
            .I(N__13260));
    LocalMux I__1520 (
            .O(N__13266),
            .I(N__13256));
    InMux I__1519 (
            .O(N__13265),
            .I(N__13251));
    InMux I__1518 (
            .O(N__13264),
            .I(N__13251));
    InMux I__1517 (
            .O(N__13263),
            .I(N__13248));
    InMux I__1516 (
            .O(N__13260),
            .I(N__13243));
    InMux I__1515 (
            .O(N__13259),
            .I(N__13243));
    Odrv4 I__1514 (
            .O(N__13256),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1513 (
            .O(N__13251),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1512 (
            .O(N__13248),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1511 (
            .O(N__13243),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    InMux I__1510 (
            .O(N__13234),
            .I(N__13231));
    LocalMux I__1509 (
            .O(N__13231),
            .I(N__13228));
    Odrv12 I__1508 (
            .O(N__13228),
            .I(\this_vga_signals.M_hcounter_d7lt4 ));
    CascadeMux I__1507 (
            .O(N__13225),
            .I(N__13219));
    InMux I__1506 (
            .O(N__13224),
            .I(N__13214));
    CascadeMux I__1505 (
            .O(N__13223),
            .I(N__13210));
    InMux I__1504 (
            .O(N__13222),
            .I(N__13204));
    InMux I__1503 (
            .O(N__13219),
            .I(N__13201));
    InMux I__1502 (
            .O(N__13218),
            .I(N__13196));
    InMux I__1501 (
            .O(N__13217),
            .I(N__13196));
    LocalMux I__1500 (
            .O(N__13214),
            .I(N__13191));
    InMux I__1499 (
            .O(N__13213),
            .I(N__13188));
    InMux I__1498 (
            .O(N__13210),
            .I(N__13181));
    InMux I__1497 (
            .O(N__13209),
            .I(N__13181));
    InMux I__1496 (
            .O(N__13208),
            .I(N__13181));
    InMux I__1495 (
            .O(N__13207),
            .I(N__13178));
    LocalMux I__1494 (
            .O(N__13204),
            .I(N__13170));
    LocalMux I__1493 (
            .O(N__13201),
            .I(N__13170));
    LocalMux I__1492 (
            .O(N__13196),
            .I(N__13170));
    InMux I__1491 (
            .O(N__13195),
            .I(N__13167));
    InMux I__1490 (
            .O(N__13194),
            .I(N__13164));
    Span4Mux_h I__1489 (
            .O(N__13191),
            .I(N__13161));
    LocalMux I__1488 (
            .O(N__13188),
            .I(N__13154));
    LocalMux I__1487 (
            .O(N__13181),
            .I(N__13154));
    LocalMux I__1486 (
            .O(N__13178),
            .I(N__13154));
    InMux I__1485 (
            .O(N__13177),
            .I(N__13151));
    Span4Mux_v I__1484 (
            .O(N__13170),
            .I(N__13146));
    LocalMux I__1483 (
            .O(N__13167),
            .I(N__13146));
    LocalMux I__1482 (
            .O(N__13164),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1481 (
            .O(N__13161),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1480 (
            .O(N__13154),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__1479 (
            .O(N__13151),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1478 (
            .O(N__13146),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__1477 (
            .O(N__13135),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    CascadeMux I__1476 (
            .O(N__13132),
            .I(N__13123));
    CascadeMux I__1475 (
            .O(N__13131),
            .I(N__13120));
    CascadeMux I__1474 (
            .O(N__13130),
            .I(N__13115));
    CascadeMux I__1473 (
            .O(N__13129),
            .I(N__13112));
    CascadeMux I__1472 (
            .O(N__13128),
            .I(N__13107));
    CascadeMux I__1471 (
            .O(N__13127),
            .I(N__13101));
    InMux I__1470 (
            .O(N__13126),
            .I(N__13094));
    InMux I__1469 (
            .O(N__13123),
            .I(N__13094));
    InMux I__1468 (
            .O(N__13120),
            .I(N__13094));
    InMux I__1467 (
            .O(N__13119),
            .I(N__13087));
    InMux I__1466 (
            .O(N__13118),
            .I(N__13087));
    InMux I__1465 (
            .O(N__13115),
            .I(N__13087));
    InMux I__1464 (
            .O(N__13112),
            .I(N__13084));
    InMux I__1463 (
            .O(N__13111),
            .I(N__13081));
    InMux I__1462 (
            .O(N__13110),
            .I(N__13078));
    InMux I__1461 (
            .O(N__13107),
            .I(N__13075));
    InMux I__1460 (
            .O(N__13106),
            .I(N__13068));
    InMux I__1459 (
            .O(N__13105),
            .I(N__13068));
    InMux I__1458 (
            .O(N__13104),
            .I(N__13068));
    InMux I__1457 (
            .O(N__13101),
            .I(N__13063));
    LocalMux I__1456 (
            .O(N__13094),
            .I(N__13052));
    LocalMux I__1455 (
            .O(N__13087),
            .I(N__13052));
    LocalMux I__1454 (
            .O(N__13084),
            .I(N__13052));
    LocalMux I__1453 (
            .O(N__13081),
            .I(N__13052));
    LocalMux I__1452 (
            .O(N__13078),
            .I(N__13052));
    LocalMux I__1451 (
            .O(N__13075),
            .I(N__13049));
    LocalMux I__1450 (
            .O(N__13068),
            .I(N__13046));
    CascadeMux I__1449 (
            .O(N__13067),
            .I(N__13043));
    InMux I__1448 (
            .O(N__13066),
            .I(N__13039));
    LocalMux I__1447 (
            .O(N__13063),
            .I(N__13036));
    Span4Mux_v I__1446 (
            .O(N__13052),
            .I(N__13031));
    Span4Mux_h I__1445 (
            .O(N__13049),
            .I(N__13031));
    Span4Mux_h I__1444 (
            .O(N__13046),
            .I(N__13028));
    InMux I__1443 (
            .O(N__13043),
            .I(N__13023));
    InMux I__1442 (
            .O(N__13042),
            .I(N__13023));
    LocalMux I__1441 (
            .O(N__13039),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1440 (
            .O(N__13036),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1439 (
            .O(N__13031),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1438 (
            .O(N__13028),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1437 (
            .O(N__13023),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__1436 (
            .O(N__13012),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    CascadeMux I__1435 (
            .O(N__13009),
            .I(N__13006));
    InMux I__1434 (
            .O(N__13006),
            .I(N__12992));
    InMux I__1433 (
            .O(N__13005),
            .I(N__12992));
    InMux I__1432 (
            .O(N__13004),
            .I(N__12989));
    InMux I__1431 (
            .O(N__13003),
            .I(N__12986));
    InMux I__1430 (
            .O(N__13002),
            .I(N__12981));
    InMux I__1429 (
            .O(N__13001),
            .I(N__12981));
    InMux I__1428 (
            .O(N__13000),
            .I(N__12978));
    InMux I__1427 (
            .O(N__12999),
            .I(N__12973));
    InMux I__1426 (
            .O(N__12998),
            .I(N__12973));
    InMux I__1425 (
            .O(N__12997),
            .I(N__12967));
    LocalMux I__1424 (
            .O(N__12992),
            .I(N__12962));
    LocalMux I__1423 (
            .O(N__12989),
            .I(N__12962));
    LocalMux I__1422 (
            .O(N__12986),
            .I(N__12953));
    LocalMux I__1421 (
            .O(N__12981),
            .I(N__12953));
    LocalMux I__1420 (
            .O(N__12978),
            .I(N__12953));
    LocalMux I__1419 (
            .O(N__12973),
            .I(N__12953));
    InMux I__1418 (
            .O(N__12972),
            .I(N__12943));
    InMux I__1417 (
            .O(N__12971),
            .I(N__12943));
    InMux I__1416 (
            .O(N__12970),
            .I(N__12943));
    LocalMux I__1415 (
            .O(N__12967),
            .I(N__12936));
    Span4Mux_h I__1414 (
            .O(N__12962),
            .I(N__12936));
    Span4Mux_v I__1413 (
            .O(N__12953),
            .I(N__12936));
    InMux I__1412 (
            .O(N__12952),
            .I(N__12933));
    InMux I__1411 (
            .O(N__12951),
            .I(N__12928));
    InMux I__1410 (
            .O(N__12950),
            .I(N__12928));
    LocalMux I__1409 (
            .O(N__12943),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1408 (
            .O(N__12936),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1407 (
            .O(N__12933),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1406 (
            .O(N__12928),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__1405 (
            .O(N__12919),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__1404 (
            .O(N__12916),
            .I(N__12907));
    InMux I__1403 (
            .O(N__12915),
            .I(N__12907));
    InMux I__1402 (
            .O(N__12914),
            .I(N__12904));
    InMux I__1401 (
            .O(N__12913),
            .I(N__12899));
    InMux I__1400 (
            .O(N__12912),
            .I(N__12899));
    LocalMux I__1399 (
            .O(N__12907),
            .I(N__12890));
    LocalMux I__1398 (
            .O(N__12904),
            .I(N__12890));
    LocalMux I__1397 (
            .O(N__12899),
            .I(N__12890));
    InMux I__1396 (
            .O(N__12898),
            .I(N__12887));
    InMux I__1395 (
            .O(N__12897),
            .I(N__12875));
    Span4Mux_v I__1394 (
            .O(N__12890),
            .I(N__12870));
    LocalMux I__1393 (
            .O(N__12887),
            .I(N__12870));
    InMux I__1392 (
            .O(N__12886),
            .I(N__12861));
    InMux I__1391 (
            .O(N__12885),
            .I(N__12861));
    InMux I__1390 (
            .O(N__12884),
            .I(N__12861));
    InMux I__1389 (
            .O(N__12883),
            .I(N__12861));
    InMux I__1388 (
            .O(N__12882),
            .I(N__12856));
    InMux I__1387 (
            .O(N__12881),
            .I(N__12856));
    InMux I__1386 (
            .O(N__12880),
            .I(N__12849));
    InMux I__1385 (
            .O(N__12879),
            .I(N__12849));
    InMux I__1384 (
            .O(N__12878),
            .I(N__12849));
    LocalMux I__1383 (
            .O(N__12875),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__1382 (
            .O(N__12870),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1381 (
            .O(N__12861),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1380 (
            .O(N__12856),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1379 (
            .O(N__12849),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    InMux I__1378 (
            .O(N__12838),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__1377 (
            .O(N__12835),
            .I(N__12827));
    InMux I__1376 (
            .O(N__12834),
            .I(N__12827));
    InMux I__1375 (
            .O(N__12833),
            .I(N__12818));
    InMux I__1374 (
            .O(N__12832),
            .I(N__12818));
    LocalMux I__1373 (
            .O(N__12827),
            .I(N__12814));
    CascadeMux I__1372 (
            .O(N__12826),
            .I(N__12810));
    InMux I__1371 (
            .O(N__12825),
            .I(N__12805));
    InMux I__1370 (
            .O(N__12824),
            .I(N__12805));
    InMux I__1369 (
            .O(N__12823),
            .I(N__12802));
    LocalMux I__1368 (
            .O(N__12818),
            .I(N__12799));
    CascadeMux I__1367 (
            .O(N__12817),
            .I(N__12794));
    Span4Mux_v I__1366 (
            .O(N__12814),
            .I(N__12788));
    InMux I__1365 (
            .O(N__12813),
            .I(N__12785));
    InMux I__1364 (
            .O(N__12810),
            .I(N__12782));
    LocalMux I__1363 (
            .O(N__12805),
            .I(N__12779));
    LocalMux I__1362 (
            .O(N__12802),
            .I(N__12774));
    Span4Mux_h I__1361 (
            .O(N__12799),
            .I(N__12774));
    InMux I__1360 (
            .O(N__12798),
            .I(N__12771));
    InMux I__1359 (
            .O(N__12797),
            .I(N__12766));
    InMux I__1358 (
            .O(N__12794),
            .I(N__12766));
    InMux I__1357 (
            .O(N__12793),
            .I(N__12759));
    InMux I__1356 (
            .O(N__12792),
            .I(N__12759));
    InMux I__1355 (
            .O(N__12791),
            .I(N__12759));
    Odrv4 I__1354 (
            .O(N__12788),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1353 (
            .O(N__12785),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1352 (
            .O(N__12782),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1351 (
            .O(N__12779),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1350 (
            .O(N__12774),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1349 (
            .O(N__12771),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1348 (
            .O(N__12766),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1347 (
            .O(N__12759),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    InMux I__1346 (
            .O(N__12742),
            .I(N__12736));
    InMux I__1345 (
            .O(N__12741),
            .I(N__12736));
    LocalMux I__1344 (
            .O(N__12736),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0 ));
    InMux I__1343 (
            .O(N__12733),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__1342 (
            .O(N__12730),
            .I(N__12727));
    LocalMux I__1341 (
            .O(N__12727),
            .I(N__12722));
    InMux I__1340 (
            .O(N__12726),
            .I(N__12714));
    InMux I__1339 (
            .O(N__12725),
            .I(N__12711));
    Span4Mux_v I__1338 (
            .O(N__12722),
            .I(N__12708));
    InMux I__1337 (
            .O(N__12721),
            .I(N__12705));
    InMux I__1336 (
            .O(N__12720),
            .I(N__12696));
    InMux I__1335 (
            .O(N__12719),
            .I(N__12696));
    InMux I__1334 (
            .O(N__12718),
            .I(N__12696));
    InMux I__1333 (
            .O(N__12717),
            .I(N__12696));
    LocalMux I__1332 (
            .O(N__12714),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1331 (
            .O(N__12711),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__1330 (
            .O(N__12708),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1329 (
            .O(N__12705),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1328 (
            .O(N__12696),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__1327 (
            .O(N__12685),
            .I(N__12682));
    LocalMux I__1326 (
            .O(N__12682),
            .I(N__12679));
    Span4Mux_h I__1325 (
            .O(N__12679),
            .I(N__12675));
    InMux I__1324 (
            .O(N__12678),
            .I(N__12672));
    Odrv4 I__1323 (
            .O(N__12675),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0 ));
    LocalMux I__1322 (
            .O(N__12672),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0 ));
    InMux I__1321 (
            .O(N__12667),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    CascadeMux I__1320 (
            .O(N__12664),
            .I(\this_vga_signals.if_m7_0_x4_0_cascade_ ));
    CascadeMux I__1319 (
            .O(N__12661),
            .I(\this_vga_signals.if_N_9_1_cascade_ ));
    InMux I__1318 (
            .O(N__12658),
            .I(N__12653));
    InMux I__1317 (
            .O(N__12657),
            .I(N__12648));
    InMux I__1316 (
            .O(N__12656),
            .I(N__12648));
    LocalMux I__1315 (
            .O(N__12653),
            .I(\this_vga_signals.mult1_un75_sum_c2_0 ));
    LocalMux I__1314 (
            .O(N__12648),
            .I(\this_vga_signals.mult1_un75_sum_c2_0 ));
    CascadeMux I__1313 (
            .O(N__12643),
            .I(N__12640));
    InMux I__1312 (
            .O(N__12640),
            .I(N__12637));
    LocalMux I__1311 (
            .O(N__12637),
            .I(\this_vga_signals.mult1_un82_sum_c3 ));
    CascadeMux I__1310 (
            .O(N__12634),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_cascade_ ));
    InMux I__1309 (
            .O(N__12631),
            .I(N__12628));
    LocalMux I__1308 (
            .O(N__12628),
            .I(\this_vga_signals.mult1_un89_sum_c3 ));
    CascadeMux I__1307 (
            .O(N__12625),
            .I(N__12622));
    InMux I__1306 (
            .O(N__12622),
            .I(N__12619));
    LocalMux I__1305 (
            .O(N__12619),
            .I(N__12616));
    Span12Mux_h I__1304 (
            .O(N__12616),
            .I(N__12613));
    Odrv12 I__1303 (
            .O(N__12613),
            .I(M_this_vga_signals_address_0));
    InMux I__1302 (
            .O(N__12610),
            .I(N__12607));
    LocalMux I__1301 (
            .O(N__12607),
            .I(\this_vga_signals.d_N_12 ));
    InMux I__1300 (
            .O(N__12604),
            .I(N__12601));
    LocalMux I__1299 (
            .O(N__12601),
            .I(\this_vga_signals.d_N_11 ));
    CascadeMux I__1298 (
            .O(N__12598),
            .I(N__12595));
    InMux I__1297 (
            .O(N__12595),
            .I(N__12592));
    LocalMux I__1296 (
            .O(N__12592),
            .I(N__12589));
    Odrv4 I__1295 (
            .O(N__12589),
            .I(\this_vga_signals.M_hcounter_q_RNIUAKU9Z0Z_4 ));
    InMux I__1294 (
            .O(N__12586),
            .I(N__12583));
    LocalMux I__1293 (
            .O(N__12583),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_0 ));
    InMux I__1292 (
            .O(N__12580),
            .I(N__12576));
    InMux I__1291 (
            .O(N__12579),
            .I(N__12569));
    LocalMux I__1290 (
            .O(N__12576),
            .I(N__12566));
    InMux I__1289 (
            .O(N__12575),
            .I(N__12557));
    InMux I__1288 (
            .O(N__12574),
            .I(N__12557));
    InMux I__1287 (
            .O(N__12573),
            .I(N__12557));
    InMux I__1286 (
            .O(N__12572),
            .I(N__12557));
    LocalMux I__1285 (
            .O(N__12569),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    Odrv4 I__1284 (
            .O(N__12566),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__1283 (
            .O(N__12557),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    InMux I__1282 (
            .O(N__12550),
            .I(N__12547));
    LocalMux I__1281 (
            .O(N__12547),
            .I(\this_vga_signals.N_2_7_0 ));
    InMux I__1280 (
            .O(N__12544),
            .I(N__12540));
    InMux I__1279 (
            .O(N__12543),
            .I(N__12537));
    LocalMux I__1278 (
            .O(N__12540),
            .I(\this_vga_signals.N_236 ));
    LocalMux I__1277 (
            .O(N__12537),
            .I(\this_vga_signals.N_236 ));
    InMux I__1276 (
            .O(N__12532),
            .I(N__12529));
    LocalMux I__1275 (
            .O(N__12529),
            .I(N__12525));
    InMux I__1274 (
            .O(N__12528),
            .I(N__12520));
    Span4Mux_v I__1273 (
            .O(N__12525),
            .I(N__12517));
    InMux I__1272 (
            .O(N__12524),
            .I(N__12514));
    InMux I__1271 (
            .O(N__12523),
            .I(N__12511));
    LocalMux I__1270 (
            .O(N__12520),
            .I(\this_vga_signals.SUM_3_i_0_0_3 ));
    Odrv4 I__1269 (
            .O(N__12517),
            .I(\this_vga_signals.SUM_3_i_0_0_3 ));
    LocalMux I__1268 (
            .O(N__12514),
            .I(\this_vga_signals.SUM_3_i_0_0_3 ));
    LocalMux I__1267 (
            .O(N__12511),
            .I(\this_vga_signals.SUM_3_i_0_0_3 ));
    CascadeMux I__1266 (
            .O(N__12502),
            .I(N__12499));
    InMux I__1265 (
            .O(N__12499),
            .I(N__12496));
    LocalMux I__1264 (
            .O(N__12496),
            .I(N__12493));
    Span4Mux_v I__1263 (
            .O(N__12493),
            .I(N__12490));
    Odrv4 I__1262 (
            .O(N__12490),
            .I(\this_vga_signals.g0_1 ));
    CascadeMux I__1261 (
            .O(N__12487),
            .I(\this_vga_signals.un6_vvisibilitylt8_cascade_ ));
    CascadeMux I__1260 (
            .O(N__12484),
            .I(\this_vga_signals.vvisibility_1_cascade_ ));
    InMux I__1259 (
            .O(N__12481),
            .I(N__12478));
    LocalMux I__1258 (
            .O(N__12478),
            .I(N__12475));
    Odrv4 I__1257 (
            .O(N__12475),
            .I(\this_vga_signals.vsync_1_3 ));
    CascadeMux I__1256 (
            .O(N__12472),
            .I(\this_vga_signals.vsync_1_2_cascade_ ));
    IoInMux I__1255 (
            .O(N__12469),
            .I(N__12466));
    LocalMux I__1254 (
            .O(N__12466),
            .I(N__12463));
    IoSpan4Mux I__1253 (
            .O(N__12463),
            .I(N__12460));
    Span4Mux_s2_v I__1252 (
            .O(N__12460),
            .I(N__12457));
    Sp12to4 I__1251 (
            .O(N__12457),
            .I(N__12454));
    Span12Mux_s10_v I__1250 (
            .O(N__12454),
            .I(N__12451));
    Odrv12 I__1249 (
            .O(N__12451),
            .I(this_vga_signals_vsync_1_i));
    InMux I__1248 (
            .O(N__12448),
            .I(N__12440));
    InMux I__1247 (
            .O(N__12447),
            .I(N__12437));
    CascadeMux I__1246 (
            .O(N__12446),
            .I(N__12434));
    InMux I__1245 (
            .O(N__12445),
            .I(N__12431));
    CascadeMux I__1244 (
            .O(N__12444),
            .I(N__12428));
    CascadeMux I__1243 (
            .O(N__12443),
            .I(N__12425));
    LocalMux I__1242 (
            .O(N__12440),
            .I(N__12420));
    LocalMux I__1241 (
            .O(N__12437),
            .I(N__12420));
    InMux I__1240 (
            .O(N__12434),
            .I(N__12417));
    LocalMux I__1239 (
            .O(N__12431),
            .I(N__12414));
    InMux I__1238 (
            .O(N__12428),
            .I(N__12409));
    InMux I__1237 (
            .O(N__12425),
            .I(N__12409));
    Odrv4 I__1236 (
            .O(N__12420),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9 ));
    LocalMux I__1235 (
            .O(N__12417),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9 ));
    Odrv4 I__1234 (
            .O(N__12414),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9 ));
    LocalMux I__1233 (
            .O(N__12409),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9 ));
    InMux I__1232 (
            .O(N__12400),
            .I(N__12397));
    LocalMux I__1231 (
            .O(N__12397),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1 ));
    InMux I__1230 (
            .O(N__12394),
            .I(N__12391));
    LocalMux I__1229 (
            .O(N__12391),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_7 ));
    CascadeMux I__1228 (
            .O(N__12388),
            .I(N__12384));
    InMux I__1227 (
            .O(N__12387),
            .I(N__12381));
    InMux I__1226 (
            .O(N__12384),
            .I(N__12378));
    LocalMux I__1225 (
            .O(N__12381),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_8 ));
    LocalMux I__1224 (
            .O(N__12378),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_8 ));
    CascadeMux I__1223 (
            .O(N__12373),
            .I(N__12370));
    InMux I__1222 (
            .O(N__12370),
            .I(N__12367));
    LocalMux I__1221 (
            .O(N__12367),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_9 ));
    InMux I__1220 (
            .O(N__12364),
            .I(N__12360));
    InMux I__1219 (
            .O(N__12363),
            .I(N__12357));
    LocalMux I__1218 (
            .O(N__12360),
            .I(N__12354));
    LocalMux I__1217 (
            .O(N__12357),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_6 ));
    Odrv4 I__1216 (
            .O(N__12354),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_6 ));
    CascadeMux I__1215 (
            .O(N__12349),
            .I(\this_vga_signals.SUM_3_i_0_0_3_cascade_ ));
    InMux I__1214 (
            .O(N__12346),
            .I(N__12342));
    InMux I__1213 (
            .O(N__12345),
            .I(N__12339));
    LocalMux I__1212 (
            .O(N__12342),
            .I(N__12333));
    LocalMux I__1211 (
            .O(N__12339),
            .I(N__12333));
    InMux I__1210 (
            .O(N__12338),
            .I(N__12330));
    Odrv4 I__1209 (
            .O(N__12333),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ));
    LocalMux I__1208 (
            .O(N__12330),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ));
    CascadeMux I__1207 (
            .O(N__12325),
            .I(N__12321));
    CascadeMux I__1206 (
            .O(N__12324),
            .I(N__12317));
    InMux I__1205 (
            .O(N__12321),
            .I(N__12314));
    InMux I__1204 (
            .O(N__12320),
            .I(N__12310));
    InMux I__1203 (
            .O(N__12317),
            .I(N__12307));
    LocalMux I__1202 (
            .O(N__12314),
            .I(N__12304));
    InMux I__1201 (
            .O(N__12313),
            .I(N__12301));
    LocalMux I__1200 (
            .O(N__12310),
            .I(N__12296));
    LocalMux I__1199 (
            .O(N__12307),
            .I(N__12296));
    Odrv12 I__1198 (
            .O(N__12304),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    LocalMux I__1197 (
            .O(N__12301),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    Odrv4 I__1196 (
            .O(N__12296),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    CascadeMux I__1195 (
            .O(N__12289),
            .I(\this_vga_signals.mult1_un61_sum_axb1_cascade_ ));
    CascadeMux I__1194 (
            .O(N__12286),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_cascade_ ));
    InMux I__1193 (
            .O(N__12283),
            .I(N__12280));
    LocalMux I__1192 (
            .O(N__12280),
            .I(\this_vga_signals.mult1_un75_sum_axb2_1 ));
    CascadeMux I__1191 (
            .O(N__12277),
            .I(\this_vga_signals.N_236_cascade_ ));
    InMux I__1190 (
            .O(N__12274),
            .I(N__12271));
    LocalMux I__1189 (
            .O(N__12271),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_0 ));
    CascadeMux I__1188 (
            .O(N__12268),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_ ));
    CascadeMux I__1187 (
            .O(N__12265),
            .I(\this_vga_signals.N_3_2_1_cascade_ ));
    InMux I__1186 (
            .O(N__12262),
            .I(N__12259));
    LocalMux I__1185 (
            .O(N__12259),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0 ));
    CascadeMux I__1184 (
            .O(N__12256),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_0_0_cascade_ ));
    InMux I__1183 (
            .O(N__12253),
            .I(N__12250));
    LocalMux I__1182 (
            .O(N__12250),
            .I(\this_vga_signals.g2_0_0 ));
    InMux I__1181 (
            .O(N__12247),
            .I(N__12244));
    LocalMux I__1180 (
            .O(N__12244),
            .I(\this_vga_signals.if_N_9_0_0 ));
    InMux I__1179 (
            .O(N__12241),
            .I(N__12237));
    InMux I__1178 (
            .O(N__12240),
            .I(N__12234));
    LocalMux I__1177 (
            .O(N__12237),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    LocalMux I__1176 (
            .O(N__12234),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    CascadeMux I__1175 (
            .O(N__12229),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ));
    CascadeMux I__1174 (
            .O(N__12226),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_cascade_ ));
    IoInMux I__1173 (
            .O(N__12223),
            .I(N__12220));
    LocalMux I__1172 (
            .O(N__12220),
            .I(N__12217));
    Odrv12 I__1171 (
            .O(N__12217),
            .I(this_vga_signals_vvisibility_i));
    InMux I__1170 (
            .O(N__12214),
            .I(N__12210));
    InMux I__1169 (
            .O(N__12213),
            .I(N__12207));
    LocalMux I__1168 (
            .O(N__12210),
            .I(N__12204));
    LocalMux I__1167 (
            .O(N__12207),
            .I(\this_vga_signals.N_5_i_5 ));
    Odrv4 I__1166 (
            .O(N__12204),
            .I(\this_vga_signals.N_5_i_5 ));
    InMux I__1165 (
            .O(N__12199),
            .I(N__12196));
    LocalMux I__1164 (
            .O(N__12196),
            .I(N__12193));
    Odrv4 I__1163 (
            .O(N__12193),
            .I(\this_vga_signals.mult1_un82_sum_c3_0 ));
    CascadeMux I__1162 (
            .O(N__12190),
            .I(\this_vga_signals.g0_4_cascade_ ));
    CascadeMux I__1161 (
            .O(N__12187),
            .I(\this_vga_signals.g0_7_0_cascade_ ));
    CascadeMux I__1160 (
            .O(N__12184),
            .I(N__12181));
    InMux I__1159 (
            .O(N__12181),
            .I(N__12178));
    LocalMux I__1158 (
            .O(N__12178),
            .I(N__12175));
    Span4Mux_v I__1157 (
            .O(N__12175),
            .I(N__12172));
    Sp12to4 I__1156 (
            .O(N__12172),
            .I(N__12169));
    Span12Mux_h I__1155 (
            .O(N__12169),
            .I(N__12166));
    Odrv12 I__1154 (
            .O(N__12166),
            .I(M_this_vga_signals_address_1));
    InMux I__1153 (
            .O(N__12163),
            .I(N__12160));
    LocalMux I__1152 (
            .O(N__12160),
            .I(N__12157));
    Odrv4 I__1151 (
            .O(N__12157),
            .I(\this_vga_ramdac.N_24_mux ));
    InMux I__1150 (
            .O(N__12154),
            .I(N__12150));
    InMux I__1149 (
            .O(N__12153),
            .I(N__12147));
    LocalMux I__1148 (
            .O(N__12150),
            .I(N__12144));
    LocalMux I__1147 (
            .O(N__12147),
            .I(N__12141));
    Odrv4 I__1146 (
            .O(N__12144),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ));
    Odrv4 I__1145 (
            .O(N__12141),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ));
    InMux I__1144 (
            .O(N__12136),
            .I(N__12133));
    LocalMux I__1143 (
            .O(N__12133),
            .I(\this_vga_signals.g1 ));
    InMux I__1142 (
            .O(N__12130),
            .I(N__12127));
    LocalMux I__1141 (
            .O(N__12127),
            .I(N__12124));
    Odrv4 I__1140 (
            .O(N__12124),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_0_0 ));
    InMux I__1139 (
            .O(N__12121),
            .I(N__12118));
    LocalMux I__1138 (
            .O(N__12118),
            .I(\this_vga_signals.un2_hsynclt6_0 ));
    InMux I__1137 (
            .O(N__12115),
            .I(N__12109));
    InMux I__1136 (
            .O(N__12114),
            .I(N__12109));
    LocalMux I__1135 (
            .O(N__12109),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_1 ));
    CascadeMux I__1134 (
            .O(N__12106),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_ ));
    CascadeMux I__1133 (
            .O(N__12103),
            .I(\this_vga_signals.M_hcounter_d7lt7_0_cascade_ ));
    InMux I__1132 (
            .O(N__12100),
            .I(N__12097));
    LocalMux I__1131 (
            .O(N__12097),
            .I(\this_vga_signals.M_hcounter_d7lto7_1 ));
    CascadeMux I__1130 (
            .O(N__12094),
            .I(\this_vga_signals.mult1_un61_sum_0_3_cascade_ ));
    IoInMux I__1129 (
            .O(N__12091),
            .I(N__12088));
    LocalMux I__1128 (
            .O(N__12088),
            .I(N__12085));
    Odrv12 I__1127 (
            .O(N__12085),
            .I(\this_vga_signals.N_614_1 ));
    InMux I__1126 (
            .O(N__12082),
            .I(N__12079));
    LocalMux I__1125 (
            .O(N__12079),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_0 ));
    CascadeMux I__1124 (
            .O(N__12076),
            .I(\this_vga_signals.g0_i_x4_0_cascade_ ));
    InMux I__1123 (
            .O(N__12073),
            .I(N__12070));
    LocalMux I__1122 (
            .O(N__12070),
            .I(N__12067));
    Odrv4 I__1121 (
            .O(N__12067),
            .I(\this_vga_signals.g0_i_x4_2 ));
    CascadeMux I__1120 (
            .O(N__12064),
            .I(\this_vga_signals.N_931_1_cascade_ ));
    IoInMux I__1119 (
            .O(N__12061),
            .I(N__12058));
    LocalMux I__1118 (
            .O(N__12058),
            .I(N__12055));
    Span12Mux_s8_v I__1117 (
            .O(N__12055),
            .I(N__12052));
    Span12Mux_h I__1116 (
            .O(N__12052),
            .I(N__12048));
    InMux I__1115 (
            .O(N__12051),
            .I(N__12045));
    Odrv12 I__1114 (
            .O(N__12048),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI0JBR6Z0Z_9 ));
    LocalMux I__1113 (
            .O(N__12045),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI0JBR6Z0Z_9 ));
    InMux I__1112 (
            .O(N__12040),
            .I(N__12037));
    LocalMux I__1111 (
            .O(N__12037),
            .I(\this_vga_signals.un4_hsynclto3_0 ));
    CascadeMux I__1110 (
            .O(N__12034),
            .I(\this_vga_signals.un2_hsynclt7_cascade_ ));
    InMux I__1109 (
            .O(N__12031),
            .I(N__12028));
    LocalMux I__1108 (
            .O(N__12028),
            .I(\this_vga_signals.hsync_1_0 ));
    IoInMux I__1107 (
            .O(N__12025),
            .I(N__12022));
    LocalMux I__1106 (
            .O(N__12022),
            .I(N__12019));
    Span4Mux_s0_v I__1105 (
            .O(N__12019),
            .I(N__12016));
    Span4Mux_v I__1104 (
            .O(N__12016),
            .I(N__12013));
    Span4Mux_v I__1103 (
            .O(N__12013),
            .I(N__12010));
    Span4Mux_v I__1102 (
            .O(N__12010),
            .I(N__12007));
    Odrv4 I__1101 (
            .O(N__12007),
            .I(this_vga_signals_hvisibility_i));
    CascadeMux I__1100 (
            .O(N__12004),
            .I(\this_vga_signals.if_N_8_i_0_cascade_ ));
    CascadeMux I__1099 (
            .O(N__12001),
            .I(\this_vga_signals.if_N_9_0_0_cascade_ ));
    InMux I__1098 (
            .O(N__11998),
            .I(N__11994));
    InMux I__1097 (
            .O(N__11997),
            .I(N__11991));
    LocalMux I__1096 (
            .O(N__11994),
            .I(N__11988));
    LocalMux I__1095 (
            .O(N__11991),
            .I(\this_pixel_clk.M_counter_q_i_1 ));
    Odrv4 I__1094 (
            .O(N__11988),
            .I(\this_pixel_clk.M_counter_q_i_1 ));
    InMux I__1093 (
            .O(N__11983),
            .I(N__11978));
    InMux I__1092 (
            .O(N__11982),
            .I(N__11975));
    InMux I__1091 (
            .O(N__11981),
            .I(N__11972));
    LocalMux I__1090 (
            .O(N__11978),
            .I(\this_pixel_clk.M_counter_qZ0Z_0 ));
    LocalMux I__1089 (
            .O(N__11975),
            .I(\this_pixel_clk.M_counter_qZ0Z_0 ));
    LocalMux I__1088 (
            .O(N__11972),
            .I(\this_pixel_clk.M_counter_qZ0Z_0 ));
    IoInMux I__1087 (
            .O(N__11965),
            .I(N__11962));
    LocalMux I__1086 (
            .O(N__11962),
            .I(N__11959));
    Span4Mux_s2_h I__1085 (
            .O(N__11959),
            .I(N__11956));
    Sp12to4 I__1084 (
            .O(N__11956),
            .I(N__11953));
    Odrv12 I__1083 (
            .O(N__11953),
            .I(rgb_c_3));
    IoInMux I__1082 (
            .O(N__11950),
            .I(N__11947));
    LocalMux I__1081 (
            .O(N__11947),
            .I(N__11944));
    Span4Mux_s2_h I__1080 (
            .O(N__11944),
            .I(N__11941));
    Span4Mux_v I__1079 (
            .O(N__11941),
            .I(N__11938));
    Span4Mux_v I__1078 (
            .O(N__11938),
            .I(N__11935));
    Odrv4 I__1077 (
            .O(N__11935),
            .I(rgb_c_4));
    CascadeMux I__1076 (
            .O(N__11932),
            .I(N__11928));
    InMux I__1075 (
            .O(N__11931),
            .I(N__11925));
    InMux I__1074 (
            .O(N__11928),
            .I(N__11922));
    LocalMux I__1073 (
            .O(N__11925),
            .I(\this_vga_ramdac.N_2870_reto ));
    LocalMux I__1072 (
            .O(N__11922),
            .I(\this_vga_ramdac.N_2870_reto ));
    IoInMux I__1071 (
            .O(N__11917),
            .I(N__11914));
    LocalMux I__1070 (
            .O(N__11914),
            .I(N__11911));
    Odrv12 I__1069 (
            .O(N__11911),
            .I(rgb_c_2));
    InMux I__1068 (
            .O(N__11908),
            .I(N__11905));
    LocalMux I__1067 (
            .O(N__11905),
            .I(\this_vga_ramdac.i2_mux_0 ));
    InMux I__1066 (
            .O(N__11902),
            .I(N__11898));
    CascadeMux I__1065 (
            .O(N__11901),
            .I(N__11895));
    LocalMux I__1064 (
            .O(N__11898),
            .I(N__11892));
    InMux I__1063 (
            .O(N__11895),
            .I(N__11889));
    Odrv4 I__1062 (
            .O(N__11892),
            .I(\this_vga_ramdac.N_2875_reto ));
    LocalMux I__1061 (
            .O(N__11889),
            .I(\this_vga_ramdac.N_2875_reto ));
    CascadeMux I__1060 (
            .O(N__11884),
            .I(\this_vga_signals.un4_hsynclto7_0_cascade_ ));
    IoInMux I__1059 (
            .O(N__11881),
            .I(N__11878));
    LocalMux I__1058 (
            .O(N__11878),
            .I(N__11875));
    IoSpan4Mux I__1057 (
            .O(N__11875),
            .I(N__11872));
    Span4Mux_s3_v I__1056 (
            .O(N__11872),
            .I(N__11869));
    Sp12to4 I__1055 (
            .O(N__11869),
            .I(N__11866));
    Odrv12 I__1054 (
            .O(N__11866),
            .I(this_vga_signals_hsync_1_i));
    IoInMux I__1053 (
            .O(N__11863),
            .I(N__11860));
    LocalMux I__1052 (
            .O(N__11860),
            .I(N__11857));
    Span4Mux_s0_h I__1051 (
            .O(N__11857),
            .I(N__11854));
    Span4Mux_v I__1050 (
            .O(N__11854),
            .I(N__11851));
    Odrv4 I__1049 (
            .O(N__11851),
            .I(port_nmib_0_i));
    InMux I__1048 (
            .O(N__11848),
            .I(N__11845));
    LocalMux I__1047 (
            .O(N__11845),
            .I(N__11842));
    Span4Mux_v I__1046 (
            .O(N__11842),
            .I(N__11839));
    Odrv4 I__1045 (
            .O(N__11839),
            .I(port_clk_c));
    InMux I__1044 (
            .O(N__11836),
            .I(N__11833));
    LocalMux I__1043 (
            .O(N__11833),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    IoInMux I__1042 (
            .O(N__11830),
            .I(N__11827));
    LocalMux I__1041 (
            .O(N__11827),
            .I(N__11824));
    IoSpan4Mux I__1040 (
            .O(N__11824),
            .I(N__11821));
    Span4Mux_s1_h I__1039 (
            .O(N__11821),
            .I(N__11818));
    Span4Mux_v I__1038 (
            .O(N__11818),
            .I(N__11815));
    Odrv4 I__1037 (
            .O(N__11815),
            .I(rgb_c_5));
    IoInMux I__1036 (
            .O(N__11812),
            .I(N__11809));
    LocalMux I__1035 (
            .O(N__11809),
            .I(N__11806));
    IoSpan4Mux I__1034 (
            .O(N__11806),
            .I(N__11803));
    Span4Mux_s1_h I__1033 (
            .O(N__11803),
            .I(N__11800));
    Odrv4 I__1032 (
            .O(N__11800),
            .I(port_data_rw_0_i));
    IoInMux I__1031 (
            .O(N__11797),
            .I(N__11794));
    LocalMux I__1030 (
            .O(N__11794),
            .I(N__11791));
    Span4Mux_s2_h I__1029 (
            .O(N__11791),
            .I(N__11788));
    Sp12to4 I__1028 (
            .O(N__11788),
            .I(N__11785));
    Odrv12 I__1027 (
            .O(N__11785),
            .I(rgb_c_0));
    IoInMux I__1026 (
            .O(N__11782),
            .I(N__11779));
    LocalMux I__1025 (
            .O(N__11779),
            .I(N__11776));
    Odrv4 I__1024 (
            .O(N__11776),
            .I(rgb_c_1));
    CascadeMux I__1023 (
            .O(N__11773),
            .I(N__11770));
    CascadeBuf I__1022 (
            .O(N__11770),
            .I(N__11767));
    CascadeMux I__1021 (
            .O(N__11767),
            .I(N__11764));
    CascadeBuf I__1020 (
            .O(N__11764),
            .I(N__11761));
    CascadeMux I__1019 (
            .O(N__11761),
            .I(N__11758));
    CascadeBuf I__1018 (
            .O(N__11758),
            .I(N__11755));
    CascadeMux I__1017 (
            .O(N__11755),
            .I(N__11752));
    CascadeBuf I__1016 (
            .O(N__11752),
            .I(N__11749));
    CascadeMux I__1015 (
            .O(N__11749),
            .I(N__11746));
    CascadeBuf I__1014 (
            .O(N__11746),
            .I(N__11743));
    CascadeMux I__1013 (
            .O(N__11743),
            .I(N__11740));
    CascadeBuf I__1012 (
            .O(N__11740),
            .I(N__11737));
    CascadeMux I__1011 (
            .O(N__11737),
            .I(N__11734));
    CascadeBuf I__1010 (
            .O(N__11734),
            .I(N__11731));
    CascadeMux I__1009 (
            .O(N__11731),
            .I(N__11728));
    CascadeBuf I__1008 (
            .O(N__11728),
            .I(N__11725));
    CascadeMux I__1007 (
            .O(N__11725),
            .I(N__11722));
    CascadeBuf I__1006 (
            .O(N__11722),
            .I(N__11719));
    CascadeMux I__1005 (
            .O(N__11719),
            .I(N__11716));
    CascadeBuf I__1004 (
            .O(N__11716),
            .I(N__11713));
    CascadeMux I__1003 (
            .O(N__11713),
            .I(N__11710));
    CascadeBuf I__1002 (
            .O(N__11710),
            .I(N__11707));
    CascadeMux I__1001 (
            .O(N__11707),
            .I(N__11704));
    CascadeBuf I__1000 (
            .O(N__11704),
            .I(N__11701));
    CascadeMux I__999 (
            .O(N__11701),
            .I(N__11698));
    CascadeBuf I__998 (
            .O(N__11698),
            .I(N__11695));
    CascadeMux I__997 (
            .O(N__11695),
            .I(N__11692));
    CascadeBuf I__996 (
            .O(N__11692),
            .I(N__11689));
    CascadeMux I__995 (
            .O(N__11689),
            .I(N__11686));
    CascadeBuf I__994 (
            .O(N__11686),
            .I(N__11683));
    CascadeMux I__993 (
            .O(N__11683),
            .I(N__11680));
    InMux I__992 (
            .O(N__11680),
            .I(N__11677));
    LocalMux I__991 (
            .O(N__11677),
            .I(N__11674));
    Span12Mux_h I__990 (
            .O(N__11674),
            .I(N__11671));
    Span12Mux_h I__989 (
            .O(N__11671),
            .I(N__11668));
    Odrv12 I__988 (
            .O(N__11668),
            .I(M_this_ppu_sprites_addr_9));
    CascadeMux I__987 (
            .O(N__11665),
            .I(N__11662));
    CascadeBuf I__986 (
            .O(N__11662),
            .I(N__11659));
    CascadeMux I__985 (
            .O(N__11659),
            .I(N__11656));
    CascadeBuf I__984 (
            .O(N__11656),
            .I(N__11653));
    CascadeMux I__983 (
            .O(N__11653),
            .I(N__11650));
    CascadeBuf I__982 (
            .O(N__11650),
            .I(N__11647));
    CascadeMux I__981 (
            .O(N__11647),
            .I(N__11644));
    CascadeBuf I__980 (
            .O(N__11644),
            .I(N__11641));
    CascadeMux I__979 (
            .O(N__11641),
            .I(N__11638));
    CascadeBuf I__978 (
            .O(N__11638),
            .I(N__11635));
    CascadeMux I__977 (
            .O(N__11635),
            .I(N__11632));
    CascadeBuf I__976 (
            .O(N__11632),
            .I(N__11629));
    CascadeMux I__975 (
            .O(N__11629),
            .I(N__11626));
    CascadeBuf I__974 (
            .O(N__11626),
            .I(N__11623));
    CascadeMux I__973 (
            .O(N__11623),
            .I(N__11620));
    CascadeBuf I__972 (
            .O(N__11620),
            .I(N__11617));
    CascadeMux I__971 (
            .O(N__11617),
            .I(N__11614));
    CascadeBuf I__970 (
            .O(N__11614),
            .I(N__11611));
    CascadeMux I__969 (
            .O(N__11611),
            .I(N__11608));
    CascadeBuf I__968 (
            .O(N__11608),
            .I(N__11605));
    CascadeMux I__967 (
            .O(N__11605),
            .I(N__11602));
    CascadeBuf I__966 (
            .O(N__11602),
            .I(N__11599));
    CascadeMux I__965 (
            .O(N__11599),
            .I(N__11596));
    CascadeBuf I__964 (
            .O(N__11596),
            .I(N__11593));
    CascadeMux I__963 (
            .O(N__11593),
            .I(N__11590));
    CascadeBuf I__962 (
            .O(N__11590),
            .I(N__11587));
    CascadeMux I__961 (
            .O(N__11587),
            .I(N__11584));
    CascadeBuf I__960 (
            .O(N__11584),
            .I(N__11581));
    CascadeMux I__959 (
            .O(N__11581),
            .I(N__11578));
    CascadeBuf I__958 (
            .O(N__11578),
            .I(N__11575));
    CascadeMux I__957 (
            .O(N__11575),
            .I(N__11572));
    InMux I__956 (
            .O(N__11572),
            .I(N__11569));
    LocalMux I__955 (
            .O(N__11569),
            .I(N__11566));
    Span4Mux_h I__954 (
            .O(N__11566),
            .I(N__11563));
    Sp12to4 I__953 (
            .O(N__11563),
            .I(N__11560));
    Span12Mux_s3_v I__952 (
            .O(N__11560),
            .I(N__11557));
    Span12Mux_h I__951 (
            .O(N__11557),
            .I(N__11554));
    Odrv12 I__950 (
            .O(N__11554),
            .I(M_this_ppu_sprites_addr_8));
    CascadeMux I__949 (
            .O(N__11551),
            .I(N__11548));
    CascadeBuf I__948 (
            .O(N__11548),
            .I(N__11545));
    CascadeMux I__947 (
            .O(N__11545),
            .I(N__11542));
    CascadeBuf I__946 (
            .O(N__11542),
            .I(N__11539));
    CascadeMux I__945 (
            .O(N__11539),
            .I(N__11536));
    CascadeBuf I__944 (
            .O(N__11536),
            .I(N__11533));
    CascadeMux I__943 (
            .O(N__11533),
            .I(N__11530));
    CascadeBuf I__942 (
            .O(N__11530),
            .I(N__11527));
    CascadeMux I__941 (
            .O(N__11527),
            .I(N__11524));
    CascadeBuf I__940 (
            .O(N__11524),
            .I(N__11521));
    CascadeMux I__939 (
            .O(N__11521),
            .I(N__11518));
    CascadeBuf I__938 (
            .O(N__11518),
            .I(N__11515));
    CascadeMux I__937 (
            .O(N__11515),
            .I(N__11512));
    CascadeBuf I__936 (
            .O(N__11512),
            .I(N__11509));
    CascadeMux I__935 (
            .O(N__11509),
            .I(N__11506));
    CascadeBuf I__934 (
            .O(N__11506),
            .I(N__11503));
    CascadeMux I__933 (
            .O(N__11503),
            .I(N__11500));
    CascadeBuf I__932 (
            .O(N__11500),
            .I(N__11497));
    CascadeMux I__931 (
            .O(N__11497),
            .I(N__11494));
    CascadeBuf I__930 (
            .O(N__11494),
            .I(N__11491));
    CascadeMux I__929 (
            .O(N__11491),
            .I(N__11488));
    CascadeBuf I__928 (
            .O(N__11488),
            .I(N__11485));
    CascadeMux I__927 (
            .O(N__11485),
            .I(N__11482));
    CascadeBuf I__926 (
            .O(N__11482),
            .I(N__11479));
    CascadeMux I__925 (
            .O(N__11479),
            .I(N__11476));
    CascadeBuf I__924 (
            .O(N__11476),
            .I(N__11473));
    CascadeMux I__923 (
            .O(N__11473),
            .I(N__11470));
    CascadeBuf I__922 (
            .O(N__11470),
            .I(N__11467));
    CascadeMux I__921 (
            .O(N__11467),
            .I(N__11464));
    CascadeBuf I__920 (
            .O(N__11464),
            .I(N__11461));
    CascadeMux I__919 (
            .O(N__11461),
            .I(N__11458));
    InMux I__918 (
            .O(N__11458),
            .I(N__11455));
    LocalMux I__917 (
            .O(N__11455),
            .I(N__11452));
    Span4Mux_s2_v I__916 (
            .O(N__11452),
            .I(N__11449));
    Sp12to4 I__915 (
            .O(N__11449),
            .I(N__11446));
    Span12Mux_s6_h I__914 (
            .O(N__11446),
            .I(N__11443));
    Span12Mux_h I__913 (
            .O(N__11443),
            .I(N__11440));
    Odrv12 I__912 (
            .O(N__11440),
            .I(M_this_ppu_sprites_addr_7));
    CascadeMux I__911 (
            .O(N__11437),
            .I(N__11434));
    CascadeBuf I__910 (
            .O(N__11434),
            .I(N__11431));
    CascadeMux I__909 (
            .O(N__11431),
            .I(N__11428));
    CascadeBuf I__908 (
            .O(N__11428),
            .I(N__11425));
    CascadeMux I__907 (
            .O(N__11425),
            .I(N__11422));
    CascadeBuf I__906 (
            .O(N__11422),
            .I(N__11419));
    CascadeMux I__905 (
            .O(N__11419),
            .I(N__11416));
    CascadeBuf I__904 (
            .O(N__11416),
            .I(N__11413));
    CascadeMux I__903 (
            .O(N__11413),
            .I(N__11410));
    CascadeBuf I__902 (
            .O(N__11410),
            .I(N__11407));
    CascadeMux I__901 (
            .O(N__11407),
            .I(N__11404));
    CascadeBuf I__900 (
            .O(N__11404),
            .I(N__11401));
    CascadeMux I__899 (
            .O(N__11401),
            .I(N__11398));
    CascadeBuf I__898 (
            .O(N__11398),
            .I(N__11395));
    CascadeMux I__897 (
            .O(N__11395),
            .I(N__11392));
    CascadeBuf I__896 (
            .O(N__11392),
            .I(N__11389));
    CascadeMux I__895 (
            .O(N__11389),
            .I(N__11386));
    CascadeBuf I__894 (
            .O(N__11386),
            .I(N__11383));
    CascadeMux I__893 (
            .O(N__11383),
            .I(N__11380));
    CascadeBuf I__892 (
            .O(N__11380),
            .I(N__11377));
    CascadeMux I__891 (
            .O(N__11377),
            .I(N__11374));
    CascadeBuf I__890 (
            .O(N__11374),
            .I(N__11371));
    CascadeMux I__889 (
            .O(N__11371),
            .I(N__11368));
    CascadeBuf I__888 (
            .O(N__11368),
            .I(N__11365));
    CascadeMux I__887 (
            .O(N__11365),
            .I(N__11362));
    CascadeBuf I__886 (
            .O(N__11362),
            .I(N__11359));
    CascadeMux I__885 (
            .O(N__11359),
            .I(N__11356));
    CascadeBuf I__884 (
            .O(N__11356),
            .I(N__11353));
    CascadeMux I__883 (
            .O(N__11353),
            .I(N__11350));
    CascadeBuf I__882 (
            .O(N__11350),
            .I(N__11347));
    CascadeMux I__881 (
            .O(N__11347),
            .I(N__11344));
    InMux I__880 (
            .O(N__11344),
            .I(N__11341));
    LocalMux I__879 (
            .O(N__11341),
            .I(N__11338));
    Span4Mux_s2_v I__878 (
            .O(N__11338),
            .I(N__11335));
    Sp12to4 I__877 (
            .O(N__11335),
            .I(N__11332));
    Span12Mux_h I__876 (
            .O(N__11332),
            .I(N__11329));
    Odrv12 I__875 (
            .O(N__11329),
            .I(M_this_ppu_sprites_addr_6));
    CascadeMux I__874 (
            .O(N__11326),
            .I(N__11323));
    CascadeBuf I__873 (
            .O(N__11323),
            .I(N__11320));
    CascadeMux I__872 (
            .O(N__11320),
            .I(N__11317));
    CascadeBuf I__871 (
            .O(N__11317),
            .I(N__11314));
    CascadeMux I__870 (
            .O(N__11314),
            .I(N__11311));
    CascadeBuf I__869 (
            .O(N__11311),
            .I(N__11308));
    CascadeMux I__868 (
            .O(N__11308),
            .I(N__11305));
    CascadeBuf I__867 (
            .O(N__11305),
            .I(N__11302));
    CascadeMux I__866 (
            .O(N__11302),
            .I(N__11299));
    CascadeBuf I__865 (
            .O(N__11299),
            .I(N__11296));
    CascadeMux I__864 (
            .O(N__11296),
            .I(N__11293));
    CascadeBuf I__863 (
            .O(N__11293),
            .I(N__11290));
    CascadeMux I__862 (
            .O(N__11290),
            .I(N__11287));
    CascadeBuf I__861 (
            .O(N__11287),
            .I(N__11284));
    CascadeMux I__860 (
            .O(N__11284),
            .I(N__11281));
    CascadeBuf I__859 (
            .O(N__11281),
            .I(N__11278));
    CascadeMux I__858 (
            .O(N__11278),
            .I(N__11275));
    CascadeBuf I__857 (
            .O(N__11275),
            .I(N__11272));
    CascadeMux I__856 (
            .O(N__11272),
            .I(N__11269));
    CascadeBuf I__855 (
            .O(N__11269),
            .I(N__11266));
    CascadeMux I__854 (
            .O(N__11266),
            .I(N__11263));
    CascadeBuf I__853 (
            .O(N__11263),
            .I(N__11260));
    CascadeMux I__852 (
            .O(N__11260),
            .I(N__11257));
    CascadeBuf I__851 (
            .O(N__11257),
            .I(N__11254));
    CascadeMux I__850 (
            .O(N__11254),
            .I(N__11251));
    CascadeBuf I__849 (
            .O(N__11251),
            .I(N__11248));
    CascadeMux I__848 (
            .O(N__11248),
            .I(N__11245));
    CascadeBuf I__847 (
            .O(N__11245),
            .I(N__11242));
    CascadeMux I__846 (
            .O(N__11242),
            .I(N__11239));
    CascadeBuf I__845 (
            .O(N__11239),
            .I(N__11236));
    CascadeMux I__844 (
            .O(N__11236),
            .I(N__11233));
    InMux I__843 (
            .O(N__11233),
            .I(N__11230));
    LocalMux I__842 (
            .O(N__11230),
            .I(N__11227));
    Span4Mux_v I__841 (
            .O(N__11227),
            .I(N__11224));
    Span4Mux_h I__840 (
            .O(N__11224),
            .I(N__11221));
    Sp12to4 I__839 (
            .O(N__11221),
            .I(N__11218));
    Span12Mux_h I__838 (
            .O(N__11218),
            .I(N__11215));
    Odrv12 I__837 (
            .O(N__11215),
            .I(M_this_map_ram_read_data_4));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_23_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_17_0_));
    defparam IN_MUX_bfv_23_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_18_0_ (
            .carryinitin(M_this_data_count_q_cry_7),
            .carryinitout(bfn_23_18_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(un1_M_this_sprites_address_q_cry_7),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_19_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_22_0_));
    defparam IN_MUX_bfv_19_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_23_0_ (
            .carryinitin(un1_M_this_map_address_q_cry_7),
            .carryinitout(bfn_19_23_0_));
    defparam IN_MUX_bfv_22_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_20_0_));
    defparam IN_MUX_bfv_22_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_21_0_ (
            .carryinitin(un1_M_this_external_address_q_cry_7),
            .carryinitout(bfn_22_21_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNILD847_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__12091),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_614_1_g ));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNI0JBR6_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__12061),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_931_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_9  (
            .USERSIGNALTOGLOBALBUFFER(N__27493),
            .GLOBALBUFFEROUTPUT(M_this_reset_cond_out_g_0));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__21412),
            .GLOBALBUFFEROUTPUT(N_989_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOJ6UA_8_LC_2_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOJ6UA_8_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOJ6UA_8_LC_2_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIOJ6UA_8_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__17008),
            .in2(_gnd_net_),
            .in3(N__21642),
            .lcout(port_nmib_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_2_17_1 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_2_17_1 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_2_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11848),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32047),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_2_17_3 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_2_17_3 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_2_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11836),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32047),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_2_18_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_2_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_2_18_6  (
            .in0(N__13834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11902),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.port_data_rw_0_i_LC_2_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.port_data_rw_0_i_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.port_data_rw_0_i_LC_2_21_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_vga_signals.port_data_rw_0_i_LC_2_21_5  (
            .in0(N__25287),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21652),
            .lcout(port_data_rw_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_16_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_16_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_16_4  (
            .in0(N__13847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11931),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(N__15373),
            .in2(_gnd_net_),
            .in3(N__13825),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_19_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_19_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_19_3  (
            .in0(N__13848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15841),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_19_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_19_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_19_6  (
            .in0(N__13873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13849),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_0_LC_4_15_6 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_4_15_6 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_4_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11982),
            .lcout(\this_pixel_clk.M_counter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32028),
            .ce(),
            .sr(N__32393));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_4_16_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_4_16_0 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_4_16_0  (
            .in0(N__12163),
            .in1(N__27502),
            .in2(N__11932),
            .in3(N__15886),
            .lcout(\this_vga_ramdac.N_2870_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32037),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_17_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_17_1 .LUT_INIT=16'b0100011100100101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_17_1  (
            .in0(N__16868),
            .in1(N__16816),
            .in2(N__16678),
            .in3(N__16753),
            .lcout(\this_vga_ramdac.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_2  (
            .in0(N__15349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13846),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_4_18_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_4_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_4_18_3 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_4_18_3  (
            .in0(N__11908),
            .in1(N__27497),
            .in2(N__11901),
            .in3(N__15885),
            .lcout(\this_vga_ramdac.N_2875_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32045),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_2_LC_4_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_2_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_2_LC_4_19_0 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIADGD1_2_LC_4_19_0  (
            .in0(N__12040),
            .in1(N__13005),
            .in2(N__13225),
            .in3(N__12915),
            .lcout(),
            .ltout(\this_vga_signals.un4_hsynclto7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIF7AC4_8_LC_4_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIF7AC4_8_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIF7AC4_8_LC_4_19_1 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIF7AC4_8_LC_4_19_1  (
            .in0(N__13614),
            .in1(N__12031),
            .in2(N__11884),
            .in3(N__12834),
            .lcout(this_vga_signals_hsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNINT9T1_6_LC_4_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNINT9T1_6_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNINT9T1_6_LC_4_19_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNINT9T1_6_LC_4_19_3  (
            .in0(N__12916),
            .in1(N__12121),
            .in2(N__13009),
            .in3(N__12835),
            .lcout(),
            .ltout(\this_vga_signals.un2_hsynclt7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI73DH2_9_LC_4_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI73DH2_9_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI73DH2_9_LC_4_19_4 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI73DH2_9_LC_4_19_4  (
            .in0(N__13534),
            .in1(N__13613),
            .in2(N__12034),
            .in3(N__12726),
            .lcout(\this_vga_signals.hsync_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_4_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_4_20_0 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_4_20_0  (
            .in0(N__13533),
            .in1(N__13612),
            .in2(_gnd_net_),
            .in3(N__12725),
            .lcout(this_vga_signals_hvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_5_15_1 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_5_15_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_5_15_1  (
            .in0(N__11997),
            .in1(N__11983),
            .in2(_gnd_net_),
            .in3(N__32437),
            .lcout(\this_pixel_clk.M_counter_q_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32025),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_16_2 .LUT_INIT=16'b0010110110110100;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_16_2  (
            .in0(N__13000),
            .in1(N__13111),
            .in2(N__12324),
            .in3(N__14010),
            .lcout(),
            .ltout(\this_vga_signals.if_N_8_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_16_3 .LUT_INIT=16'b0011000011110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(N__13217),
            .in2(N__12004),
            .in3(N__13330),
            .lcout(\this_vga_signals.if_N_9_0_0 ),
            .ltout(\this_vga_signals.if_N_9_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_m2_LC_5_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_m2_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_m2_LC_5_16_4 .LUT_INIT=16'b0100011100011101;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_m2_LC_5_16_4  (
            .in0(N__13218),
            .in1(N__12213),
            .in2(N__12001),
            .in3(N__12073),
            .lcout(\this_vga_signals.mult1_un82_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_RNILQS8_1_LC_5_16_7 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_RNILQS8_1_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \this_pixel_clk.M_counter_q_RNILQS8_1_LC_5_16_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_pixel_clk.M_counter_q_RNILQS8_1_LC_5_16_7  (
            .in0(N__11998),
            .in1(N__11981),
            .in2(_gnd_net_),
            .in3(N__32427),
            .lcout(M_counter_q_RNILQS8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_3_LC_5_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_3_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_3_LC_5_17_0 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_3_LC_5_17_0  (
            .in0(N__12345),
            .in1(N__12448),
            .in2(_gnd_net_),
            .in3(N__12153),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_8_LC_5_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_8_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_8_LC_5_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_8_LC_5_17_1  (
            .in0(N__12115),
            .in1(N__12082),
            .in2(N__12094),
            .in3(N__14396),
            .lcout(\this_vga_signals.N_5_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILD847_9_LC_5_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILD847_9_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILD847_9_LC_5_17_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILD847_9_LC_5_17_2  (
            .in0(N__14636),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12051),
            .lcout(\this_vga_signals.N_614_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_5_LC_5_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_5_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_5_LC_5_17_3 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \this_vga_signals.un4_haddress_g0_5_LC_5_17_3  (
            .in0(N__12114),
            .in1(N__12914),
            .in2(_gnd_net_),
            .in3(N__12998),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_17_6 .LUT_INIT=16'b1001001111001001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_17_6  (
            .in0(N__12999),
            .in1(N__12313),
            .in2(N__13129),
            .in3(N__14011),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_x4_0_LC_5_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_x4_0_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_x4_0_LC_5_18_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_x4_0_LC_5_18_0  (
            .in0(N__12913),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13104),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_x4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_x4_2_LC_5_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_x4_2_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_x4_2_LC_5_18_1 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_x4_2_LC_5_18_1  (
            .in0(N__12833),
            .in1(N__12543),
            .in2(N__12076),
            .in3(N__12532),
            .lcout(\this_vga_signals.g0_i_x4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIST9Q2_9_LC_5_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIST9Q2_9_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIST9Q2_9_LC_5_18_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIST9Q2_9_LC_5_18_2  (
            .in0(N__14650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14475),
            .lcout(\this_vga_signals.N_931_1 ),
            .ltout(\this_vga_signals.N_931_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI0JBR6_9_LC_5_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI0JBR6_9_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI0JBR6_9_LC_5_18_3 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI0JBR6_9_LC_5_18_3  (
            .in0(N__14259),
            .in1(N__17433),
            .in2(N__12064),
            .in3(N__15999),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNI0JBR6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m5_i_a4_0_1_LC_5_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m5_i_a4_0_1_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m5_i_a4_0_1_LC_5_18_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_m5_i_a4_0_1_LC_5_18_5  (
            .in0(N__13106),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13329),
            .lcout(\this_vga_signals.un4_hsynclto3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_5_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_5_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_5_18_6  (
            .in0(N__13328),
            .in1(N__13222),
            .in2(N__13273),
            .in3(N__13105),
            .lcout(\this_vga_signals.un2_hsynclt6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_LC_5_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_LC_5_18_7 .LUT_INIT=16'b1111001010110000;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_LC_5_18_7  (
            .in0(N__12832),
            .in1(N__12912),
            .in2(N__12446),
            .in3(N__14304),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHO633_9_LC_5_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHO633_9_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHO633_9_LC_5_19_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIHO633_9_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__13415),
            .in2(_gnd_net_),
            .in3(N__14664),
            .lcout(\this_vga_signals.N_614_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_5_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_5_19_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_5_19_3  (
            .in0(N__12523),
            .in1(N__12262),
            .in2(_gnd_net_),
            .in3(N__12400),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_5_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_5_19_4 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_5_19_4  (
            .in0(N__12338),
            .in1(_gnd_net_),
            .in2(N__12106),
            .in3(N__12445),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_5_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_5_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_5_19_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_5_19_5  (
            .in0(N__13195),
            .in1(N__13234),
            .in2(N__13128),
            .in3(N__13004),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_d7lt7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI73DH2_0_9_LC_5_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI73DH2_0_9_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI73DH2_0_9_LC_5_19_6 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI73DH2_0_9_LC_5_19_6  (
            .in0(N__12100),
            .in1(N__13608),
            .in2(N__12103),
            .in3(N__13532),
            .lcout(\this_vga_signals.M_hcounter_d7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI11GM_7_LC_5_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI11GM_7_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI11GM_7_LC_5_19_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI11GM_7_LC_5_19_7  (
            .in0(N__12898),
            .in1(N__12721),
            .in2(_gnd_net_),
            .in3(N__12823),
            .lcout(\this_vga_signals.M_hcounter_d7lto7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_7_LC_5_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_7_LC_5_20_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_7_LC_5_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_7_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12685),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32048),
            .ce(N__13472),
            .sr(N__13431));
    defparam \this_vga_signals.M_hcounter_q_esr_8_LC_5_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_8_LC_5_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_8_LC_5_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_8_LC_5_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13570),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32048),
            .ce(N__13472),
            .sr(N__13431));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_8_LC_5_28_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_8_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_8_LC_5_28_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_8_LC_5_28_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17029),
            .lcout(this_vga_signals_vvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_4_LC_6_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_4_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_4_LC_6_15_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_4_LC_6_15_2  (
            .in0(N__12136),
            .in1(N__12320),
            .in2(N__12502),
            .in3(N__12214),
            .lcout(),
            .ltout(\this_vga_signals.g0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_7_LC_6_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_7_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_7_LC_6_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_7_LC_6_15_3  (
            .in0(N__12199),
            .in1(N__12658),
            .in2(N__12190),
            .in3(N__13384),
            .lcout(),
            .ltout(\this_vga_signals.g0_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIQFEIV5_9_LC_6_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIQFEIV5_9_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIQFEIV5_9_LC_6_15_4 .LUT_INIT=16'b0000101010000010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIQFEIV5_9_LC_6_15_4  (
            .in0(N__20963),
            .in1(N__12130),
            .in2(N__12187),
            .in3(N__13348),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_6_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_6_16_0 .LUT_INIT=16'b0010001010111011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_6_16_0  (
            .in0(N__13119),
            .in1(N__13207),
            .in2(_gnd_net_),
            .in3(N__12580),
            .lcout(\this_vga_signals.mult1_un75_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_16_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_16_2 .LUT_INIT=16'b0011001101000100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_16_2  (
            .in0(N__16815),
            .in1(N__16666),
            .in2(_gnd_net_),
            .in3(N__16751),
            .lcout(\this_vga_ramdac.N_24_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_LC_6_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_LC_6_16_4 .LUT_INIT=16'b0000001000101111;
    LogicCell40 \this_vga_signals.un4_haddress_g1_LC_6_16_4  (
            .in0(N__12253),
            .in1(N__12154),
            .in2(N__13130),
            .in3(N__13001),
            .lcout(\this_vga_signals.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIUAKU9_4_LC_6_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIUAKU9_4_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIUAKU9_4_LC_6_16_5 .LUT_INIT=16'b1101001001001011;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIUAKU9_4_LC_6_16_5  (
            .in0(N__13002),
            .in1(N__13118),
            .in2(N__12325),
            .in3(N__14013),
            .lcout(\this_vga_signals.M_hcounter_q_RNIUAKU9Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_0_LC_6_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_0_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_0_LC_6_17_0 .LUT_INIT=16'b1110010111011010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_0_LC_6_17_0  (
            .in0(N__13003),
            .in1(N__12572),
            .in2(N__13131),
            .in3(N__14012),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_3_0_0 ),
            .ltout(\this_vga_signals.mult1_un75_sum_ac0_3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1 .LUT_INIT=16'b0110011010010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1  (
            .in0(N__12573),
            .in1(N__12241),
            .in2(N__12256),
            .in3(N__13341),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g2_0_LC_6_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g2_0_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g2_0_LC_6_17_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.un4_haddress_g2_0_LC_6_17_2  (
            .in0(_gnd_net_),
            .in1(N__12447),
            .in2(_gnd_net_),
            .in3(N__12346),
            .lcout(\this_vga_signals.g2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_6_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_6_17_3 .LUT_INIT=16'b0000100101101111;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_6_17_3  (
            .in0(N__12575),
            .in1(N__13126),
            .in2(N__13223),
            .in3(N__12247),
            .lcout(\this_vga_signals.mult1_un82_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIB3UCP_1_LC_6_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIB3UCP_1_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIB3UCP_1_LC_6_17_4 .LUT_INIT=16'b1010010101011100;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIB3UCP_1_LC_6_17_4  (
            .in0(N__13317),
            .in1(N__13209),
            .in2(N__13132),
            .in3(N__12574),
            .lcout(\this_vga_signals.d_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIVPQGA_1_LC_6_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIVPQGA_1_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIVPQGA_1_LC_6_17_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIVPQGA_1_LC_6_17_6  (
            .in0(N__13318),
            .in1(N__13208),
            .in2(_gnd_net_),
            .in3(N__12240),
            .lcout(\this_vga_signals.d_N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_17_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_17_7 .LUT_INIT=16'b0110010100101011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_17_7  (
            .in0(N__16873),
            .in1(N__16814),
            .in2(N__16674),
            .in3(N__16747),
            .lcout(\this_vga_ramdac.m19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_1_LC_6_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_1_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_1_LC_6_18_0 .LUT_INIT=16'b1101001010110100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_1_LC_6_18_0  (
            .in0(N__12886),
            .in1(N__20912),
            .in2(N__13067),
            .in3(N__12971),
            .lcout(\this_vga_signals.mult1_un75_sum_axb2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_1 .LUT_INIT=16'b1111001010110000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_1  (
            .in0(N__12824),
            .in1(N__12883),
            .in2(N__12443),
            .in3(N__14302),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_6_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_6_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_6_18_2 .LUT_INIT=16'b0000101010101111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_6_18_2  (
            .in0(N__12885),
            .in1(_gnd_net_),
            .in2(N__12229),
            .in3(N__12972),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_6_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_6_18_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_6_18_3  (
            .in0(N__13110),
            .in1(N__14392),
            .in2(N__12226),
            .in3(N__14366),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_18_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_18_4  (
            .in0(N__14367),
            .in1(_gnd_net_),
            .in2(N__14400),
            .in3(N__14415),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_6_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_6_18_5 .LUT_INIT=16'b1100000110000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_6_18_5  (
            .in0(N__12825),
            .in1(N__12884),
            .in2(N__12444),
            .in3(N__14303),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_18_6 .LUT_INIT=16'b1100011111000001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_18_6  (
            .in0(N__13042),
            .in1(N__12970),
            .in2(N__12289),
            .in3(N__13994),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_LC_6_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_LC_6_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_LC_6_18_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_LC_6_18_7  (
            .in0(N__20913),
            .in1(N__12274),
            .in2(N__12286),
            .in3(N__12283),
            .lcout(\this_vga_signals.mult1_un75_sum_axb2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_6_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_6_19_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_6_19_0  (
            .in0(N__12719),
            .in1(N__12793),
            .in2(N__13626),
            .in3(N__13509),
            .lcout(\this_vga_signals.N_236 ),
            .ltout(\this_vga_signals.N_236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_6_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_6_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_6_19_1 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_6_19_1  (
            .in0(N__12880),
            .in1(N__12797),
            .in2(N__12277),
            .in3(N__12524),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_3_0 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_6_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_6_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_6_19_2  (
            .in0(_gnd_net_),
            .in1(N__20911),
            .in2(N__12268),
            .in3(N__13993),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIOIVT_6_LC_6_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIOIVT_6_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIOIVT_6_LC_6_19_3 .LUT_INIT=16'b1100011100011111;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNIOIVT_6_LC_6_19_3  (
            .in0(N__12364),
            .in1(N__13506),
            .in2(N__12388),
            .in3(N__12717),
            .lcout(\this_vga_signals.N_3_2_1 ),
            .ltout(\this_vga_signals.N_3_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_6_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_6_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_6_19_4 .LUT_INIT=16'b0010100011000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_6_19_4  (
            .in0(N__12950),
            .in1(N__12792),
            .in2(N__12265),
            .in3(N__12878),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_6_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_6_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_6_19_5 .LUT_INIT=16'b0101100101100101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_6_19_5  (
            .in0(N__12791),
            .in1(N__13507),
            .in2(N__13625),
            .in3(N__12718),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNIUFPQZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_6_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_6_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_6_19_6 .LUT_INIT=16'b0011101110000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_6_19_6  (
            .in0(N__12951),
            .in1(N__12879),
            .in2(N__12817),
            .in3(N__14301),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI43BG3_9_LC_6_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI43BG3_9_LC_6_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI43BG3_9_LC_6_19_7 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI43BG3_9_LC_6_19_7  (
            .in0(N__13618),
            .in1(N__13508),
            .in2(N__17018),
            .in3(N__12720),
            .lcout(M_this_vga_ramdac_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_8_LC_6_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_8_LC_6_20_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_8_LC_6_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_8_LC_6_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13563),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32046),
            .ce(N__13476),
            .sr(N__13436));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_7_LC_6_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_7_LC_6_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_7_LC_6_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_7_LC_6_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12678),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32046),
            .ce(N__13476),
            .sr(N__13436));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_9_LC_6_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_9_LC_6_20_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_9_LC_6_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_9_LC_6_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13546),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32046),
            .ce(N__13476),
            .sr(N__13436));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_6_LC_6_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_6_LC_6_20_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_6_LC_6_20_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_6_LC_6_20_3  (
            .in0(N__12742),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32046),
            .ce(N__13476),
            .sr(N__13436));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIIL511_7_LC_6_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIIL511_7_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIIL511_7_LC_6_20_4 .LUT_INIT=16'b0100110001001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNIIL511_7_LC_6_20_4  (
            .in0(N__12394),
            .in1(N__12387),
            .in2(N__12373),
            .in3(N__12363),
            .lcout(\this_vga_signals.SUM_3_i_0_0_3 ),
            .ltout(\this_vga_signals.SUM_3_i_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_20_5 .LUT_INIT=16'b0000100001011101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_20_5  (
            .in0(N__12881),
            .in1(N__12798),
            .in2(N__12349),
            .in3(N__12952),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_6_LC_6_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_6_LC_6_20_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_6_LC_6_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_6_LC_6_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12741),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32046),
            .ce(N__13476),
            .sr(N__13436));
    defparam \this_vga_signals.un4_haddress_g0_1_LC_6_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_1_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_1_LC_6_20_7 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_1_LC_6_20_7  (
            .in0(N__12882),
            .in1(N__12544),
            .in2(N__12826),
            .in3(N__12528),
            .lcout(\this_vga_signals.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJELD1_8_LC_7_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJELD1_8_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJELD1_8_LC_7_13_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIJELD1_8_LC_7_13_4  (
            .in0(N__15998),
            .in1(N__19230),
            .in2(N__18129),
            .in3(N__16494),
            .lcout(\this_vga_signals.vsync_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_7_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_7_15_0 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_7_15_0  (
            .in0(N__19233),
            .in1(N__18089),
            .in2(_gnd_net_),
            .in3(N__19701),
            .lcout(),
            .ltout(\this_vga_signals.un6_vvisibilitylt8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI81G42_7_LC_7_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI81G42_7_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI81G42_7_LC_7_15_1 .LUT_INIT=16'b0000110000010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI81G42_7_LC_7_15_1  (
            .in0(N__18090),
            .in1(N__16500),
            .in2(N__12487),
            .in3(N__16571),
            .lcout(),
            .ltout(\this_vga_signals.vvisibility_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_8_LC_7_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_8_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_8_LC_7_15_2 .LUT_INIT=16'b0001010100000101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_8_LC_7_15_2  (
            .in0(N__15997),
            .in1(N__16501),
            .in2(N__12484),
            .in3(N__14140),
            .lcout(this_vga_signals_vvisibility),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_7_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_7_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_7_16_0  (
            .in0(N__19708),
            .in1(N__16502),
            .in2(N__18128),
            .in3(N__16587),
            .lcout(\this_vga_signals.M_vcounter_d7lto8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_7_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_7_16_5 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_7_16_5  (
            .in0(N__17818),
            .in1(N__19246),
            .in2(N__19018),
            .in3(N__18550),
            .lcout(),
            .ltout(\this_vga_signals.vsync_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIUAQ3_7_LC_7_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIUAQ3_7_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIUAQ3_7_LC_7_16_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIUAQ3_7_LC_7_16_6  (
            .in0(N__19709),
            .in1(N__12481),
            .in2(N__12472),
            .in3(N__16588),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_7_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_7_17_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__13379),
            .in2(_gnd_net_),
            .in3(N__13360),
            .lcout(),
            .ltout(\this_vga_signals.if_m7_0_x4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_17_1 .LUT_INIT=16'b0111000100010111;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_17_1  (
            .in0(N__13315),
            .in1(N__13263),
            .in2(N__12664),
            .in3(N__12656),
            .lcout(),
            .ltout(\this_vga_signals.if_N_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_17_2 .LUT_INIT=16'b0010011100011011;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_17_2  (
            .in0(N__13914),
            .in1(N__13316),
            .in2(N__12661),
            .in3(N__13224),
            .lcout(\this_vga_signals.mult1_un89_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_17_3  (
            .in0(N__13380),
            .in1(N__12657),
            .in2(N__12643),
            .in3(N__13913),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI32C8PD_9_LC_7_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI32C8PD_9_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI32C8PD_9_LC_7_17_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI32C8PD_9_LC_7_17_4  (
            .in0(N__20962),
            .in1(N__12586),
            .in2(N__12634),
            .in3(N__12631),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_17_5 .LUT_INIT=16'b0000111101000100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_17_5  (
            .in0(N__12610),
            .in1(N__12604),
            .in2(N__12598),
            .in3(N__12550),
            .lcout(\this_vga_signals.mult1_un89_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m5_i_LC_7_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m5_i_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m5_i_LC_7_17_7 .LUT_INIT=16'b0100011001100010;
    LogicCell40 \this_vga_signals.un4_haddress_if_m5_i_LC_7_17_7  (
            .in0(N__13314),
            .in1(N__13213),
            .in2(N__13127),
            .in3(N__12579),
            .lcout(\this_vga_signals.N_2_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_7_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_7_18_1 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(N__13264),
            .in2(N__14718),
            .in3(N__13319),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32029),
            .ce(),
            .sr(N__13432));
    defparam \this_vga_signals.M_hcounter_q_0_LC_7_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_7_18_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_7_18_2  (
            .in0(N__13265),
            .in1(N__14706),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32029),
            .ce(),
            .sr(N__13432));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_d_LC_7_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_d_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_d_LC_7_18_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_d_LC_7_18_7  (
            .in0(N__13177),
            .in1(N__13378),
            .in2(_gnd_net_),
            .in3(N__13359),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_3_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_7_19_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_7_19_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_7_19_0  (
            .in0(N__13259),
            .in1(N__13310),
            .in2(N__13269),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_d7lt4 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_7_19_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_7_19_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_7_19_1  (
            .in0(N__14691),
            .in1(N__13194),
            .in2(_gnd_net_),
            .in3(N__13135),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__32038),
            .ce(),
            .sr(N__13443));
    defparam \this_vga_signals.M_hcounter_q_3_LC_7_19_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_7_19_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_7_19_2  (
            .in0(N__14689),
            .in1(N__13066),
            .in2(_gnd_net_),
            .in3(N__13012),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__32038),
            .ce(),
            .sr(N__13443));
    defparam \this_vga_signals.M_hcounter_q_4_LC_7_19_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_7_19_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_7_19_3  (
            .in0(N__14692),
            .in1(N__12997),
            .in2(_gnd_net_),
            .in3(N__12919),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__32038),
            .ce(),
            .sr(N__13443));
    defparam \this_vga_signals.M_hcounter_q_5_LC_7_19_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_7_19_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_7_19_4  (
            .in0(N__14690),
            .in1(N__12897),
            .in2(_gnd_net_),
            .in3(N__12838),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__32038),
            .ce(),
            .sr(N__13443));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_7_19_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_7_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__12813),
            .in2(_gnd_net_),
            .in3(N__12733),
            .lcout(\this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_7_19_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_7_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__12730),
            .in2(_gnd_net_),
            .in3(N__12667),
            .lcout(\this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_7_19_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_7_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__13627),
            .in2(_gnd_net_),
            .in3(N__13552),
            .lcout(\this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_7_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_7_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__13525),
            .in2(_gnd_net_),
            .in3(N__13549),
            .lcout(\this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_7_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_7_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_7_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13545),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32041),
            .ce(N__13477),
            .sr(N__13444));
    defparam \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_9_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_9_12_2 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_9_12_2  (
            .in0(N__17305),
            .in1(N__15072),
            .in2(_gnd_net_),
            .in3(N__15325),
            .lcout(\this_vga_signals.g0_31_N_4L6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_3_LC_9_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_3_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_3_LC_9_12_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_3_LC_9_12_3  (
            .in0(N__19475),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17306),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_9_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_9_12_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_11_LC_9_12_4  (
            .in0(N__19750),
            .in1(N__16140),
            .in2(N__13387),
            .in3(N__17225),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_9_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_9_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__14998),
            .in2(_gnd_net_),
            .in3(N__14968),
            .lcout(\this_vga_signals.vaddress_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_9_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_9_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14788),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31980),
            .ce(N__15140),
            .sr(N__15114));
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_9_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_9_13_3 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_34_LC_9_13_3  (
            .in0(N__16578),
            .in1(N__15081),
            .in2(N__16504),
            .in3(N__15960),
            .lcout(),
            .ltout(\this_vga_signals.if_m8_0_a3_1_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_9_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_9_13_4 .LUT_INIT=16'b0010111000011101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_9_13_4  (
            .in0(N__13657),
            .in1(N__13648),
            .in2(N__13651),
            .in3(N__17179),
            .lcout(\this_vga_signals.g0_31_N_5L8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_31_N_3L3_LC_9_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_3L3_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_3L3_LC_9_13_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_N_3L3_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__19615),
            .in2(_gnd_net_),
            .in3(N__19474),
            .lcout(\this_vga_signals.g0_31_N_3L3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_9_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_9_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14787),
            .lcout(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31980),
            .ce(N__15140),
            .sr(N__15114));
    defparam \this_vga_signals.un5_vaddress_g3_3_0_LC_9_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_3_0_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_3_0_LC_9_14_0 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_3_0_LC_9_14_0  (
            .in0(N__18042),
            .in1(N__19617),
            .in2(_gnd_net_),
            .in3(N__19458),
            .lcout(\this_vga_signals.g3_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_9_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_9_14_1 .LUT_INIT=16'b0110110110110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_32_LC_9_14_1  (
            .in0(N__16498),
            .in1(N__16585),
            .in2(N__18115),
            .in3(N__15975),
            .lcout(),
            .ltout(\this_vga_signals.if_m8_0_a3_1_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_8_0_LC_9_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_8_0_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_8_0_LC_9_14_2 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_8_0_LC_9_14_2  (
            .in0(N__13761),
            .in1(N__13642),
            .in2(N__13636),
            .in3(N__17211),
            .lcout(),
            .ltout(\this_vga_signals.g0_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_9_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_9_14_3 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_27_LC_9_14_3  (
            .in0(N__19131),
            .in1(N__17675),
            .in2(N__13633),
            .in3(N__18394),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_9_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_9_14_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__19616),
            .in2(_gnd_net_),
            .in3(N__19462),
            .lcout(\this_vga_signals.vaddress_2_5 ),
            .ltout(\this_vga_signals.vaddress_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_9_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_9_14_5 .LUT_INIT=16'b0110000101001001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_LC_9_14_5  (
            .in0(N__17943),
            .in1(N__17224),
            .in2(N__13630),
            .in3(N__16054),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_9_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_9_14_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__17303),
            .in2(_gnd_net_),
            .in3(N__15322),
            .lcout(\this_vga_signals.g1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_9_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_9_14_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_9_14_7  (
            .in0(N__17304),
            .in1(_gnd_net_),
            .in2(N__19508),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.vaddress_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_9_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_9_15_0 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_19_LC_9_15_0  (
            .in0(N__15990),
            .in1(N__16469),
            .in2(N__18083),
            .in3(N__16570),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_9_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_9_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14812),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31992),
            .ce(N__15138),
            .sr(N__15115));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_9_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_9_15_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_9_15_2  (
            .in0(N__14839),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31992),
            .ce(N__15138),
            .sr(N__15115));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_9_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_9_15_3 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_9_15_3  (
            .in0(N__18031),
            .in1(N__19463),
            .in2(_gnd_net_),
            .in3(N__17331),
            .lcout(\this_vga_signals.vaddress_3_0_6 ),
            .ltout(\this_vga_signals.vaddress_3_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_33_LC_9_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_33_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_33_LC_9_15_4 .LUT_INIT=16'b1100111111110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_33_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__17204),
            .in2(N__13669),
            .in3(N__17942),
            .lcout(),
            .ltout(\this_vga_signals.g2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_1_LC_9_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_1_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_1_LC_9_15_5 .LUT_INIT=16'b0001110111001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_1_LC_9_15_5  (
            .in0(N__18395),
            .in1(N__19228),
            .in2(N__13666),
            .in3(N__19643),
            .lcout(\this_vga_signals.g1_1_1 ),
            .ltout(\this_vga_signals.g1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_2_LC_9_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_2_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_2_LC_9_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_2_LC_9_15_6  (
            .in0(N__13750),
            .in1(N__18231),
            .in2(N__13663),
            .in3(N__18396),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_x4_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_9_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_9_15_7 .LUT_INIT=16'b0100101100101101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_9_15_7  (
            .in0(N__19229),
            .in1(N__18991),
            .in2(N__13660),
            .in3(N__14182),
            .lcout(\this_vga_signals.g0_i_x4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_9_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_9_16_2 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_LC_9_16_2  (
            .in0(N__18026),
            .in1(N__19641),
            .in2(_gnd_net_),
            .in3(N__19455),
            .lcout(\this_vga_signals.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_9_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_9_16_3 .LUT_INIT=16'b0010010010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_28_LC_9_16_3  (
            .in0(N__13765),
            .in1(N__17219),
            .in2(N__13744),
            .in3(N__17940),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_9_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_9_16_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__19642),
            .in2(_gnd_net_),
            .in3(N__19457),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_9_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_9_16_5 .LUT_INIT=16'b0010010011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_36_LC_9_16_5  (
            .in0(N__13743),
            .in1(N__17218),
            .in2(N__13729),
            .in3(N__17941),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i_1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_1_LC_9_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_1_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_1_LC_9_16_6 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_1_LC_9_16_6  (
            .in0(N__18027),
            .in1(N__19456),
            .in2(_gnd_net_),
            .in3(N__17330),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_3_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_9_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_9_16_7 .LUT_INIT=16'b0100010101010000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_22_LC_9_16_7  (
            .in0(N__16198),
            .in1(N__17217),
            .in2(N__13726),
            .in3(N__17939),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_9_17_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_9_17_0 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_9_17_0  (
            .in0(N__23196),
            .in1(N__13675),
            .in2(N__14059),
            .in3(N__29674),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_9_17_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_9_17_1 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_9_17_1  (
            .in0(N__14023),
            .in1(N__23197),
            .in2(N__13723),
            .in3(N__13771),
            .lcout(M_this_ppu_vram_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_9_17_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_9_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_9_17_2  (
            .in0(N__27804),
            .in1(N__13702),
            .in2(_gnd_net_),
            .in3(N__13687),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_9_17_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_9_17_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_9_17_3  (
            .in0(N__27801),
            .in1(N__14086),
            .in2(_gnd_net_),
            .in3(N__14077),
            .lcout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_9_17_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_9_17_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_9_17_4  (
            .in0(N__14050),
            .in1(N__14038),
            .in2(_gnd_net_),
            .in3(N__27802),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIL26KA_9_LC_9_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIL26KA_9_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIL26KA_9_LC_9_17_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIL26KA_9_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__20982),
            .in2(_gnd_net_),
            .in3(N__14017),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_9_17_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_9_17_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_9_17_6  (
            .in0(N__13948),
            .in1(N__13930),
            .in2(_gnd_net_),
            .in3(N__27803),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC813H3_9_LC_9_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC813H3_9_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC813H3_9_LC_9_17_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIC813H3_9_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__20981),
            .in2(_gnd_net_),
            .in3(N__13918),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_0 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_0  (
            .in0(N__13885),
            .in1(N__27489),
            .in2(N__13866),
            .in3(N__15874),
            .lcout(\this_vga_ramdac.N_2874_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32015),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_18_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_18_4 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_ret_LC_9_18_4  (
            .in0(N__20999),
            .in1(N__13813),
            .in2(N__27501),
            .in3(N__15875),
            .lcout(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32015),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_9_18_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_9_18_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_9_18_7  (
            .in0(N__13798),
            .in1(N__13780),
            .in2(_gnd_net_),
            .in3(N__27805),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_10_11_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_10_11_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_10_11_0  (
            .in0(N__14693),
            .in1(N__18572),
            .in2(N__14536),
            .in3(N__14535),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__31954),
            .ce(),
            .sr(N__15108));
    defparam \this_vga_signals.M_vcounter_q_1_LC_10_11_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_10_11_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_10_11_1  (
            .in0(N__14714),
            .in1(N__18513),
            .in2(_gnd_net_),
            .in3(N__14113),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__31954),
            .ce(),
            .sr(N__15108));
    defparam \this_vga_signals.M_vcounter_q_2_LC_10_11_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_10_11_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_10_11_2  (
            .in0(N__14694),
            .in1(N__17789),
            .in2(_gnd_net_),
            .in3(N__14110),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__31954),
            .ce(),
            .sr(N__15108));
    defparam \this_vga_signals.M_vcounter_q_3_LC_10_11_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_10_11_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_10_11_3  (
            .in0(N__14715),
            .in1(N__18913),
            .in2(_gnd_net_),
            .in3(N__14107),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__31954),
            .ce(),
            .sr(N__15108));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_11_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__19203),
            .in2(_gnd_net_),
            .in3(N__14104),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_11_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__19700),
            .in2(_gnd_net_),
            .in3(N__14101),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_11_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__18105),
            .in2(_gnd_net_),
            .in3(N__14098),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_11_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__16584),
            .in2(_gnd_net_),
            .in3(N__14095),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_12_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__16499),
            .in2(_gnd_net_),
            .in3(N__14092),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_10_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_10_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__15964),
            .in2(_gnd_net_),
            .in3(N__14089),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31962),
            .ce(N__15142),
            .sr(N__15110));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_10_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_10_13_0 .LUT_INIT=16'b0000101100011101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_10_13_0  (
            .in0(N__14939),
            .in1(N__15938),
            .in2(N__14758),
            .in3(N__14891),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_13_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__15158),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31967),
            .ce(N__15141),
            .sr(N__15112));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_13_2  (
            .in0(N__15159),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31967),
            .ce(N__15141),
            .sr(N__15112));
    defparam \this_vga_signals.un5_vaddress_g1_1_0_LC_10_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_0_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_0_LC_10_13_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_0_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__19130),
            .in2(_gnd_net_),
            .in3(N__18362),
            .lcout(this_vga_signals_un5_vaddress_g1_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_10_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_10_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14834),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31967),
            .ce(N__15141),
            .sr(N__15112));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_13_7  (
            .in0(N__14835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31967),
            .ce(N__15141),
            .sr(N__15112));
    defparam \this_vga_signals.un5_vaddress_g2_3_LC_10_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_3_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_3_LC_10_14_0 .LUT_INIT=16'b0110111111111001;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_3_LC_10_14_0  (
            .in0(N__17199),
            .in1(N__18038),
            .in2(N__19231),
            .in3(N__19663),
            .lcout(\this_vga_signals.g2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_10_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_10_14_1 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_10_14_1  (
            .in0(N__14940),
            .in1(N__14892),
            .in2(N__15076),
            .in3(N__15965),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_10_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_10_14_2 .LUT_INIT=16'b1110011100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_10_14_2  (
            .in0(N__14136),
            .in1(N__15064),
            .in2(N__14122),
            .in3(N__14119),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_LC_10_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_LC_10_14_3 .LUT_INIT=16'b1011100111100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_LC_10_14_3  (
            .in0(N__17887),
            .in1(N__18084),
            .in2(N__14176),
            .in3(N__14173),
            .lcout(\this_vga_signals.g2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_LC_10_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_LC_10_14_4 .LUT_INIT=16'b0010110110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_LC_10_14_4  (
            .in0(N__16138),
            .in1(N__16166),
            .in2(N__19512),
            .in3(N__17883),
            .lcout(\this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJHZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_0_LC_10_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_0_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_0_LC_10_14_5 .LUT_INIT=16'b0011100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5_0_LC_10_14_5  (
            .in0(N__16167),
            .in1(N__19470),
            .in2(N__17917),
            .in3(N__16139),
            .lcout(\this_vga_signals.M_vcounter_q_4_rep2_esr_RNIBUJH5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_10_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_10_14_6 .LUT_INIT=16'b0011001000110011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_LC_10_14_6  (
            .in0(N__17679),
            .in1(N__14164),
            .in2(N__19232),
            .in3(N__18372),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_10_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_10_14_7 .LUT_INIT=16'b0111111011100111;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_0_LC_10_14_7  (
            .in0(N__19664),
            .in1(N__19471),
            .in2(N__18088),
            .in3(N__17200),
            .lcout(\this_vga_signals.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_10_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_10_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_20_LC_10_15_0  (
            .in0(N__17673),
            .in1(N__15265),
            .in2(N__14158),
            .in3(N__18232),
            .lcout(\this_vga_signals.N_4_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_LC_10_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_LC_10_15_1 .LUT_INIT=16'b0101001101001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_LC_10_15_1  (
            .in0(N__17177),
            .in1(N__19644),
            .in2(N__18100),
            .in3(N__19507),
            .lcout(\this_vga_signals.g2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICU8TI_6_LC_10_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICU8TI_6_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICU8TI_6_LC_10_15_2 .LUT_INIT=16'b0011011001100011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICU8TI_6_LC_10_15_2  (
            .in0(N__17920),
            .in1(N__16280),
            .in2(N__18127),
            .in3(N__18141),
            .lcout(),
            .ltout(\this_vga_signals.m9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVKPDR_5_LC_10_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVKPDR_5_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVKPDR_5_LC_10_15_3 .LUT_INIT=16'b1001011010100101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIVKPDR_5_LC_10_15_3  (
            .in0(N__19703),
            .in1(N__18156),
            .in2(N__14149),
            .in3(N__17921),
            .lcout(\this_vga_signals.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_10_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_10_15_4 .LUT_INIT=16'b0001110011011101;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_3_LC_10_15_4  (
            .in0(N__18361),
            .in1(N__19202),
            .in2(N__19692),
            .in3(N__14146),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_10_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_10_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_30_LC_10_15_5  (
            .in0(N__18960),
            .in1(N__14227),
            .in2(N__14221),
            .in3(N__17672),
            .lcout(\this_vga_signals.g0_1_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_2_LC_10_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_2_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_2_LC_10_15_6 .LUT_INIT=16'b1110111001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_2_LC_10_15_6  (
            .in0(N__17919),
            .in1(N__14215),
            .in2(_gnd_net_),
            .in3(N__17178),
            .lcout(),
            .ltout(\this_vga_signals.g2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_10_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_10_15_7 .LUT_INIT=16'b0001101110101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_0_LC_10_15_7  (
            .in0(N__19201),
            .in1(N__18360),
            .in2(N__14218),
            .in3(N__19648),
            .lcout(\this_vga_signals.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_10_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_10_16_0 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_10_16_0  (
            .in0(N__17335),
            .in1(N__15077),
            .in2(_gnd_net_),
            .in3(N__15323),
            .lcout(\this_vga_signals.vaddress_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_10_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_10_16_1 .LUT_INIT=16'b1010100000100010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_LC_10_16_1  (
            .in0(N__15244),
            .in1(N__14209),
            .in2(N__19004),
            .in3(N__15214),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_10_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_10_16_2 .LUT_INIT=16'b1101010001001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_LC_10_16_2  (
            .in0(N__18526),
            .in1(N__17813),
            .in2(N__14203),
            .in3(N__14200),
            .lcout(\this_vga_signals.if_i1_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_10_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_10_16_3 .LUT_INIT=16'b0111100010000111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_5_LC_10_16_3  (
            .in0(N__15324),
            .in1(N__17337),
            .in2(N__15082),
            .in3(N__17220),
            .lcout(),
            .ltout(\this_vga_signals.g1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_10_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_10_16_4 .LUT_INIT=16'b1110001010111000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_29_LC_10_16_4  (
            .in0(N__15199),
            .in1(N__19241),
            .in2(N__14194),
            .in3(N__19702),
            .lcout(),
            .ltout(\this_vga_signals.g0_2_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_10_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_10_16_5 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_35_LC_10_16_5  (
            .in0(N__19242),
            .in1(N__14191),
            .in2(N__14185),
            .in3(N__18397),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_10_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_10_16_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_10_16_6  (
            .in0(N__17336),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19472),
            .lcout(\this_vga_signals.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIT8RA8_LC_10_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIT8RA8_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIT8RA8_LC_10_16_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIT8RA8_LC_10_16_7  (
            .in0(N__19473),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17680),
            .lcout(\this_vga_signals.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNICEV1S_9_LC_10_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICEV1S_9_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICEV1S_9_LC_10_17_1 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNICEV1S_9_LC_10_17_1  (
            .in0(N__14422),
            .in1(N__14404),
            .in2(N__21001),
            .in3(N__14374),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_10_17_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_10_17_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_sprites_ram.mem_mem_4_0_wclke_3_LC_10_17_2  (
            .in0(N__20801),
            .in1(N__25732),
            .in2(N__23348),
            .in3(N__24577),
            .lcout(\this_sprites_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNISLAE4_6_LC_10_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNISLAE4_6_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNISLAE4_6_LC_10_17_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNISLAE4_6_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__20998),
            .in2(_gnd_net_),
            .in3(N__14311),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_0_LC_10_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_0_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_0_LC_10_17_7 .LUT_INIT=16'b0110010011001100;
    LogicCell40 \this_vga_signals.M_lcounter_q_0_LC_10_17_7  (
            .in0(N__14716),
            .in1(N__16018),
            .in2(N__14239),
            .in3(N__14531),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31994),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_e_0_RNIR1JA4_1_LC_10_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_e_0_RNIR1JA4_1_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_e_0_RNIR1JA4_1_LC_10_18_0 .LUT_INIT=16'b0010000000110011;
    LogicCell40 \this_vga_signals.M_lcounter_q_e_0_RNIR1JA4_1_LC_10_18_0  (
            .in0(N__17434),
            .in1(N__16032),
            .in2(N__14263),
            .in3(N__15994),
            .lcout(\this_vga_signals.M_lcounter_d_0_sqmuxa ),
            .ltout(\this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_e_0_1_LC_10_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_e_0_1_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_e_0_1_LC_10_18_1 .LUT_INIT=16'b0110000010101010;
    LogicCell40 \this_vga_signals.M_lcounter_q_e_0_1_LC_10_18_1  (
            .in0(N__16033),
            .in1(N__16017),
            .in2(N__14230),
            .in3(N__14528),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32002),
            .ce(N__14717),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_10_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_10_18_3 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_1_LC_10_18_3  (
            .in0(N__14566),
            .in1(N__14737),
            .in2(N__14590),
            .in3(N__14530),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32002),
            .ce(N__14717),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_10_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_10_18_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_0_LC_10_18_6  (
            .in0(N__14529),
            .in1(N__14548),
            .in2(_gnd_net_),
            .in3(N__14565),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32002),
            .ce(N__14717),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIOB8H3_0_LC_10_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIOB8H3_0_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIOB8H3_0_LC_10_19_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNIOB8H3_0_LC_10_19_0  (
            .in0(N__14736),
            .in1(_gnd_net_),
            .in2(N__14719),
            .in3(N__14452),
            .lcout(N_2_0),
            .ltout(N_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_10_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_10_19_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14740),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_pcounter_q_i_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32007),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_RNI5JMN3_LC_10_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_RNI5JMN3_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_RNI5JMN3_LC_10_19_2 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_RNI5JMN3_LC_10_19_2  (
            .in0(N__14505),
            .in1(N__14735),
            .in2(N__14589),
            .in3(N__14564),
            .lcout(),
            .ltout(\this_vga_signals.M_pcounter_q_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNILGGG4_1_LC_10_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNILGGG4_1_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNILGGG4_1_LC_10_19_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNILGGG4_1_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__14710),
            .in2(N__14593),
            .in3(N__14585),
            .lcout(N_3_0),
            .ltout(N_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_LC_10_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_10_19_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14569),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_pcounter_q_i_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32007),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNI9FEO2_LC_10_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNI9FEO2_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNI9FEO2_LC_10_19_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_RNI9FEO2_LC_10_19_7  (
            .in0(N__14563),
            .in1(N__14547),
            .in2(_gnd_net_),
            .in3(N__14504),
            .lcout(\this_vga_signals.M_pcounter_q_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_10_20_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_10_20_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_5_0_wclke_3_LC_10_20_1  (
            .in0(N__25728),
            .in1(N__24568),
            .in2(N__23347),
            .in3(N__20809),
            .lcout(\this_sprites_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14804),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31950),
            .ce(N__15145),
            .sr(N__15107));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_12_2 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_12_2  (
            .in0(N__15039),
            .in1(N__17342),
            .in2(_gnd_net_),
            .in3(N__15291),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14833),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31955),
            .ce(N__15144),
            .sr(N__15109));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_11_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_11_12_4 .LUT_INIT=16'b1111100000000111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_11_12_4  (
            .in0(N__14993),
            .in1(N__15290),
            .in2(N__15060),
            .in3(N__14890),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_11_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_11_12_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_11_12_5  (
            .in0(N__14805),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31955),
            .ce(N__15144),
            .sr(N__15109));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14778),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31955),
            .ce(N__15144),
            .sr(N__15109));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_12_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_12_7  (
            .in0(N__14909),
            .in1(N__14994),
            .in2(N__14767),
            .in3(N__14967),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_11_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_11_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15183),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31963),
            .ce(N__15143),
            .sr(N__15111));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_11_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_11_13_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_11_13_1  (
            .in0(N__14992),
            .in1(N__14966),
            .in2(_gnd_net_),
            .in3(N__14749),
            .lcout(),
            .ltout(\this_vga_signals.N_1_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_11_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_11_13_2 .LUT_INIT=16'b1010111111101111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_11_13_2  (
            .in0(N__14911),
            .in1(N__14938),
            .in2(N__14743),
            .in3(N__15937),
            .lcout(),
            .ltout(\this_vga_signals.SUM_2_i_1_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_11_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_11_13_3 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_11_13_3  (
            .in0(N__15007),
            .in1(N__14863),
            .in2(N__15001),
            .in3(N__14947),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_11_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_11_13_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_11_13_4  (
            .in0(N__15935),
            .in1(N__14991),
            .in2(N__14941),
            .in3(N__14886),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_11_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_11_13_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14971),
            .in3(N__14965),
            .lcout(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15182),
            .lcout(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31963),
            .ce(N__15143),
            .sr(N__15111));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_13_7 .LUT_INIT=16'b1010101001111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_13_7  (
            .in0(N__14937),
            .in1(N__14910),
            .in2(N__14893),
            .in3(N__15936),
            .lcout(\this_vga_signals.SUM_2_i_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_11_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_11_14_0 .LUT_INIT=16'b0010010011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m2_1_LC_11_14_0  (
            .in0(N__17171),
            .in1(N__16136),
            .in2(N__16178),
            .in3(N__17901),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI87FSD_LC_11_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI87FSD_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI87FSD_LC_11_14_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI87FSD_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__17170),
            .in2(N__14857),
            .in3(N__14848),
            .lcout(\this_vga_signals.d_N_3_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_14_2 .LUT_INIT=16'b0100001010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_14_2  (
            .in0(N__17172),
            .in1(N__16137),
            .in2(N__16179),
            .in3(N__17902),
            .lcout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i),
            .ltout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam m18x_N_3L3_LC_11_14_3.C_ON=1'b0;
    defparam m18x_N_3L3_LC_11_14_3.SEQ_MODE=4'b0000;
    defparam m18x_N_3L3_LC_11_14_3.LUT_INIT=16'b0011011111001000;
    LogicCell40 m18x_N_3L3_LC_11_14_3 (
            .in0(N__16950),
            .in1(N__17593),
            .in2(N__14842),
            .in3(N__18267),
            .lcout(m18x_N_3LZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_11_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_11_14_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_15_LC_11_14_4  (
            .in0(N__17174),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18116),
            .lcout(\this_vga_signals.N_5_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM43JE1_5_LC_11_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM43JE1_5_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM43JE1_5_LC_11_14_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIM43JE1_5_LC_11_14_5  (
            .in0(N__15208),
            .in1(N__17467),
            .in2(N__16069),
            .in3(N__17594),
            .lcout(\this_vga_signals.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_1_LC_11_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_1_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_1_LC_11_14_6 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_1_LC_11_14_6  (
            .in0(N__17344),
            .in1(N__15066),
            .in2(_gnd_net_),
            .in3(N__15310),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_11_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_11_14_7 .LUT_INIT=16'b1111101001011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_1_LC_11_14_7  (
            .in0(N__17903),
            .in1(_gnd_net_),
            .in2(N__15202),
            .in3(N__17173),
            .lcout(\this_vga_signals.g2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_37_LC_11_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_37_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_37_LC_11_15_0 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_37_LC_11_15_0  (
            .in0(N__15996),
            .in1(N__16442),
            .in2(N__18123),
            .in3(N__16539),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_11_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_11_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15187),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31972),
            .ce(N__15139),
            .sr(N__15113));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_11_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_11_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15166),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31972),
            .ce(N__15139),
            .sr(N__15113));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_11_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_11_15_3 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_11_15_3  (
            .in0(N__16538),
            .in1(N__15065),
            .in2(N__16468),
            .in3(N__15995),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_1 ),
            .ltout(\this_vga_signals.if_m8_0_a3_1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_15_4 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__17341),
            .in2(N__15010),
            .in3(N__15309),
            .lcout(),
            .ltout(\this_vga_signals.if_N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_11_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_11_15_5 .LUT_INIT=16'b0000110100001110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_LC_11_15_5  (
            .in0(N__16134),
            .in1(N__16168),
            .in2(N__15328),
            .in3(N__17175),
            .lcout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_11_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_11_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__17340),
            .in2(_gnd_net_),
            .in3(N__15308),
            .lcout(\this_vga_signals.vaddress_5 ),
            .ltout(\this_vga_signals.vaddress_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_11_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_11_15_7 .LUT_INIT=16'b0000110100001010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_11_15_7  (
            .in0(N__16135),
            .in1(N__17176),
            .in2(N__15268),
            .in3(N__17918),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_11_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_11_16_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_2_LC_11_16_0  (
            .in0(N__18996),
            .in1(N__15264),
            .in2(N__19257),
            .in3(N__17678),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_11_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_11_16_1 .LUT_INIT=16'b1111110101111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_26_LC_11_16_1  (
            .in0(N__17812),
            .in1(N__15253),
            .in2(N__15247),
            .in3(N__18228),
            .lcout(\this_vga_signals.g1_0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIB3A8M_LC_11_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIB3A8M_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIB3A8M_LC_11_16_2 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIB3A8M_LC_11_16_2  (
            .in0(N__15238),
            .in1(N__16347),
            .in2(N__19360),
            .in3(N__18391),
            .lcout(\this_vga_signals.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_LC_11_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_LC_11_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x2_LC_11_16_3  (
            .in0(N__15229),
            .in1(N__16288),
            .in2(_gnd_net_),
            .in3(N__18229),
            .lcout(\this_vga_signals.N_5_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_2_x1_LC_11_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_2_x1_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_2_x1_LC_11_16_4 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_2_x1_LC_11_16_4  (
            .in0(N__16310),
            .in1(N__19237),
            .in2(N__19013),
            .in3(N__17676),
            .lcout(\this_vga_signals.g0_2_0_2_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_2_x0_LC_11_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_2_x0_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_2_x0_LC_11_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_2_x0_LC_11_16_5  (
            .in0(N__17677),
            .in1(N__18995),
            .in2(N__19255),
            .in3(N__16309),
            .lcout(),
            .ltout(\this_vga_signals.g0_2_0_2_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_2_ns_LC_11_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_2_ns_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_2_ns_LC_11_16_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_2_ns_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__15481),
            .in2(N__15475),
            .in3(N__18390),
            .lcout(\this_vga_signals.g0_2_0_2 ),
            .ltout(\this_vga_signals.g0_2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_11_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_11_16_7 .LUT_INIT=16'b1101111111110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_LC_11_16_7  (
            .in0(N__17811),
            .in1(N__16224),
            .in2(N__15472),
            .in3(N__17563),
            .lcout(\this_vga_signals.g1_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_11_17_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_11_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_11_17_2  (
            .in0(N__15469),
            .in1(N__15451),
            .in2(_gnd_net_),
            .in3(N__27822),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_11_17_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_11_17_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_11_17_4  (
            .in0(N__15436),
            .in1(N__15421),
            .in2(_gnd_net_),
            .in3(N__27821),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_11_17_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_11_17_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_wclke_3_LC_11_17_5  (
            .in0(N__25723),
            .in1(N__24576),
            .in2(N__23350),
            .in3(N__20800),
            .lcout(\this_sprites_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6 .LUT_INIT=16'b0101011101010011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6  (
            .in0(N__16869),
            .in1(N__16803),
            .in2(N__16673),
            .in3(N__16739),
            .lcout(\this_vga_ramdac.m6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_18_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_18_0 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_18_0  (
            .in0(N__15379),
            .in1(N__27459),
            .in2(N__15369),
            .in3(N__15861),
            .lcout(\this_vga_ramdac.N_2871_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31995),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.G_384_LC_11_18_1 .C_ON=1'b0;
    defparam \this_ppu.G_384_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.G_384_LC_11_18_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.G_384_LC_11_18_1  (
            .in0(N__15799),
            .in1(N__15816),
            .in2(_gnd_net_),
            .in3(N__15807),
            .lcout(G_384),
            .ltout(G_384_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_18_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_18_2 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_18_2  (
            .in0(N__15339),
            .in1(N__16594),
            .in2(N__15352),
            .in3(N__27461),
            .lcout(\this_vga_ramdac.N_2872_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31995),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_11_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_11_18_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_11_18_5  (
            .in0(N__16031),
            .in1(N__16016),
            .in2(_gnd_net_),
            .in3(N__16000),
            .lcout(\this_vga_signals.line_clk_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_11_18_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_11_18_6 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_11_18_6  (
            .in0(N__16879),
            .in1(N__27460),
            .in2(N__15834),
            .in3(N__15862),
            .lcout(\this_vga_ramdac.N_2873_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31995),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_11_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_11_18_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__15817),
            .in2(_gnd_net_),
            .in3(N__15808),
            .lcout(M_this_vga_signals_pixel_clk_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31995),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIBSKN5_1_LC_11_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIBSKN5_1_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIBSKN5_1_LC_11_19_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIBSKN5_1_LC_11_19_1  (
            .in0(N__15659),
            .in1(N__15513),
            .in2(_gnd_net_),
            .in3(N__21972),
            .lcout(\this_ppu.un1_M_vaddress_q_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_11_20_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_11_20_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_6_0_wclke_3_LC_11_20_5  (
            .in0(N__25716),
            .in1(N__24567),
            .in2(N__23349),
            .in3(N__20808),
            .lcout(\this_sprites_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_0_LC_11_21_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_0_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_0_LC_11_21_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_ppu.M_vaddress_q_0_LC_11_21_2  (
            .in0(N__22008),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15648),
            .lcout(M_this_ppu_vram_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32016),
            .ce(),
            .sr(N__21466));
    defparam \this_ppu.M_vaddress_q_1_LC_11_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_1_LC_11_21_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_1_LC_11_21_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_ppu.M_vaddress_q_1_LC_11_21_4  (
            .in0(N__22009),
            .in1(N__15647),
            .in2(_gnd_net_),
            .in3(N__15505),
            .lcout(M_this_ppu_sprites_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32016),
            .ce(),
            .sr(N__21466));
    defparam \this_ppu.M_vaddress_q_2_LC_11_23_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_2_LC_11_23_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_2_LC_11_23_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_vaddress_q_2_LC_11_23_3  (
            .in0(N__15655),
            .in1(N__15512),
            .in2(N__20352),
            .in3(N__22023),
            .lcout(M_this_ppu_sprites_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32032),
            .ce(),
            .sr(N__21492));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGE761_6_LC_12_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGE761_6_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGE761_6_LC_12_11_1 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGE761_6_LC_12_11_1  (
            .in0(N__18104),
            .in1(N__19693),
            .in2(_gnd_net_),
            .in3(N__19513),
            .lcout(\this_vga_signals.vaddress_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_2_LC_12_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_2_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_2_LC_12_12_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_2_LC_12_12_0  (
            .in0(N__19520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17343),
            .lcout(\this_vga_signals.vaddress_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_12_4 .LUT_INIT=16'b1011001000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_12_4  (
            .in0(N__16183),
            .in1(N__17235),
            .in2(N__16141),
            .in3(N__17915),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_12_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_12_12_5 .LUT_INIT=16'b0011001110100101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_LC_12_12_5  (
            .in0(N__19707),
            .in1(N__16087),
            .in2(N__16078),
            .in3(N__17461),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_12_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_12_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_12_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNINM635_5_LC_12_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNINM635_5_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNINM635_5_LC_12_13_0 .LUT_INIT=16'b0001011110110010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNINM635_5_LC_12_13_0  (
            .in0(N__19141),
            .in1(N__19752),
            .in2(N__19706),
            .in3(N__16075),
            .lcout(\this_vga_signals.i2_mux ),
            .ltout(\this_vga_signals.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5BS7N_5_LC_12_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5BS7N_5_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5BS7N_5_LC_12_13_1 .LUT_INIT=16'b0000111101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5BS7N_5_LC_12_13_1  (
            .in0(N__19675),
            .in1(N__17836),
            .in2(N__16060),
            .in3(N__17465),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNI5BS7NZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m4_0_LC_12_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m4_0_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m4_0_LC_12_13_2 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m4_0_LC_12_13_2  (
            .in0(N__18972),
            .in1(N__19525),
            .in2(_gnd_net_),
            .in3(N__18330),
            .lcout(\this_vga_signals.if_i2_mux ),
            .ltout(\this_vga_signals.if_i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_12_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_12_13_3 .LUT_INIT=16'b0000100111111001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_17_LC_12_13_3  (
            .in0(N__17092),
            .in1(N__19680),
            .in2(N__16057),
            .in3(N__17350),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_7_LC_12_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_7_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_7_LC_12_13_4 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_7_LC_12_13_4  (
            .in0(N__19138),
            .in1(N__17650),
            .in2(_gnd_net_),
            .in3(N__18328),
            .lcout(\this_vga_signals.g1_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_12_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_12_13_5 .LUT_INIT=16'b1011001001010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_LC_12_13_5  (
            .in0(N__16050),
            .in1(N__17234),
            .in2(N__17508),
            .in3(N__17916),
            .lcout(\this_vga_signals.g1_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_12_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_12_13_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_23_LC_12_13_6  (
            .in0(N__19139),
            .in1(N__19671),
            .in2(_gnd_net_),
            .in3(N__19751),
            .lcout(\this_vga_signals.if_N_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_12_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_12_13_7 .LUT_INIT=16'b0001110011011101;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_LC_12_13_7  (
            .in0(N__18329),
            .in1(N__19140),
            .in2(N__19704),
            .in3(N__16246),
            .lcout(\this_vga_signals.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVRE454_5_LC_12_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVRE454_5_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVRE454_5_LC_12_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIVRE454_5_LC_12_14_0  (
            .in0(N__16240),
            .in1(N__16234),
            .in2(N__16228),
            .in3(N__16971),
            .lcout(\this_vga_signals.i14_mux_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x0_LC_12_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x0_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x0_LC_12_14_1 .LUT_INIT=16'b0110011000110110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x0_LC_12_14_1  (
            .in0(N__16311),
            .in1(N__19000),
            .in2(N__18389),
            .in3(N__19523),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_axb1_0_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_ns_LC_12_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_ns_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_ns_LC_12_14_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_ns_LC_12_14_2  (
            .in0(N__17658),
            .in1(_gnd_net_),
            .in2(N__16210),
            .in3(N__16204),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_0 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axb1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_6_LC_12_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_6_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_6_LC_12_14_3 .LUT_INIT=16'b0111111111110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_6_LC_12_14_3  (
            .in0(N__17804),
            .in1(N__16252),
            .in2(N__16207),
            .in3(N__17518),
            .lcout(\this_vga_signals.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_14_4 .LUT_INIT=16'b0110000011111001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_14_4  (
            .in0(N__19521),
            .in1(N__18964),
            .in2(N__16282),
            .in3(N__17589),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_4_LC_12_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_4_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_4_LC_12_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_4_LC_12_14_5  (
            .in0(N__18965),
            .in1(N__19522),
            .in2(_gnd_net_),
            .in3(N__17657),
            .lcout(\this_vga_signals.g0_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x1_LC_12_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x1_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x1_LC_12_14_6 .LUT_INIT=16'b1111000001001011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_0_x1_LC_12_14_6  (
            .in0(N__19524),
            .in1(N__18356),
            .in2(N__19014),
            .in3(N__16312),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_0_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_12_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_12_14_7 .LUT_INIT=16'b1111100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_LC_12_14_7  (
            .in0(N__16384),
            .in1(N__16375),
            .in2(N__19005),
            .in3(N__18421),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHM0ARA_5_LC_12_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHM0ARA_5_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHM0ARA_5_LC_12_15_0 .LUT_INIT=16'b0110100111000011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHM0ARA_5_LC_12_15_0  (
            .in0(N__16366),
            .in1(N__16360),
            .in2(N__17689),
            .in3(N__16354),
            .lcout(\this_vga_signals.i13_mux_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI3HO5K_LC_12_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI3HO5K_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI3HO5K_LC_12_15_1 .LUT_INIT=16'b0011011100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNI3HO5K_LC_12_15_1  (
            .in0(N__17647),
            .in1(N__16348),
            .in2(N__19527),
            .in3(N__18355),
            .lcout(),
            .ltout(\this_vga_signals.g1_N_4L5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5E1_LC_12_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5E1_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5E1_LC_12_15_2 .LUT_INIT=16'b1100100100110110;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5E1_LC_12_15_2  (
            .in0(N__19356),
            .in1(N__16327),
            .in2(N__16318),
            .in3(N__17649),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_4_rep2_esr_RNIREU5EZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIAO8TO2_2_LC_12_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIAO8TO2_2_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIAO8TO2_2_LC_12_15_3 .LUT_INIT=16'b0010101101001101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIAO8TO2_2_LC_12_15_3  (
            .in0(N__17805),
            .in1(N__19010),
            .in2(N__16315),
            .in3(N__18230),
            .lcout(\this_vga_signals.m21_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_520_LC_12_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_520_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_520_LC_12_15_4 .LUT_INIT=16'b1001110010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_520_LC_12_15_4  (
            .in0(N__16308),
            .in1(N__17646),
            .in2(N__19526),
            .in3(N__18327),
            .lcout(if_generate_plus_mult1_un68_sum_axb1_520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_12_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_12_15_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_1_LC_12_15_5  (
            .in0(N__17648),
            .in1(_gnd_net_),
            .in2(N__19253),
            .in3(N__19009),
            .lcout(\this_vga_signals.g0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_15_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_15_6  (
            .in0(N__18354),
            .in1(N__16281),
            .in2(_gnd_net_),
            .in3(N__16261),
            .lcout(\this_vga_signals.mult1_un61_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_12_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_12_15_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_LC_12_15_7  (
            .in0(N__19221),
            .in1(N__19008),
            .in2(N__16255),
            .in3(N__18264),
            .lcout(\this_vga_signals.g0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_LC_12_16_0 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.line_clk.M_last_q_LC_12_16_0 .LUT_INIT=16'b1011000011010000;
    LogicCell40 \this_ppu.line_clk.M_last_q_LC_12_16_0  (
            .in0(N__17403),
            .in1(N__16467),
            .in2(N__16402),
            .in3(N__16560),
            .lcout(\this_ppu.line_clk.M_last_qZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31973),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_12_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_12_16_1 .LUT_INIT=16'b0101011010101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_LC_12_16_1  (
            .in0(N__16972),
            .in1(N__16957),
            .in2(N__16939),
            .in3(N__17595),
            .lcout(\this_vga_signals.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKBOI74_4_LC_12_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKBOI74_4_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKBOI74_4_LC_12_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIKBOI74_4_LC_12_16_5  (
            .in0(N__16924),
            .in1(N__18268),
            .in2(N__19258),
            .in3(N__16918),
            .lcout(\this_vga_signals.m21_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_17_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_17_4 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_17_4  (
            .in0(N__16912),
            .in1(N__16900),
            .in2(N__23203),
            .in3(N__19312),
            .lcout(M_this_ppu_vram_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_5_LC_12_18_0 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_5_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_5_LC_12_18_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIMRAD5_5_LC_12_18_0  (
            .in0(N__20099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20028),
            .lcout(\this_ppu.M_last_q_RNIMRAD5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_18_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_18_1 .LUT_INIT=16'b0010110100010111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_18_1  (
            .in0(N__16644),
            .in1(N__16743),
            .in2(N__16804),
            .in3(N__16855),
            .lcout(\this_vga_ramdac.m16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_12_18_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_12_18_2 .LUT_INIT=16'b0001001101011101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_12_18_2  (
            .in0(N__16854),
            .in1(N__16791),
            .in2(N__16752),
            .in3(N__16645),
            .lcout(\this_vga_ramdac.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUNVB4_7_LC_12_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUNVB4_7_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUNVB4_7_LC_12_18_4 .LUT_INIT=16'b1101101100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIUNVB4_7_LC_12_18_4  (
            .in0(N__16586),
            .in1(N__17404),
            .in2(N__16503),
            .in3(N__16395),
            .lcout(M_this_vga_signals_line_clk_0),
            .ltout(M_this_vga_signals_line_clk_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_LC_12_18_5 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_LC_12_18_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIMRAD5_LC_12_18_5  (
            .in0(N__18750),
            .in1(N__20608),
            .in2(N__17086),
            .in3(N__20098),
            .lcout(\this_ppu.M_state_d_0_sqmuxa ),
            .ltout(\this_ppu.M_state_d_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_1_LC_12_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_1_LC_12_18_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_1_LC_12_18_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_ppu.M_count_q_1_LC_12_18_6  (
            .in0(N__18457),
            .in1(N__20184),
            .in2(N__17083),
            .in3(N__27482),
            .lcout(\this_ppu.M_count_qZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31988),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_0_LC_12_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_0_LC_12_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_0_LC_12_18_7 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \this_ppu.M_state_q_0_LC_12_18_7  (
            .in0(N__27481),
            .in1(N__20100),
            .in2(_gnd_net_),
            .in3(N__21994),
            .lcout(\this_ppu.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31988),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_12_19_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_12_19_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_12_19_1  (
            .in0(N__17080),
            .in1(N__17065),
            .in2(_gnd_net_),
            .in3(N__27820),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_4_LC_12_19_3 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_4_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_4_LC_12_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIMRAD5_4_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__20107),
            .in2(_gnd_net_),
            .in3(N__20023),
            .lcout(\this_ppu.M_last_q_RNIMRAD5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_0_c_RNO_LC_12_19_5 .C_ON=1'b0;
    defparam \this_ppu.un1_M_count_q_1_cry_0_0_c_RNO_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_0_c_RNO_LC_12_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_0_c_RNO_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__20106),
            .in2(_gnd_net_),
            .in3(N__20022),
            .lcout(\this_ppu.un1_M_count_q_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_12_20_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_12_20_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_12_20_4  (
            .in0(N__17053),
            .in1(N__17041),
            .in2(_gnd_net_),
            .in3(N__27800),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIQKTIG_LC_12_21_5 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIQKTIG_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIQKTIG_LC_12_21_5 .LUT_INIT=16'b1111111110001010;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIQKTIG_LC_12_21_5  (
            .in0(N__22001),
            .in1(N__21641),
            .in2(N__17028),
            .in3(N__27480),
            .lcout(\this_ppu.M_last_q_RNIQKTIG ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_13_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_13_12_0 .LUT_INIT=16'b1010000001011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_LC_13_12_0  (
            .in0(N__19217),
            .in1(_gnd_net_),
            .in2(N__19714),
            .in3(N__18103),
            .lcout(),
            .ltout(\this_vga_signals.g1_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_13_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_13_12_1 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_LC_13_12_1  (
            .in0(N__17509),
            .in1(N__17386),
            .in2(N__17482),
            .in3(N__17236),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_12_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__18527),
            .in2(_gnd_net_),
            .in3(N__18579),
            .lcout(\this_vga_signals.M_vcounter_d7lt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_LC_13_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_LC_13_13_0 .LUT_INIT=16'b0101010111000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_LC_13_13_0  (
            .in0(N__17479),
            .in1(N__17473),
            .in2(N__19705),
            .in3(N__17466),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIJPU72_2_LC_13_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIJPU72_2_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIJPU72_2_LC_13_13_1 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIJPU72_2_LC_13_13_1  (
            .in0(N__17801),
            .in1(N__17440),
            .in2(N__19006),
            .in3(N__19517),
            .lcout(\this_vga_signals.M_vcounter_d7lt9_1 ),
            .ltout(\this_vga_signals.M_vcounter_d7lt9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIAEPU2_6_LC_13_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIAEPU2_6_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIAEPU2_6_LC_13_13_2 .LUT_INIT=16'b0000000011110101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIAEPU2_6_LC_13_13_2  (
            .in0(N__19676),
            .in1(_gnd_net_),
            .in2(N__17407),
            .in3(N__18102),
            .lcout(\this_vga_signals.un4_lvisibility_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_1_LC_13_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_1_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_1_LC_13_13_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_1_LC_13_13_4  (
            .in0(N__19518),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17338),
            .lcout(\this_vga_signals.vaddress_1_5 ),
            .ltout(\this_vga_signals.vaddress_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_13_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_13_13_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_18_LC_13_13_5  (
            .in0(N__17382),
            .in1(N__17365),
            .in2(N__17353),
            .in3(N__17233),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_0_LC_13_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_0_LC_13_13_6 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_0_LC_13_13_6  (
            .in0(N__19519),
            .in1(N__18101),
            .in2(_gnd_net_),
            .in3(N__17339),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_13_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_13_13_7 .LUT_INIT=16'b1011001000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_4_LC_13_13_7  (
            .in0(N__17242),
            .in1(N__17232),
            .in2(N__17095),
            .in3(N__17929),
            .lcout(\this_vga_signals.g1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNITP439_0_2_LC_13_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNITP439_0_2_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNITP439_0_2_LC_13_14_0 .LUT_INIT=16'b1001101001100101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNITP439_0_2_LC_13_14_0  (
            .in0(N__18371),
            .in1(N__18978),
            .in2(N__19249),
            .in3(N__17803),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_RNITP439_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIFPMH71_2_LC_13_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIFPMH71_2_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIFPMH71_2_LC_13_14_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIFPMH71_2_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__18834),
            .in2(N__17692),
            .in3(N__17551),
            .lcout(\this_vga_signals.m16_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_13_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_13_14_3 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_13_14_3  (
            .in0(N__17674),
            .in1(N__18368),
            .in2(N__19247),
            .in3(N__17599),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_13_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_13_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__18976),
            .in2(N__17566),
            .in3(N__18262),
            .lcout(\this_vga_signals.g0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNITP439_2_LC_13_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNITP439_2_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNITP439_2_LC_13_14_5 .LUT_INIT=16'b1100011000111001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNITP439_2_LC_13_14_5  (
            .in0(N__18977),
            .in1(N__17802),
            .in2(N__19248),
            .in3(N__18369),
            .lcout(\this_vga_signals.M_vcounter_q_RNITP439Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_14_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_14_6  (
            .in0(N__18370),
            .in1(N__18263),
            .in2(N__18842),
            .in3(N__18217),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_13_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_13_14_7 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_0_LC_13_14_7  (
            .in0(N__17545),
            .in1(N__17536),
            .in2(N__17530),
            .in3(N__18218),
            .lcout(\this_vga_signals.g0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_13_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_13_15_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_13_15_0  (
            .in0(N__18835),
            .in1(N__18265),
            .in2(_gnd_net_),
            .in3(N__18219),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_1_LC_13_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_1_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_1_LC_13_15_1 .LUT_INIT=16'b0011100110011100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_1_LC_13_15_1  (
            .in0(N__19012),
            .in1(N__19216),
            .in2(N__17512),
            .in3(N__17806),
            .lcout(\this_vga_signals.mult1_un82_sum_c3_0_N_4L5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_3_LC_13_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_3_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_3_LC_13_15_3 .LUT_INIT=16'b1001110010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_3_LC_13_15_3  (
            .in0(N__18439),
            .in1(N__18427),
            .in2(N__19254),
            .in3(N__18393),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_13_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_13_15_4 .LUT_INIT=16'b1010110111011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_21_LC_13_15_4  (
            .in0(N__18420),
            .in1(N__19011),
            .in2(N__18409),
            .in3(N__18221),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_LC_13_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_LC_13_15_5 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_LC_13_15_5  (
            .in0(N__18406),
            .in1(N__17807),
            .in2(N__18400),
            .in3(N__18169),
            .lcout(\this_vga_signals.N_5_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_15_6  (
            .in0(N__18392),
            .in1(N__18266),
            .in2(N__18843),
            .in3(N__18220),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_15_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(N__18805),
            .in2(N__18178),
            .in3(N__18175),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_LC_13_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_LC_13_16_0 .LUT_INIT=16'b1010101011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_LC_13_16_0  (
            .in0(N__18163),
            .in1(N__18145),
            .in2(N__18130),
            .in3(N__17944),
            .lcout(\this_vga_signals.g1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI1RPOO2_1_LC_13_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI1RPOO2_1_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI1RPOO2_1_LC_13_16_1 .LUT_INIT=16'b0001010000101000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI1RPOO2_1_LC_13_16_1  (
            .in0(N__17824),
            .in1(N__17817),
            .in2(N__18548),
            .in3(N__17722),
            .lcout(),
            .ltout(\this_vga_signals.N_25_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5P1Q0M_4_LC_13_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5P1Q0M_4_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5P1Q0M_4_LC_13_16_2 .LUT_INIT=16'b1010100101011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5P1Q0M_4_LC_13_16_2  (
            .in0(N__17713),
            .in1(N__17707),
            .in2(N__17695),
            .in3(N__18625),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGBAMTL1_9_LC_13_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGBAMTL1_9_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGBAMTL1_9_LC_13_16_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIGBAMTL1_9_LC_13_16_3  (
            .in0(N__21000),
            .in1(N__18619),
            .in2(N__18610),
            .in3(N__18481),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_LC_13_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_LC_13_16_5 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_N_4L5_LC_13_16_5  (
            .in0(N__18586),
            .in1(N__18844),
            .in2(N__18549),
            .in3(N__18556),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_N_4L5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_13_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_13_16_6 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_m2_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(N__18544),
            .in2(N__18490),
            .in3(N__18487),
            .lcout(\this_vga_signals.mult1_un82_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_2_LC_13_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_2_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_2_LC_13_17_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_count_q_2_LC_13_17_4  (
            .in0(N__27450),
            .in1(N__21990),
            .in2(N__20188),
            .in3(N__18448),
            .lcout(\this_ppu.M_count_qZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31974),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_13_17_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_13_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18475),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31974),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_0_c_LC_13_18_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_0_c_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_0_c_LC_13_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_0_c_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__18463),
            .in2(N__19812),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\this_ppu.un1_M_count_q_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_1_LC_13_18_1 .C_ON=1'b1;
    defparam \this_ppu.M_count_q_RNO_0_1_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_1_LC_13_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_count_q_RNO_0_1_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__18721),
            .in2(N__19851),
            .in3(N__18451),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_0 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_2_LC_13_18_2 .C_ON=1'b1;
    defparam \this_ppu.M_count_q_RNO_0_2_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_2_LC_13_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_count_q_RNO_0_2_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__18637),
            .in2(N__19834),
            .in3(N__18442),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_3_LC_13_18_3 .C_ON=1'b1;
    defparam \this_ppu.M_count_q_RNO_0_3_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_3_LC_13_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_count_q_RNO_0_3_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__20272),
            .in2(N__20259),
            .in3(N__18670),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_2 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_4_LC_13_18_4 .C_ON=1'b1;
    defparam \this_ppu.M_count_q_RNO_0_4_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_4_LC_13_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_count_q_RNO_0_4_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__18667),
            .in2(N__20242),
            .in3(N__18661),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_3 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_5_LC_13_18_5 .C_ON=1'b1;
    defparam \this_ppu.M_count_q_RNO_0_5_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_5_LC_13_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_count_q_RNO_0_5_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__18643),
            .in2(N__20122),
            .in3(N__18658),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_4 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_6_LC_13_18_6 .C_ON=1'b1;
    defparam \this_ppu.M_count_q_RNO_0_6_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_6_LC_13_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_count_q_RNO_0_6_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__18655),
            .in2(N__20227),
            .in3(N__18649),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_5 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_7_LC_13_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_7_LC_13_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_7_LC_13_18_7 .LUT_INIT=16'b0101000101010100;
    LogicCell40 \this_ppu.M_count_q_7_LC_13_18_7  (
            .in0(N__20159),
            .in1(N__19990),
            .in2(N__22011),
            .in3(N__18646),
            .lcout(\this_ppu.M_count_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31981),
            .ce(),
            .sr(N__32392));
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_1_LC_13_19_0 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_1_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_1_LC_13_19_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIMRAD5_1_LC_13_19_0  (
            .in0(N__20025),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20094),
            .lcout(\this_ppu.M_last_q_RNIMRAD5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_0_LC_13_19_1 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_0_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_0_LC_13_19_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIMRAD5_0_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__20092),
            .in2(_gnd_net_),
            .in3(N__20024),
            .lcout(\this_ppu.M_last_q_RNIMRAD5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_4_LC_13_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_4_LC_13_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_4_LC_13_19_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_count_q_4_LC_13_19_2  (
            .in0(N__27452),
            .in1(N__21988),
            .in2(N__20177),
            .in3(N__18631),
            .lcout(\this_ppu.M_count_qZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31989),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_0_LC_13_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNO_0_0_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_0_LC_13_19_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_count_q_RNO_0_0_LC_13_19_3  (
            .in0(N__19813),
            .in1(N__20093),
            .in2(_gnd_net_),
            .in3(N__20026),
            .lcout(),
            .ltout(\this_ppu.un1_M_count_q_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_0_LC_13_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_0_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_0_LC_13_19_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_ppu.M_count_q_0_LC_13_19_4  (
            .in0(N__27451),
            .in1(N__20160),
            .in2(N__18760),
            .in3(N__21989),
            .lcout(\this_ppu.M_count_qZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31989),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_6_LC_13_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_6_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_6_LC_13_19_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_count_q_6_LC_13_19_5  (
            .in0(N__21987),
            .in1(N__27453),
            .in2(N__20175),
            .in3(N__18757),
            .lcout(\this_ppu.M_count_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31989),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIMMU35_LC_13_19_6 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIMMU35_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIMMU35_LC_13_19_6 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIMMU35_LC_13_19_6  (
            .in0(N__18751),
            .in1(N__20601),
            .in2(_gnd_net_),
            .in3(N__18730),
            .lcout(\this_ppu.N_82_i ),
            .ltout(\this_ppu.N_82_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_3_LC_13_19_7 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_3_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_3_LC_13_19_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIMRAD5_3_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18724),
            .in3(N__20091),
            .lcout(\this_ppu.M_last_q_RNIMRAD5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_3_LC_13_22_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_3_LC_13_22_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_3_LC_13_22_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_vaddress_q_3_LC_13_22_7  (
            .in0(N__20357),
            .in1(N__20482),
            .in2(_gnd_net_),
            .in3(N__20304),
            .lcout(M_this_ppu_map_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32008),
            .ce(),
            .sr(N__21467));
    defparam \this_ppu.M_vaddress_q_4_LC_13_23_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_4_LC_13_23_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_4_LC_13_23_4 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_ppu.M_vaddress_q_4_LC_13_23_4  (
            .in0(N__20525),
            .in1(N__20483),
            .in2(N__20356),
            .in3(N__20305),
            .lcout(M_this_ppu_map_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32017),
            .ce(),
            .sr(N__21493));
    defparam \this_reset_cond.M_stage_q_4_LC_14_12_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_4_LC_14_12_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_4_LC_14_12_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_4_LC_14_12_1  (
            .in0(N__28471),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18715),
            .lcout(\this_reset_cond.M_stage_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31945),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_14_12_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_14_12_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_14_12_3  (
            .in0(N__28470),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20710),
            .lcout(\this_reset_cond.M_stage_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31945),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_14_13_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_14_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_14_13_2  (
            .in0(N__27823),
            .in1(N__18709),
            .in2(_gnd_net_),
            .in3(N__18691),
            .lcout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_14_13_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_14_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_14_13_3  (
            .in0(N__27824),
            .in1(N__19789),
            .in2(_gnd_net_),
            .in3(N__19768),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_14_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_14_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_13_LC_14_14_1  (
            .in0(N__19753),
            .in1(N__19710),
            .in2(_gnd_net_),
            .in3(N__19528),
            .lcout(\this_vga_signals.if_N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_5_LC_14_14_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_5_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_5_LC_14_14_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_5_LC_14_14_2  (
            .in0(N__28481),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19333),
            .lcout(\this_reset_cond.M_stage_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31951),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_14_14_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_14_14_3 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_14_14_3  (
            .in0(N__23185),
            .in1(N__19324),
            .in2(N__29672),
            .in3(N__19318),
            .lcout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_6_LC_14_14_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_6_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_6_LC_14_14_4 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \this_reset_cond.M_stage_q_6_LC_14_14_4  (
            .in0(N__19300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28482),
            .lcout(\this_reset_cond.M_stage_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31951),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_14_14_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_14_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_14_14_6  (
            .in0(N__27825),
            .in1(N__19294),
            .in2(_gnd_net_),
            .in3(N__19279),
            .lcout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_14_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_14_15_1 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_14_15_1  (
            .in0(N__19256),
            .in1(N__19007),
            .in2(_gnd_net_),
            .in3(N__18830),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_14_15_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_14_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_14_15_2  (
            .in0(N__27762),
            .in1(N__18799),
            .in2(_gnd_net_),
            .in3(N__18781),
            .lcout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_14_16_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_14_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_14_16_4  (
            .in0(N__27826),
            .in1(N__19978),
            .in2(_gnd_net_),
            .in3(N__19960),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_14_16_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_14_16_5 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_14_16_5  (
            .in0(N__29645),
            .in1(N__23161),
            .in2(N__19945),
            .in3(N__19942),
            .lcout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_14_17_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_14_17_3 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_14_17_3  (
            .in0(N__23198),
            .in1(N__20668),
            .in2(N__29673),
            .in3(N__19936),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_14_17_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_14_17_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_14_17_4  (
            .in0(N__23192),
            .in1(N__19927),
            .in2(N__19915),
            .in3(N__19861),
            .lcout(M_this_ppu_vram_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_14_17_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_14_17_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_14_17_7  (
            .in0(N__19897),
            .in1(N__19882),
            .in2(_gnd_net_),
            .in3(N__27819),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_1_LC_14_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_14_18_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_state_q_RNO_0_1_LC_14_18_0  (
            .in0(N__20203),
            .in1(N__20209),
            .in2(_gnd_net_),
            .in3(N__20097),
            .lcout(),
            .ltout(\this_ppu.N_91_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_1_LC_14_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_1_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_1_LC_14_18_1 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \this_ppu.M_state_q_1_LC_14_18_1  (
            .in0(N__20613),
            .in1(N__20577),
            .in2(N__19855),
            .in3(N__32436),
            .lcout(\this_ppu.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31975),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNI230G_0_LC_14_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNI230G_0_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNI230G_0_LC_14_18_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_count_q_RNI230G_0_LC_14_18_2  (
            .in0(N__19852),
            .in1(N__19833),
            .in2(N__20260),
            .in3(N__19808),
            .lcout(\this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI05C9_1_LC_14_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI05C9_1_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI05C9_1_LC_14_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.M_state_q_RNI05C9_1_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20576),
            .lcout(\this_ppu.M_state_q_i_1 ),
            .ltout(\this_ppu.M_state_q_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_2_LC_14_18_4 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_2_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIMRAD5_2_LC_14_18_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIMRAD5_2_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20275),
            .in3(N__20027),
            .lcout(\this_ppu.M_last_q_RNIMRAD5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_3_LC_14_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_3_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_3_LC_14_18_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_count_q_3_LC_14_18_6  (
            .in0(N__27496),
            .in1(N__22010),
            .in2(N__20176),
            .in3(N__20266),
            .lcout(\this_ppu.M_count_qZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31975),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIIJ0G_7_LC_14_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIIJ0G_7_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIIJ0G_7_LC_14_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_count_q_RNIIJ0G_7_LC_14_19_0  (
            .in0(N__20238),
            .in1(N__20220),
            .in2(N__20041),
            .in3(N__20118),
            .lcout(\this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4 ),
            .ltout(\this_ppu.M_state_d_0_sqmuxa_1_0_a3_8_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIJVOI1_0_LC_14_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIJVOI1_0_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIJVOI1_0_LC_14_19_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_state_q_RNIJVOI1_0_LC_14_19_1  (
            .in0(N__20202),
            .in1(N__20617),
            .in2(N__20191),
            .in3(N__20095),
            .lcout(\this_ppu.M_state_d_0_sqmuxa_1 ),
            .ltout(\this_ppu.M_state_d_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_5_LC_14_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_5_LC_14_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_5_LC_14_19_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_count_q_5_LC_14_19_2  (
            .in0(N__27495),
            .in1(N__22022),
            .in2(N__20131),
            .in3(N__20128),
            .lcout(\this_ppu.M_count_qZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31982),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_7_LC_14_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_14_19_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_count_q_RNO_0_7_LC_14_19_3  (
            .in0(N__20096),
            .in1(N__20040),
            .in2(_gnd_net_),
            .in3(N__20029),
            .lcout(\this_ppu.un1_M_count_q_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_15_11_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_15_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28467),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31941),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_15_11_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_15_11_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_15_11_1  (
            .in0(N__28468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19984),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31941),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_15_11_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_15_11_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_15_11_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_15_11_5  (
            .in0(N__28469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20716),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31941),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_15_16_3.C_ON=1'b0;
    defparam M_this_state_q_4_LC_15_16_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_15_16_3.LUT_INIT=16'b0000101011001110;
    LogicCell40 M_this_state_q_4_LC_15_16_3 (
            .in0(N__25789),
            .in1(N__27554),
            .in2(N__27002),
            .in3(N__32830),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31956),
            .ce(),
            .sr(N__32390));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_15_17_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_15_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_15_17_2  (
            .in0(N__27818),
            .in1(N__20704),
            .in2(_gnd_net_),
            .in3(N__20686),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_15_17_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_15_17_4 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_15_17_4  (
            .in0(N__20662),
            .in1(N__20653),
            .in2(N__23199),
            .in3(N__20641),
            .lcout(M_this_ppu_vram_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIV8OI_1_LC_15_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIV8OI_1_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIV8OI_1_LC_15_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_state_q_RNIV8OI_1_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__20612),
            .in2(_gnd_net_),
            .in3(N__20578),
            .lcout(M_this_ppu_vram_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_15_19_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_15_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_7_0_wclke_3_LC_15_19_3  (
            .in0(N__25708),
            .in1(N__24561),
            .in2(N__23319),
            .in3(N__20788),
            .lcout(\this_sprites_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_m_2_LC_15_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_2_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_2_LC_15_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_2_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__30306),
            .in2(_gnd_net_),
            .in3(N__30597),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNI25476_4_LC_15_23_0 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI25476_4_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI25476_4_LC_15_23_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNI25476_4_LC_15_23_0  (
            .in0(N__20529),
            .in1(N__20493),
            .in2(N__20364),
            .in3(N__20303),
            .lcout(\this_ppu.un1_M_vaddress_q_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_6_LC_15_24_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_6_LC_15_24_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_6_LC_15_24_7 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_ppu.M_vaddress_q_6_LC_15_24_7  (
            .in0(N__21551),
            .in1(N__21522),
            .in2(_gnd_net_),
            .in3(N__23885),
            .lcout(\this_ppu.M_vaddress_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32009),
            .ce(),
            .sr(N__21503));
    defparam \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(N__23712),
            .in2(_gnd_net_),
            .in3(N__24469),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_16_14_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_16_14_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_16_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20878),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31944),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_en_0_LC_16_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_en_0_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_en_0_LC_16_15_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_en_0_LC_16_15_0  (
            .in0(N__27924),
            .in1(N__27207),
            .in2(_gnd_net_),
            .in3(N__32638),
            .lcout(M_this_sprites_ram_write_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI2S2S_13_LC_16_15_2.C_ON=1'b0;
    defparam M_this_state_q_RNI2S2S_13_LC_16_15_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI2S2S_13_LC_16_15_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_state_q_RNI2S2S_13_LC_16_15_2 (
            .in0(N__27925),
            .in1(N__27208),
            .in2(N__31327),
            .in3(N__28017),
            .lcout(M_this_state_q_RNI2S2SZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_fast_15_LC_16_16_0.C_ON=1'b0;
    defparam M_this_state_q_fast_15_LC_16_16_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_fast_15_LC_16_16_0.LUT_INIT=16'b0010001000100000;
    LogicCell40 M_this_state_q_fast_15_LC_16_16_0 (
            .in0(N__27216),
            .in1(N__27169),
            .in2(N__27096),
            .in3(N__27052),
            .lcout(M_this_state_q_fastZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31949),
            .ce(),
            .sr(N__32388));
    defparam M_this_state_q_14_LC_16_16_1.C_ON=1'b0;
    defparam M_this_state_q_14_LC_16_16_1.SEQ_MODE=4'b1000;
    defparam M_this_state_q_14_LC_16_16_1.LUT_INIT=16'b0000101100001010;
    LogicCell40 M_this_state_q_14_LC_16_16_1 (
            .in0(N__27226),
            .in1(N__28528),
            .in2(N__32851),
            .in3(N__25768),
            .lcout(M_this_state_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31949),
            .ce(),
            .sr(N__32388));
    defparam \this_vga_signals.M_this_state_q_tr43_LC_16_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_tr43_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_tr43_LC_16_16_2 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_vga_signals.M_this_state_q_tr43_LC_16_16_2  (
            .in0(N__27215),
            .in1(N__27168),
            .in2(N__27097),
            .in3(N__27051),
            .lcout(\this_vga_signals.M_this_state_q_ns_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_16_16_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_16_16_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_wclke_3_LC_16_16_4  (
            .in0(N__25725),
            .in1(N__24562),
            .in2(N__23339),
            .in3(N__20769),
            .lcout(\this_sprites_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_16_16_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_16_16_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_wclke_3_LC_16_16_5  (
            .in0(N__20770),
            .in1(N__23323),
            .in2(N__24575),
            .in3(N__25726),
            .lcout(\this_sprites_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_16_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_16_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_16_6  (
            .in0(N__25727),
            .in1(N__24566),
            .in2(N__23340),
            .in3(N__20771),
            .lcout(\this_sprites_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_0_LC_16_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_0_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_0_LC_16_17_0 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_0_LC_16_17_0  (
            .in0(N__22653),
            .in1(N__33818),
            .in2(N__33340),
            .in3(N__21104),
            .lcout(M_this_sprites_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_LC_16_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_LC_16_17_1 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_1_LC_16_17_1  (
            .in0(N__21105),
            .in1(N__33982),
            .in2(N__33642),
            .in3(N__22654),
            .lcout(M_this_sprites_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_16_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_16_17_2 .LUT_INIT=16'b0000000101010101;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_16_17_2  (
            .in0(N__27945),
            .in1(N__25392),
            .in2(N__27227),
            .in3(N__32786),
            .lcout(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ),
            .ltout(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_2_LC_16_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_2_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_2_LC_16_17_3 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_2_LC_16_17_3  (
            .in0(N__33512),
            .in1(N__34212),
            .in2(N__21205),
            .in3(N__22655),
            .lcout(M_this_sprites_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_16_18_4.C_ON=1'b0;
    defparam M_this_state_q_5_LC_16_18_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_16_18_4.LUT_INIT=16'b1011001110100000;
    LogicCell40 M_this_state_q_5_LC_16_18_4 (
            .in0(N__24594),
            .in1(N__32785),
            .in2(N__24042),
            .in3(N__30598),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31961),
            .ce(),
            .sr(N__32389));
    defparam M_this_state_q_12_LC_16_18_7.C_ON=1'b0;
    defparam M_this_state_q_12_LC_16_18_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_12_LC_16_18_7.LUT_INIT=16'b0101010100010000;
    LogicCell40 M_this_state_q_12_LC_16_18_7 (
            .in0(N__32784),
            .in1(N__28524),
            .in2(N__23995),
            .in3(N__27994),
            .lcout(M_this_state_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31961),
            .ce(),
            .sr(N__32389));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_3_LC_16_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_3_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_3_LC_16_19_3 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_3_LC_16_19_3  (
            .in0(N__34347),
            .in1(N__22662),
            .in2(N__33427),
            .in3(N__21109),
            .lcout(M_this_sprites_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNICRTO5_9_LC_16_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICRTO5_9_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICRTO5_9_LC_16_19_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNICRTO5_9_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(N__20991),
            .in2(_gnd_net_),
            .in3(N__20920),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_5_LC_16_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_5_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_5_LC_16_20_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_0_5_LC_16_20_7  (
            .in0(N__27003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26856),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_0_LC_16_22_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_0_LC_16_22_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_0_LC_16_22_2 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \this_ppu.M_haddress_q_0_LC_16_22_2  (
            .in0(N__22252),
            .in1(N__22219),
            .in2(_gnd_net_),
            .in3(N__22027),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31987),
            .ce(),
            .sr(N__25036));
    defparam \this_ppu.M_haddress_q_1_LC_16_22_7 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_1_LC_16_22_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_1_LC_16_22_7 .LUT_INIT=16'b0011110001111000;
    LogicCell40 \this_ppu.M_haddress_q_1_LC_16_22_7  (
            .in0(N__22026),
            .in1(N__22251),
            .in2(N__22066),
            .in3(N__22220),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31987),
            .ce(),
            .sr(N__25036));
    defparam \this_ppu.M_vaddress_q_5_LC_16_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_5_LC_16_23_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_5_LC_16_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_vaddress_q_5_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(N__21521),
            .in2(_gnd_net_),
            .in3(N__21547),
            .lcout(M_this_ppu_map_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31993),
            .ce(),
            .sr(N__21505));
    defparam \this_ppu.M_vaddress_q_7_LC_16_24_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_7_LC_16_24_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_7_LC_16_24_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_ppu.M_vaddress_q_7_LC_16_24_2  (
            .in0(N__21445),
            .in1(N__23886),
            .in2(N__21555),
            .in3(N__21523),
            .lcout(\this_ppu.M_vaddress_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32001),
            .ce(),
            .sr(N__21504));
    defparam \this_ppu.M_vaddress_q_RNI1DAA_7_LC_16_25_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI1DAA_7_LC_16_25_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI1DAA_7_LC_16_25_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_vaddress_q_RNI1DAA_7_LC_16_25_6  (
            .in0(_gnd_net_),
            .in1(N__21444),
            .in2(_gnd_net_),
            .in3(N__23881),
            .lcout(M_this_ppu_map_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_17_13_7.C_ON=1'b0;
    defparam M_this_state_q_2_LC_17_13_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_17_13_7.LUT_INIT=16'b1010000011101100;
    LogicCell40 M_this_state_q_2_LC_17_13_7 (
            .in0(N__24016),
            .in1(N__28198),
            .in2(N__26877),
            .in3(N__32790),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31946),
            .ce(),
            .sr(N__32391));
    defparam \this_vga_signals.M_this_sprites_address_q_m_1_LC_17_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_1_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_1_LC_17_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_1_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__25501),
            .in2(_gnd_net_),
            .in3(N__24474),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_14_1.C_ON=1'b0;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_14_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32431),
            .lcout(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_17_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_17_14_2 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_17_14_2  (
            .in0(N__22855),
            .in1(N__24473),
            .in2(N__34213),
            .in3(N__32777),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_8_LC_17_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_8_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_8_LC_17_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_8_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(N__23002),
            .in2(_gnd_net_),
            .in3(N__28161),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_8_LC_17_15_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_8_LC_17_15_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_8_LC_17_15_4.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_8_LC_17_15_4 (
            .in0(N__21673),
            .in1(N__24151),
            .in2(N__21664),
            .in3(N__22978),
            .lcout(M_this_sprites_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31952),
            .ce(),
            .sr(N__27289));
    defparam \this_vga_signals.un23_i_a2_x1_0_LC_17_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un23_i_a2_x1_0_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un23_i_a2_x1_0_LC_17_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.un23_i_a2_x1_0_LC_17_16_0  (
            .in0(N__31202),
            .in1(N__29616),
            .in2(N__31323),
            .in3(N__25382),
            .lcout(),
            .ltout(\this_vga_signals.un23_i_a2_x1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un23_i_a2_ns_0_LC_17_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un23_i_a2_ns_0_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un23_i_a2_ns_0_LC_17_16_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vga_signals.un23_i_a2_ns_0_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21655),
            .in3(N__21685),
            .lcout(dma_axb0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dma_ac0_5_LC_17_16_3.C_ON=1'b0;
    defparam dma_ac0_5_LC_17_16_3.SEQ_MODE=4'b0000;
    defparam dma_ac0_5_LC_17_16_3.LUT_INIT=16'b0001001100110011;
    LogicCell40 dma_ac0_5_LC_17_16_3 (
            .in0(N__31252),
            .in1(N__21592),
            .in2(N__25447),
            .in3(N__21607),
            .lcout(dma_ac0Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un23_i_a2_4_2_LC_17_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un23_i_a2_4_2_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un23_i_a2_4_2_LC_17_16_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.un23_i_a2_4_2_LC_17_16_4  (
            .in0(N__29617),
            .in1(N__30784),
            .in2(N__27607),
            .in3(N__30609),
            .lcout(this_vga_signals_un23_i_a2_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un23_i_a2_1_3_LC_17_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un23_i_a2_1_3_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un23_i_a2_1_3_LC_17_16_5 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \this_vga_signals.un23_i_a2_1_3_LC_17_16_5  (
            .in0(N__25383),
            .in1(_gnd_net_),
            .in2(N__28040),
            .in3(N__32924),
            .lcout(this_vga_signals_un23_i_a2_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un23_i_a2_3_2_LC_17_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un23_i_a2_3_2_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un23_i_a2_3_2_LC_17_16_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.un23_i_a2_3_2_LC_17_16_6  (
            .in0(N__31316),
            .in1(N__27206),
            .in2(N__27946),
            .in3(N__28027),
            .lcout(),
            .ltout(this_vga_signals_un23_i_a2_3_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dma_c3_LC_17_16_7.C_ON=1'b0;
    defparam dma_c3_LC_17_16_7.SEQ_MODE=4'b0000;
    defparam dma_c3_LC_17_16_7.LUT_INIT=16'b1010000010000000;
    LogicCell40 dma_c3_LC_17_16_7 (
            .in0(N__21601),
            .in1(N__24061),
            .in2(N__21595),
            .in3(N__21585),
            .lcout(dma_c3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNITS9I4_7_LC_17_17_0.C_ON=1'b0;
    defparam M_this_state_q_RNITS9I4_7_LC_17_17_0.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNITS9I4_7_LC_17_17_0.LUT_INIT=16'b0101011101110111;
    LogicCell40 M_this_state_q_RNITS9I4_7_LC_17_17_0 (
            .in0(N__21679),
            .in1(N__21586),
            .in2(N__24076),
            .in3(N__25445),
            .lcout(),
            .ltout(M_this_state_q_RNITS9I4Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIV6UJ7_8_LC_17_17_1.C_ON=1'b0;
    defparam M_this_state_q_RNIV6UJ7_8_LC_17_17_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIV6UJ7_8_LC_17_17_1.LUT_INIT=16'b0000101011001110;
    LogicCell40 M_this_state_q_RNIV6UJ7_8_LC_17_17_1 (
            .in0(N__21910),
            .in1(N__25446),
            .in2(N__21901),
            .in3(N__22393),
            .lcout(dma_ac0_5_i),
            .ltout(dma_ac0_5_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIV6UJ7_0_8_LC_17_17_2.C_ON=1'b0;
    defparam M_this_state_q_RNIV6UJ7_0_8_LC_17_17_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIV6UJ7_0_8_LC_17_17_2.LUT_INIT=16'b0000111100001111;
    LogicCell40 M_this_state_q_RNIV6UJ7_0_8_LC_17_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21874),
            .in3(_gnd_net_),
            .lcout(dma_ac0_5_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_3_LC_17_17_5.C_ON=1'b0;
    defparam M_this_state_q_3_LC_17_17_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_17_17_5.LUT_INIT=16'b1010000011101100;
    LogicCell40 M_this_state_q_3_LC_17_17_5 (
            .in0(N__24052),
            .in1(N__26399),
            .in2(N__22387),
            .in3(N__32788),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31964),
            .ce(),
            .sr(N__32382));
    defparam \this_vga_signals.un23_i_a2_4_0_LC_17_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un23_i_a2_4_0_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un23_i_a2_4_0_LC_17_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.un23_i_a2_4_0_LC_17_17_6  (
            .in0(N__24403),
            .in1(N__30578),
            .in2(N__26425),
            .in3(N__25461),
            .lcout(\this_vga_signals.un23_i_a2_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_17_17_7.C_ON=1'b0;
    defparam M_this_state_q_1_LC_17_17_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_17_17_7.LUT_INIT=16'b0010001011110010;
    LogicCell40 M_this_state_q_1_LC_17_17_7 (
            .in0(N__24012),
            .in1(N__26873),
            .in2(N__24467),
            .in3(N__32787),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31964),
            .ce(),
            .sr(N__32382));
    defparam M_this_state_q_RNI6Q0S_7_LC_17_18_1.C_ON=1'b0;
    defparam M_this_state_q_RNI6Q0S_7_LC_17_18_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI6Q0S_7_LC_17_18_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_state_q_RNI6Q0S_7_LC_17_18_1 (
            .in0(N__29620),
            .in1(N__27621),
            .in2(N__30648),
            .in3(N__30847),
            .lcout(M_this_state_q_RNI6Q0SZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_17_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_17_18_2 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_17_18_2  (
            .in0(N__32774),
            .in1(N__23009),
            .in2(N__33981),
            .in3(N__24431),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_17_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_17_18_3 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_17_18_3  (
            .in0(N__22715),
            .in1(N__34333),
            .in2(N__24466),
            .in3(N__32776),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_17_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_17_18_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_17_18_4  (
            .in0(N__32775),
            .in1(N__23271),
            .in2(N__33538),
            .in3(N__24435),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_3_LC_17_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_3_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_3_LC_17_18_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_0_3_LC_17_18_7  (
            .in0(N__27004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26863),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_13_LC_17_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_13_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_13_LC_17_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_13_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__23272),
            .in2(_gnd_net_),
            .in3(N__28211),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_10_LC_17_19_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_10_LC_17_19_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_10_LC_17_19_7.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_10_LC_17_19_7 (
            .in0(N__22378),
            .in1(N__24175),
            .in2(N__22408),
            .in3(N__22681),
            .lcout(M_this_sprites_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31976),
            .ce(),
            .sr(N__27284));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_17_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_17_20_2 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_17_20_2  (
            .in0(N__25663),
            .in1(N__24455),
            .in2(N__33641),
            .in3(N__32826),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_4_LC_17_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_4_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_4_LC_17_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_4_LC_17_20_7  (
            .in0(N__24454),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26165),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNI21NK5_LC_17_24_1 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNI21NK5_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNI21NK5_LC_17_24_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNI21NK5_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(N__27494),
            .in2(_gnd_net_),
            .in3(N__22024),
            .lcout(\this_ppu.M_last_q_RNI21NK5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIEKA06_1_LC_17_24_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIEKA06_1_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIEKA06_1_LC_17_24_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \this_ppu.M_haddress_q_RNIEKA06_1_LC_17_24_3  (
            .in0(N__22262),
            .in1(N__22224),
            .in2(N__22076),
            .in3(N__22025),
            .lcout(\this_ppu.un1_M_haddress_q_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_2_LC_17_25_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_2_LC_17_25_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_2_LC_17_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_haddress_q_2_LC_17_25_0  (
            .in0(_gnd_net_),
            .in1(N__23428),
            .in2(_gnd_net_),
            .in3(N__23976),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32018),
            .ce(),
            .sr(N__25030));
    defparam \this_vga_signals.M_this_sprites_address_q_m_9_LC_18_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_9_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_9_LC_18_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_9_LC_18_12_0  (
            .in0(N__22859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28160),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_3_LC_18_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_3_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_3_LC_18_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_3_LC_18_12_2  (
            .in0(N__28258),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24480),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_1_LC_18_14_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_1_LC_18_14_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_1_LC_18_14_4.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_1_LC_18_14_4 (
            .in0(N__25474),
            .in1(N__24170),
            .in2(N__22456),
            .in3(N__22630),
            .lcout(M_this_sprites_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31953),
            .ce(),
            .sr(N__27291));
    defparam M_this_sprites_address_q_9_LC_18_14_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_9_LC_18_14_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_9_LC_18_14_7.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_9_LC_18_14_7 (
            .in0(N__24171),
            .in1(N__22447),
            .in2(N__22441),
            .in3(N__22831),
            .lcout(M_this_sprites_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31953),
            .ce(),
            .sr(N__27291));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_18_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_18_15_0 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_18_15_0  (
            .in0(N__22507),
            .in1(N__28170),
            .in2(N__34220),
            .in3(N__32639),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_2_LC_18_15_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_2_LC_18_15_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_2_LC_18_15_1.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_2_LC_18_15_1 (
            .in0(N__22426),
            .in1(N__24142),
            .in2(N__22429),
            .in3(N__22486),
            .lcout(M_this_sprites_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31957),
            .ce(),
            .sr(N__27290));
    defparam \this_vga_signals.M_this_sprites_address_q_m_2_LC_18_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_2_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_2_LC_18_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_2_LC_18_15_2  (
            .in0(N__22508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24465),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_3_LC_18_15_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_3_LC_18_15_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_3_LC_18_15_4.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_3_LC_18_15_4 (
            .in0(N__24143),
            .in1(N__28093),
            .in2(N__22420),
            .in3(N__22474),
            .lcout(M_this_sprites_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31957),
            .ce(),
            .sr(N__27290));
    defparam \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_16_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_16_0  (
            .in0(N__24859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24436),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_10_LC_18_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_10_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_10_LC_18_16_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_10_LC_18_16_1  (
            .in0(N__28163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22719),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIMJ231_8_LC_18_16_3.C_ON=1'b0;
    defparam M_this_state_q_RNIMJ231_8_LC_18_16_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIMJ231_8_LC_18_16_3.LUT_INIT=16'b1111111111101111;
    LogicCell40 M_this_state_q_RNIMJ231_8_LC_18_16_3 (
            .in0(N__25391),
            .in1(N__32923),
            .in2(N__31258),
            .in3(N__28031),
            .lcout(M_this_state_q_RNIMJ231Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_19_LC_18_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_19_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_19_LC_18_16_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_19_LC_18_16_4  (
            .in0(N__27940),
            .in1(N__25390),
            .in2(N__22663),
            .in3(N__24096),
            .lcout(\this_vga_signals.un1_M_this_state_q_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un23_i_a2_1_1_LC_18_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un23_i_a2_1_1_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un23_i_a2_1_1_LC_18_16_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.un23_i_a2_1_1_LC_18_16_6  (
            .in0(N__26400),
            .in1(N__31200),
            .in2(_gnd_net_),
            .in3(N__28162),
            .lcout(this_vga_signals_un23_i_a2_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNI1DGI7_0_LC_18_17_0.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNI1DGI7_0_LC_18_17_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNI1DGI7_0_LC_18_17_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNI1DGI7_0_LC_18_17_0 (
            .in0(_gnd_net_),
            .in1(N__25962),
            .in2(N__24097),
            .in3(N__24095),
            .lcout(M_this_sprites_address_q_RNI1DGI7Z0Z_0),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(un1_M_this_sprites_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_18_17_1.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_18_17_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_18_17_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_18_17_1 (
            .in0(_gnd_net_),
            .in1(N__25514),
            .in2(_gnd_net_),
            .in3(N__22621),
            .lcout(un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_0),
            .carryout(un1_M_this_sprites_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_18_17_2.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_18_17_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_18_17_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_18_17_2 (
            .in0(_gnd_net_),
            .in1(N__22515),
            .in2(_gnd_net_),
            .in3(N__22477),
            .lcout(un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_1),
            .carryout(un1_M_this_sprites_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_18_17_3.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_18_17_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_18_17_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_18_17_3 (
            .in0(_gnd_net_),
            .in1(N__28262),
            .in2(_gnd_net_),
            .in3(N__22465),
            .lcout(un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_2),
            .carryout(un1_M_this_sprites_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_18_17_4.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_18_17_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_18_17_4.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_18_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26166),
            .in3(N__22462),
            .lcout(un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_3),
            .carryout(un1_M_this_sprites_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_18_17_5.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_18_17_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_18_17_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_18_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24873),
            .in3(N__22459),
            .lcout(un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_4),
            .carryout(un1_M_this_sprites_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_18_17_6.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_18_17_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_18_17_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_18_17_6 (
            .in0(_gnd_net_),
            .in1(N__23711),
            .in2(_gnd_net_),
            .in3(N__23119),
            .lcout(un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_5),
            .carryout(un1_M_this_sprites_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_18_17_7.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_18_17_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_18_17_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_18_17_7 (
            .in0(_gnd_net_),
            .in1(N__24240),
            .in2(_gnd_net_),
            .in3(N__23116),
            .lcout(un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_6),
            .carryout(un1_M_this_sprites_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_18_18_0.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_18_18_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_18_18_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_18_18_0 (
            .in0(_gnd_net_),
            .in1(N__23010),
            .in2(_gnd_net_),
            .in3(N__22969),
            .lcout(un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(un1_M_this_sprites_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_18_18_1.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_18_18_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_18_18_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_18_18_1 (
            .in0(_gnd_net_),
            .in1(N__22860),
            .in2(_gnd_net_),
            .in3(N__22822),
            .lcout(un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_8),
            .carryout(un1_M_this_sprites_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_18_18_2.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_18_18_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_18_18_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_18_18_2 (
            .in0(_gnd_net_),
            .in1(N__22708),
            .in2(_gnd_net_),
            .in3(N__22675),
            .lcout(un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_9),
            .carryout(un1_M_this_sprites_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_18_18_3.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_18_18_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_18_18_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_18_18_3 (
            .in0(_gnd_net_),
            .in1(N__24523),
            .in2(_gnd_net_),
            .in3(N__22672),
            .lcout(un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_10),
            .carryout(un1_M_this_sprites_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_18_18_4.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_18_18_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_18_18_4.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_18_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25683),
            .in3(N__22669),
            .lcout(un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_11),
            .carryout(un1_M_this_sprites_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_18_18_5.C_ON=1'b0;
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_18_18_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_18_18_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_18_18_5 (
            .in0(_gnd_net_),
            .in1(N__23293),
            .in2(_gnd_net_),
            .in3(N__22666),
            .lcout(un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_0_0_0_0_LC_18_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_0_0_0_0_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_0_0_0_0_LC_18_18_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o2_0_0_0_0_LC_18_18_7  (
            .in0(N__32925),
            .in1(N__29595),
            .in2(_gnd_net_),
            .in3(N__24419),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_o2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_11_LC_18_19_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_11_LC_18_19_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_11_LC_18_19_1.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_11_LC_18_19_1 (
            .in0(N__24487),
            .in1(N__24172),
            .in2(N__24607),
            .in3(N__23392),
            .lcout(M_this_sprites_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31983),
            .ce(),
            .sr(N__27287));
    defparam M_this_sprites_address_q_12_LC_18_19_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_12_LC_18_19_3.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_12_LC_18_19_3.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_12_LC_18_19_3 (
            .in0(N__23386),
            .in1(N__24173),
            .in2(N__25633),
            .in3(N__23380),
            .lcout(M_this_sprites_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31983),
            .ce(),
            .sr(N__27287));
    defparam M_this_sprites_address_q_13_LC_18_19_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_13_LC_18_19_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_13_LC_18_19_4.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_13_LC_18_19_4 (
            .in0(N__24174),
            .in1(N__23374),
            .in2(N__23368),
            .in3(N__23356),
            .lcout(M_this_sprites_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31983),
            .ce(),
            .sr(N__27287));
    defparam \this_vga_signals.M_this_map_address_q_m_9_LC_18_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_9_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_9_LC_18_20_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_9_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__25218),
            .in2(_gnd_net_),
            .in3(N__27611),
            .lcout(\this_vga_signals.M_this_map_address_q_mZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_0_1_0_LC_18_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_0_1_0_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_0_1_0_LC_18_20_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o2_0_1_0_LC_18_20_4  (
            .in0(N__26436),
            .in1(N__25396),
            .in2(N__27625),
            .in3(N__28207),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_ns_0_o2_0_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_LC_18_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_LC_18_20_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_LC_18_20_5  (
            .in0(N__23236),
            .in1(N__27960),
            .in2(N__23227),
            .in3(N__32849),
            .lcout(N_435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_0_LC_18_21_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_0_LC_18_21_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_0_LC_18_21_4.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_0_LC_18_21_4 (
            .in0(N__25924),
            .in1(N__24181),
            .in2(N__23671),
            .in3(N__23224),
            .lcout(M_this_sprites_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31996),
            .ce(),
            .sr(N__27283));
    defparam \this_sprites_ram.mem_radreg_11_LC_18_22_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_11_LC_18_22_6 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_11_LC_18_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_sprites_ram.mem_radreg_11_LC_18_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23215),
            .lcout(\this_sprites_ram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32003),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_d_5_m_9_LC_18_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_5_m_9_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_5_m_9_LC_18_22_7 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_5_m_9_LC_18_22_7  (
            .in0(N__25210),
            .in1(N__26464),
            .in2(N__33311),
            .in3(N__32850),
            .lcout(\this_vga_signals.M_this_map_address_d_5_mZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_7_LC_18_23_1.C_ON=1'b0;
    defparam M_this_map_address_q_7_LC_18_23_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_7_LC_18_23_1.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_map_address_q_7_LC_18_23_1 (
            .in0(N__26325),
            .in1(N__25177),
            .in2(N__25129),
            .in3(N__25246),
            .lcout(M_this_map_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32010),
            .ce(),
            .sr(N__27281));
    defparam \this_vga_signals.M_this_map_address_q_m_2_LC_18_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_2_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_2_LC_18_23_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_2_LC_18_23_3  (
            .in0(N__24786),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26471),
            .lcout(),
            .ltout(\this_vga_signals.M_this_map_address_q_mZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_2_LC_18_23_4.C_ON=1'b0;
    defparam M_this_map_address_q_2_LC_18_23_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_2_LC_18_23_4.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_map_address_q_2_LC_18_23_4 (
            .in0(N__23623),
            .in1(N__26324),
            .in2(N__23626),
            .in3(N__24763),
            .lcout(M_this_map_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32010),
            .ce(),
            .sr(N__27281));
    defparam \this_vga_signals.M_this_map_address_d_8_m_2_LC_18_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_8_m_2_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_8_m_2_LC_18_23_5 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_8_m_2_LC_18_23_5  (
            .in0(N__24785),
            .in1(N__27626),
            .in2(N__34222),
            .in3(N__32848),
            .lcout(\this_vga_signals.M_this_map_address_d_8_mZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_9_LC_18_23_7.C_ON=1'b0;
    defparam M_this_map_address_q_9_LC_18_23_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_9_LC_18_23_7.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_map_address_q_9_LC_18_23_7 (
            .in0(N__26326),
            .in1(N__23617),
            .in2(N__23605),
            .in3(N__25183),
            .lcout(M_this_map_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32010),
            .ce(),
            .sr(N__27281));
    defparam \this_ppu.M_haddress_q_RNIR3M06_4_LC_18_25_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIR3M06_4_LC_18_25_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIR3M06_4_LC_18_25_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNIR3M06_4_LC_18_25_4  (
            .in0(N__23569),
            .in1(N__23919),
            .in2(N__23438),
            .in3(N__23975),
            .lcout(\this_ppu.un1_M_haddress_q_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_5_LC_18_26_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_5_LC_18_26_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_5_LC_18_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_haddress_q_5_LC_18_26_2  (
            .in0(_gnd_net_),
            .in1(N__25080),
            .in2(_gnd_net_),
            .in3(N__25049),
            .lcout(M_this_ppu_map_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32033),
            .ce(),
            .sr(N__25034));
    defparam \this_ppu.M_haddress_q_6_LC_18_26_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_6_LC_18_26_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_6_LC_18_26_3 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_ppu.M_haddress_q_6_LC_18_26_3  (
            .in0(N__25050),
            .in1(_gnd_net_),
            .in2(N__25093),
            .in3(N__33115),
            .lcout(M_this_ppu_vram_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32033),
            .ce(),
            .sr(N__25034));
    defparam \this_ppu.M_haddress_q_4_LC_18_26_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_4_LC_18_26_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_4_LC_18_26_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \this_ppu.M_haddress_q_4_LC_18_26_5  (
            .in0(N__23983),
            .in1(N__23426),
            .in2(N__23930),
            .in3(N__23570),
            .lcout(M_this_ppu_map_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32033),
            .ce(),
            .sr(N__25034));
    defparam \this_ppu.M_haddress_q_3_LC_18_26_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_3_LC_18_26_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_3_LC_18_26_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_haddress_q_3_LC_18_26_6  (
            .in0(N__23427),
            .in1(N__23920),
            .in2(_gnd_net_),
            .in3(N__23982),
            .lcout(M_this_ppu_map_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32033),
            .ce(),
            .sr(N__25034));
    defparam \this_ppu.M_vaddress_q_RNI0655_6_LC_18_29_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI0655_6_LC_18_29_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI0655_6_LC_18_29_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.M_vaddress_q_RNI0655_6_LC_18_29_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23893),
            .lcout(this_ppu_M_vaddress_q_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_19_14_6.C_ON=1'b0;
    defparam M_this_state_q_6_LC_19_14_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_19_14_6.LUT_INIT=16'b1010000011101100;
    LogicCell40 M_this_state_q_6_LC_19_14_6 (
            .in0(N__24595),
            .in1(N__30754),
            .in2(N__23638),
            .in3(N__32624),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31958),
            .ce(),
            .sr(N__32386));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_19_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_19_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_19_15_0 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_19_15_0  (
            .in0(N__23695),
            .in1(N__28220),
            .in2(N__33536),
            .in3(N__32620),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_6_LC_19_15_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_6_LC_19_15_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_6_LC_19_15_1.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_6_LC_19_15_1 (
            .in0(N__24150),
            .in1(N__23836),
            .in2(N__23824),
            .in3(N__23821),
            .lcout(M_this_sprites_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31965),
            .ce(),
            .sr(N__27292));
    defparam \this_vga_signals.M_this_sprites_address_q_m_0_LC_19_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_0_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_0_LC_19_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_0_LC_19_15_4  (
            .in0(_gnd_net_),
            .in1(N__25961),
            .in2(_gnd_net_),
            .in3(N__24475),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_5_LC_19_15_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_5_LC_19_15_6.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_5_LC_19_15_6.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_5_LC_19_15_6 (
            .in0(N__24835),
            .in1(N__24149),
            .in2(N__23656),
            .in3(N__23647),
            .lcout(M_this_sprites_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31965),
            .ce(),
            .sr(N__27292));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_6_LC_19_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_6_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_6_LC_19_16_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_0_6_LC_19_16_2  (
            .in0(N__26978),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26890),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_a2_0_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_6_0_a2_LC_19_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_a2_LC_19_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_a2_LC_19_16_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_6_0_a2_LC_19_16_3  (
            .in0(N__28199),
            .in1(N__24468),
            .in2(N__25381),
            .in3(N__25424),
            .lcout(),
            .ltout(\this_vga_signals.N_294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_14_1_LC_19_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_14_1_LC_19_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_14_1_LC_19_16_4 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_14_1_LC_19_16_4  (
            .in0(N__34058),
            .in1(N__32588),
            .in2(N__24103),
            .in3(N__29181),
            .lcout(),
            .ltout(\this_vga_signals.un1_M_this_state_q_14Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_14_LC_19_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_14_LC_19_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_14_LC_19_16_5 .LUT_INIT=16'b1010000010110000;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_14_LC_19_16_5  (
            .in0(N__32589),
            .in1(N__27231),
            .in2(N__24100),
            .in3(N__25379),
            .lcout(un1_M_this_state_q_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un23_i_a2_1_LC_19_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un23_i_a2_1_LC_19_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un23_i_a2_1_LC_19_16_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_vga_signals.un23_i_a2_1_LC_19_16_6  (
            .in0(N__25423),
            .in1(N__24072),
            .in2(N__29606),
            .in3(N__30756),
            .lcout(un23_i_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_3_LC_19_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_3_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_3_LC_19_17_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a3_3_LC_19_17_3  (
            .in0(N__26733),
            .in1(N__26791),
            .in2(N__25903),
            .in3(N__25811),
            .lcout(\this_vga_signals.N_486 ),
            .ltout(\this_vga_signals.N_486_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_19_17_4.C_ON=1'b0;
    defparam M_this_state_q_7_LC_19_17_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_19_17_4.LUT_INIT=16'b1010000011101100;
    LogicCell40 M_this_state_q_7_LC_19_17_4 (
            .in0(N__24043),
            .in1(N__29596),
            .in2(N__24019),
            .in3(N__32825),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31977),
            .ce(),
            .sr(N__32375));
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_19_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_19_17_5 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_19_17_5  (
            .in0(N__26732),
            .in1(N__26974),
            .in2(N__28578),
            .in3(N__26790),
            .lcout(N_465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_1_9_LC_19_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_1_9_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_1_9_LC_19_17_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_1_9_LC_19_17_7  (
            .in0(N__26734),
            .in1(N__26878),
            .in2(N__26991),
            .in3(N__26792),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_1_LC_19_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_1_LC_19_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_1_LC_19_18_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_1_1_LC_19_18_0  (
            .in0(N__26786),
            .in1(N__25898),
            .in2(N__24640),
            .in3(N__25812),
            .lcout(\this_vga_signals.N_438_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_i_o2_0_14_LC_19_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_i_o2_0_14_LC_19_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_i_o2_0_14_LC_19_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_i_o2_0_14_LC_19_18_1  (
            .in0(_gnd_net_),
            .in1(N__28078),
            .in2(_gnd_net_),
            .in3(N__31319),
            .lcout(this_vga_signals_M_this_state_q_ns_i_o2_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_i_o2_0_12_LC_19_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_i_o2_0_12_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_i_o2_0_12_LC_19_18_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_i_o2_0_12_LC_19_18_2  (
            .in0(N__28077),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31201),
            .lcout(this_vga_signals_M_this_state_q_ns_i_o2_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_11_LC_19_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_11_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_11_LC_19_18_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_11_LC_19_18_5  (
            .in0(N__24525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28226),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_5_LC_19_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_5_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_5_LC_19_18_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_1_5_LC_19_18_7  (
            .in0(N__25813),
            .in1(N__26716),
            .in2(N__26796),
            .in3(N__25902),
            .lcout(\this_vga_signals.N_446_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_19_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_19_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_19_19_0 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_19_19_0  (
            .in0(N__24524),
            .in1(N__24476),
            .in2(N__33336),
            .in3(N__32822),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_19_2 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_19_2  (
            .in0(N__24232),
            .in1(N__33794),
            .in2(N__24481),
            .in3(N__32823),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_7_LC_19_19_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_7_LC_19_19_3.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_7_LC_19_19_3.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_7_LC_19_19_3 (
            .in0(N__24180),
            .in1(N__24211),
            .in2(N__24352),
            .in3(N__24349),
            .lcout(M_this_sprites_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31990),
            .ce(),
            .sr(N__27288));
    defparam \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_19_4  (
            .in0(N__24233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28227),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_4_LC_19_19_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_4_LC_19_19_6.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_4_LC_19_19_6.LUT_INIT=16'b1111101011111110;
    LogicCell40 M_this_sprites_address_q_4_LC_19_19_6 (
            .in0(N__26125),
            .in1(N__24205),
            .in2(N__24196),
            .in3(N__24179),
            .lcout(M_this_sprites_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31990),
            .ce(),
            .sr(N__27288));
    defparam \this_vga_signals.M_this_map_address_d_5_m_5_LC_19_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_5_m_5_LC_19_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_5_m_5_LC_19_20_1 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_5_m_5_LC_19_20_1  (
            .in0(N__24731),
            .in1(N__26462),
            .in2(N__33841),
            .in3(N__32755),
            .lcout(\this_vga_signals.M_this_map_address_d_5_mZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_q_m_0_LC_19_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_0_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_0_LC_19_20_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_0_LC_19_20_2  (
            .in0(N__26463),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26096),
            .lcout(\this_vga_signals.M_this_map_address_q_mZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d_1_sqmuxa_LC_19_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d_1_sqmuxa_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d_1_sqmuxa_LC_19_20_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_this_state_d_1_sqmuxa_LC_19_20_3  (
            .in0(N__33692),
            .in1(N__32754),
            .in2(_gnd_net_),
            .in3(N__29190),
            .lcout(\this_vga_signals.M_this_state_d_1_sqmuxaZ0 ),
            .ltout(\this_vga_signals.M_this_state_d_1_sqmuxaZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_12_LC_19_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_12_LC_19_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_12_LC_19_20_4 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_12_LC_19_20_4  (
            .in0(N__29191),
            .in1(N__25915),
            .in2(N__24643),
            .in3(N__27871),
            .lcout(un1_M_this_state_q_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_19_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_19_20_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_19_20_5  (
            .in0(N__26953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26715),
            .lcout(\this_vga_signals.N_399_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_8_0_a2_1_LC_19_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_8_0_a2_1_LC_19_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_8_0_a2_1_LC_19_20_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_8_0_a2_1_LC_19_20_6  (
            .in0(_gnd_net_),
            .in1(N__30755),
            .in2(_gnd_net_),
            .in3(N__30636),
            .lcout(\this_vga_signals.N_293_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_q_m_6_LC_19_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_6_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_6_LC_19_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_6_LC_19_20_7  (
            .in0(N__24677),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27627),
            .lcout(\this_vga_signals.M_this_map_address_q_mZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_q_m_5_LC_19_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_5_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_5_LC_19_21_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_5_LC_19_21_0  (
            .in0(_gnd_net_),
            .in1(N__24732),
            .in2(_gnd_net_),
            .in3(N__27624),
            .lcout(),
            .ltout(\this_vga_signals.M_this_map_address_q_mZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_5_LC_19_21_1.C_ON=1'b0;
    defparam M_this_map_address_q_5_LC_19_21_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_5_LC_19_21_1.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_map_address_q_5_LC_19_21_1 (
            .in0(N__26328),
            .in1(N__24625),
            .in2(N__24619),
            .in3(N__24706),
            .lcout(M_this_map_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32004),
            .ce(),
            .sr(N__27285));
    defparam M_this_map_address_q_0_LC_19_21_4.C_ON=1'b0;
    defparam M_this_map_address_q_0_LC_19_21_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_0_LC_19_21_4.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_map_address_q_0_LC_19_21_4 (
            .in0(N__26068),
            .in1(N__26327),
            .in2(N__24616),
            .in3(N__24817),
            .lcout(M_this_map_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32004),
            .ce(),
            .sr(N__27285));
    defparam \this_vga_signals.M_this_map_address_d_5_m_6_LC_19_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_5_m_6_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_5_m_6_LC_19_21_6 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_5_m_6_LC_19_21_6  (
            .in0(N__24678),
            .in1(N__26474),
            .in2(N__33990),
            .in3(N__32824),
            .lcout(),
            .ltout(\this_vga_signals.M_this_map_address_d_5_mZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_6_LC_19_21_7.C_ON=1'b0;
    defparam M_this_map_address_q_6_LC_19_21_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_6_LC_19_21_7.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_map_address_q_6_LC_19_21_7 (
            .in0(N__26329),
            .in1(N__24829),
            .in2(N__24820),
            .in3(N__24652),
            .lcout(M_this_map_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32004),
            .ce(),
            .sr(N__27285));
    defparam M_this_map_address_q_RNICF7V6_0_LC_19_22_0.C_ON=1'b1;
    defparam M_this_map_address_q_RNICF7V6_0_LC_19_22_0.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNICF7V6_0_LC_19_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_RNICF7V6_0_LC_19_22_0 (
            .in0(_gnd_net_),
            .in1(N__26092),
            .in2(N__26362),
            .in3(N__26360),
            .lcout(M_this_map_address_q_RNICF7V6Z0Z_0),
            .ltout(),
            .carryin(bfn_19_22_0_),
            .carryout(un1_M_this_map_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_0_c_RNI6GRR_LC_19_22_1.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_0_c_RNI6GRR_LC_19_22_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_0_c_RNI6GRR_LC_19_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_map_address_q_cry_0_c_RNI6GRR_LC_19_22_1 (
            .in0(_gnd_net_),
            .in1(N__26626),
            .in2(_gnd_net_),
            .in3(N__24811),
            .lcout(un1_M_this_map_address_q_cry_0_c_RNI6GRRZ0),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_0),
            .carryout(un1_M_this_map_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_1_c_RNI8JSR_LC_19_22_2.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_1_c_RNI8JSR_LC_19_22_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_1_c_RNI8JSR_LC_19_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_map_address_q_cry_1_c_RNI8JSR_LC_19_22_2 (
            .in0(_gnd_net_),
            .in1(N__24784),
            .in2(_gnd_net_),
            .in3(N__24757),
            .lcout(un1_M_this_map_address_q_cry_1_c_RNI8JSRZ0),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_1),
            .carryout(un1_M_this_map_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_2_c_RNIAMTR_LC_19_22_3.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_2_c_RNIAMTR_LC_19_22_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_2_c_RNIAMTR_LC_19_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_map_address_q_cry_2_c_RNIAMTR_LC_19_22_3 (
            .in0(_gnd_net_),
            .in1(N__26572),
            .in2(_gnd_net_),
            .in3(N__24754),
            .lcout(un1_M_this_map_address_q_cry_2_c_RNIAMTRZ0),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_2),
            .carryout(un1_M_this_map_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_3_c_RNICPUR_LC_19_22_4.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_3_c_RNICPUR_LC_19_22_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_3_c_RNICPUR_LC_19_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_map_address_q_cry_3_c_RNICPUR_LC_19_22_4 (
            .in0(_gnd_net_),
            .in1(N__26497),
            .in2(_gnd_net_),
            .in3(N__24751),
            .lcout(un1_M_this_map_address_q_cry_3_c_RNICPURZ0),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_3),
            .carryout(un1_M_this_map_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_4_c_RNIESVR_LC_19_22_5.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_4_c_RNIESVR_LC_19_22_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_4_c_RNIESVR_LC_19_22_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_map_address_q_cry_4_c_RNIESVR_LC_19_22_5 (
            .in0(_gnd_net_),
            .in1(N__24730),
            .in2(_gnd_net_),
            .in3(N__24700),
            .lcout(un1_M_this_map_address_q_cry_4_c_RNIESVRZ0),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_4),
            .carryout(un1_M_this_map_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_5_c_RNIGV0S_LC_19_22_6.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_5_c_RNIGV0S_LC_19_22_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_5_c_RNIGV0S_LC_19_22_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_map_address_q_cry_5_c_RNIGV0S_LC_19_22_6 (
            .in0(_gnd_net_),
            .in1(N__24676),
            .in2(_gnd_net_),
            .in3(N__24646),
            .lcout(un1_M_this_map_address_q_cry_5_c_RNIGV0SZ0),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_5),
            .carryout(un1_M_this_map_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_6_c_RNII22S_LC_19_22_7.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_6_c_RNII22S_LC_19_22_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_6_c_RNII22S_LC_19_22_7.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_map_address_q_cry_6_c_RNII22S_LC_19_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25161),
            .in3(N__25240),
            .lcout(un1_M_this_map_address_q_cry_6_c_RNII22SZ0),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_6),
            .carryout(un1_M_this_map_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_7_c_RNIK53S_LC_19_23_0.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_7_c_RNIK53S_LC_19_23_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_7_c_RNIK53S_LC_19_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_map_address_q_cry_7_c_RNIK53S_LC_19_23_0 (
            .in0(_gnd_net_),
            .in1(N__27655),
            .in2(_gnd_net_),
            .in3(N__25237),
            .lcout(un1_M_this_map_address_q_cry_7_c_RNIK53SZ0),
            .ltout(),
            .carryin(bfn_19_23_0_),
            .carryout(un1_M_this_map_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_8_c_RNIM84S_LC_19_23_1.C_ON=1'b0;
    defparam un1_M_this_map_address_q_cry_8_c_RNIM84S_LC_19_23_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_8_c_RNIM84S_LC_19_23_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_M_this_map_address_q_cry_8_c_RNIM84S_LC_19_23_1 (
            .in0(_gnd_net_),
            .in1(N__25214),
            .in2(_gnd_net_),
            .in3(N__25186),
            .lcout(un1_M_this_map_address_q_cry_8_c_RNIM84SZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_d_5_m_7_LC_19_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_5_m_7_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_5_m_7_LC_19_23_2 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_5_m_7_LC_19_23_2  (
            .in0(N__32821),
            .in1(N__25156),
            .in2(N__34221),
            .in3(N__26475),
            .lcout(\this_vga_signals.M_this_map_address_d_5_mZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_q_m_7_LC_19_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_7_LC_19_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_7_LC_19_24_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_7_LC_19_24_2  (
            .in0(_gnd_net_),
            .in1(N__25157),
            .in2(_gnd_net_),
            .in3(N__27623),
            .lcout(\this_vga_signals.M_this_map_address_q_mZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_7_LC_19_26_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_7_LC_19_26_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_7_LC_19_26_6 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_ppu.M_haddress_q_7_LC_19_26_6  (
            .in0(N__33174),
            .in1(N__33116),
            .in2(N__25097),
            .in3(N__25051),
            .lcout(\this_ppu.M_haddress_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32039),
            .ce(),
            .sr(N__25035));
    defparam \this_reset_cond.M_stage_q_7_LC_20_14_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_7_LC_20_14_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_7_LC_20_14_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_7_LC_20_14_4  (
            .in0(N__28483),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24991),
            .lcout(\this_reset_cond.M_stage_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31966),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_20_14_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_20_14_6 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_20_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_20_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24982),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31966),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_20_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_20_15_2 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_20_15_2  (
            .in0(N__24866),
            .in1(N__28213),
            .in2(N__33646),
            .in3(N__32746),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_12_LC_20_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_12_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_12_LC_20_15_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_i_o3_0_12_LC_20_15_4  (
            .in0(N__27030),
            .in1(N__27119),
            .in2(_gnd_net_),
            .in3(N__27160),
            .lcout(\this_vga_signals.N_390_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_20_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_20_15_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_20_15_5  (
            .in0(N__27118),
            .in1(N__27158),
            .in2(_gnd_net_),
            .in3(N__27029),
            .lcout(N_389_0),
            .ltout(N_389_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_20_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_20_15_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_20_15_6  (
            .in0(N__33999),
            .in1(N__25518),
            .in2(N__25477),
            .in3(N__28212),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_8_LC_20_16_2.C_ON=1'b0;
    defparam M_this_state_q_8_LC_20_16_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_8_LC_20_16_2.LUT_INIT=16'b1100000011101010;
    LogicCell40 M_this_state_q_8_LC_20_16_2 (
            .in0(N__32916),
            .in1(N__25782),
            .in2(N__26995),
            .in3(N__32622),
            .lcout(M_this_state_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31978),
            .ce(),
            .sr(N__32376));
    defparam \this_vga_signals.un23_i_a2_0_1_LC_20_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un23_i_a2_0_1_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un23_i_a2_0_1_LC_20_16_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.un23_i_a2_0_1_LC_20_16_3  (
            .in0(N__29160),
            .in1(N__25462),
            .in2(_gnd_net_),
            .in3(N__25746),
            .lcout(N_297),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_9_LC_20_16_7.C_ON=1'b0;
    defparam M_this_state_q_9_LC_20_16_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_9_LC_20_16_7.LUT_INIT=16'b1101010111000000;
    LogicCell40 M_this_state_q_9_LC_20_16_7 (
            .in0(N__32621),
            .in1(N__27246),
            .in2(N__25405),
            .in3(N__25380),
            .lcout(M_this_state_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31978),
            .ce(),
            .sr(N__32376));
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_sx_9_LC_20_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_sx_9_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_sx_9_LC_20_17_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a3_sx_9_LC_20_17_0  (
            .in0(N__25332),
            .in1(N__28574),
            .in2(N__25269),
            .in3(N__28076),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_ns_0_a3_sxZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_9_LC_20_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_9_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_9_LC_20_17_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a3_9_LC_20_17_1  (
            .in0(N__25881),
            .in1(N__25839),
            .in2(N__25336),
            .in3(N__25308),
            .lcout(\this_vga_signals.N_469 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_8_3_0_LC_20_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_8_3_0_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_8_3_0_LC_20_17_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o3_8_3_0_LC_20_17_2  (
            .in0(N__25333),
            .in1(N__25309),
            .in2(N__25270),
            .in3(N__28075),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_o3_8_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_5_0_a2_LC_20_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_5_0_a2_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_5_0_a2_LC_20_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_5_0_a2_LC_20_17_4  (
            .in0(N__28036),
            .in1(N__26426),
            .in2(N__27622),
            .in3(N__29162),
            .lcout(\this_vga_signals.N_291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_1_0_LC_20_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_1_0_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_1_0_LC_20_18_0 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a3_1_0_LC_20_18_0  (
            .in0(N__25810),
            .in1(N__25852),
            .in2(N__25882),
            .in3(N__28561),
            .lcout(N_466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_1_LC_20_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_1_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_1_LC_20_18_2 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_1_LC_20_18_2  (
            .in0(N__25876),
            .in1(N__25850),
            .in2(_gnd_net_),
            .in3(N__28559),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_4_LC_20_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_4_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_4_LC_20_18_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_1_sx_4_LC_20_18_4  (
            .in0(N__25877),
            .in1(N__25851),
            .in2(N__26889),
            .in3(N__28560),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_ns_0_a2_0_1_sxZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_4_LC_20_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_4_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_1_4_LC_20_18_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_1_4_LC_20_18_5  (
            .in0(N__26717),
            .in1(N__26769),
            .in2(N__25816),
            .in3(N__25809),
            .lcout(\this_vga_signals.N_444_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_14_LC_20_19_0.C_ON=1'b0;
    defparam M_this_external_address_q_14_LC_20_19_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_14_LC_20_19_0.LUT_INIT=16'b1111011111110101;
    LogicCell40 M_this_external_address_q_14_LC_20_19_0 (
            .in0(N__26269),
            .in1(N__30470),
            .in2(N__27330),
            .in3(N__28804),
            .lcout(M_this_external_address_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31997),
            .ce(),
            .sr(N__32380));
    defparam \this_vga_signals.M_this_external_address_d_5_14_LC_20_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_5_14_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_5_14_LC_20_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_this_external_address_d_5_14_LC_20_19_2  (
            .in0(N__33537),
            .in1(N__28825),
            .in2(_gnd_net_),
            .in3(N__32756),
            .lcout(\this_vga_signals.M_this_external_address_d_5Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_fast_14_LC_20_19_3.C_ON=1'b0;
    defparam M_this_state_q_fast_14_LC_20_19_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_fast_14_LC_20_19_3.LUT_INIT=16'b0101010100010000;
    LogicCell40 M_this_state_q_fast_14_LC_20_19_3 (
            .in0(N__32757),
            .in1(N__28523),
            .in2(N__25764),
            .in3(N__25747),
            .lcout(M_this_state_q_fastZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31997),
            .ce(),
            .sr(N__32380));
    defparam \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_20_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25724),
            .in3(N__28203),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d_0_sqmuxa_1_LC_20_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d_0_sqmuxa_1_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d_0_sqmuxa_1_LC_20_20_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_this_state_d_0_sqmuxa_1_LC_20_20_2  (
            .in0(N__34057),
            .in1(N__32770),
            .in2(_gnd_net_),
            .in3(N__29188),
            .lcout(\this_vga_signals.M_this_state_d_0_sqmuxaZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_3_iv_0_14_LC_20_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_3_iv_0_14_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_3_iv_0_14_LC_20_20_3 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \this_vga_signals.M_this_external_address_q_3_iv_0_14_LC_20_20_3  (
            .in0(N__30843),
            .in1(N__26275),
            .in2(N__28838),
            .in3(N__30675),
            .lcout(\this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_20_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_20_20_4 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_20_20_4  (
            .in0(N__26152),
            .in1(N__33319),
            .in2(N__28222),
            .in3(N__32771),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_m_5_LC_20_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_5_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_5_LC_20_20_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_5_LC_20_20_5  (
            .in0(_gnd_net_),
            .in1(N__28744),
            .in2(_gnd_net_),
            .in3(N__30676),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_d_8_m_1_LC_20_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_8_m_1_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_8_m_1_LC_20_21_0 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_8_m_1_LC_20_21_0  (
            .in0(N__32759),
            .in1(N__26627),
            .in2(N__33991),
            .in3(N__27599),
            .lcout(\this_vga_signals.M_this_map_address_d_8_mZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_d_8_m_0_LC_20_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_8_m_0_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_8_m_0_LC_20_21_1 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_8_m_0_LC_20_21_1  (
            .in0(N__26100),
            .in1(N__27597),
            .in2(N__33836),
            .in3(N__32760),
            .lcout(\this_vga_signals.M_this_map_address_d_8_mZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_q_m_4_LC_20_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_4_LC_20_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_4_LC_20_21_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_4_LC_20_21_3  (
            .in0(N__26499),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26453),
            .lcout(\this_vga_signals.M_this_map_address_q_mZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_d_8_m_4_LC_20_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_8_m_4_LC_20_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_8_m_4_LC_20_21_5 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_8_m_4_LC_20_21_5  (
            .in0(N__26498),
            .in1(N__27598),
            .in2(N__33329),
            .in3(N__32761),
            .lcout(\this_vga_signals.M_this_map_address_d_8_mZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_6 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_6  (
            .in0(N__32758),
            .in1(N__25951),
            .in2(N__28228),
            .in3(N__33827),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_q_m_1_LC_20_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_1_LC_20_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_1_LC_20_22_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_1_LC_20_22_0  (
            .in0(N__26473),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26628),
            .lcout(),
            .ltout(\this_vga_signals.M_this_map_address_q_mZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_1_LC_20_22_1.C_ON=1'b0;
    defparam M_this_map_address_q_1_LC_20_22_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_1_LC_20_22_1.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_map_address_q_1_LC_20_22_1 (
            .in0(N__26662),
            .in1(N__26306),
            .in2(N__26656),
            .in3(N__26653),
            .lcout(M_this_map_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32019),
            .ce(),
            .sr(N__27286));
    defparam \this_vga_signals.M_this_map_address_d_8_m_3_LC_20_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_8_m_3_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_8_m_3_LC_20_22_3 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_8_m_3_LC_20_22_3  (
            .in0(N__26574),
            .in1(N__27603),
            .in2(N__34362),
            .in3(N__32772),
            .lcout(),
            .ltout(\this_vga_signals.M_this_map_address_d_8_mZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_3_LC_20_22_4.C_ON=1'b0;
    defparam M_this_map_address_q_3_LC_20_22_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_3_LC_20_22_4.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_map_address_q_3_LC_20_22_4 (
            .in0(N__26307),
            .in1(N__26548),
            .in2(N__26602),
            .in3(N__26599),
            .lcout(M_this_map_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32019),
            .ce(),
            .sr(N__27286));
    defparam \this_vga_signals.M_this_map_address_q_m_3_LC_20_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_3_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_3_LC_20_22_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_3_LC_20_22_5  (
            .in0(_gnd_net_),
            .in1(N__26573),
            .in2(_gnd_net_),
            .in3(N__26472),
            .lcout(\this_vga_signals.M_this_map_address_q_mZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_4_LC_20_22_7.C_ON=1'b0;
    defparam M_this_map_address_q_4_LC_20_22_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_4_LC_20_22_7.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_map_address_q_4_LC_20_22_7 (
            .in0(N__26542),
            .in1(N__26308),
            .in2(N__26536),
            .in3(N__26524),
            .lcout(M_this_map_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32019),
            .ce(),
            .sr(N__27286));
    defparam \this_vga_signals.M_this_map_address_d_5_m_8_LC_20_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_d_5_m_8_LC_20_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_d_5_m_8_LC_20_23_1 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_map_address_d_5_m_8_LC_20_23_1  (
            .in0(N__27656),
            .in1(N__26476),
            .in2(N__34332),
            .in3(N__32854),
            .lcout(\this_vga_signals.M_this_map_address_d_5_mZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_map_ram_write_en_LC_20_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_map_ram_write_en_LC_20_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_map_ram_write_en_LC_20_23_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.un1_M_this_map_ram_write_en_LC_20_23_3  (
            .in0(_gnd_net_),
            .in1(N__33001),
            .in2(_gnd_net_),
            .in3(N__26361),
            .lcout(\this_vga_signals.un1_M_this_map_ram_write_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_8_LC_20_24_5.C_ON=1'b0;
    defparam M_this_map_address_q_8_LC_20_24_5.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_8_LC_20_24_5.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_map_address_q_8_LC_20_24_5 (
            .in0(N__26335),
            .in1(N__26309),
            .in2(N__27511),
            .in3(N__26281),
            .lcout(M_this_map_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32034),
            .ce(),
            .sr(N__27282));
    defparam M_this_state_q_10_LC_21_14_7.C_ON=1'b0;
    defparam M_this_state_q_10_LC_21_14_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_10_LC_21_14_7.LUT_INIT=16'b0011101100001010;
    LogicCell40 M_this_state_q_10_LC_21_14_7 (
            .in0(N__27250),
            .in1(N__32623),
            .in2(N__26674),
            .in3(N__29159),
            .lcout(M_this_state_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31968),
            .ce(),
            .sr(N__32381));
    defparam M_this_state_q_15_LC_21_15_4.C_ON=1'b0;
    defparam M_this_state_q_15_LC_21_15_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_15_LC_21_15_4.LUT_INIT=16'b0010001000100000;
    LogicCell40 M_this_state_q_15_LC_21_15_4 (
            .in0(N__27235),
            .in1(N__27167),
            .in2(N__27126),
            .in3(N__27042),
            .lcout(M_this_state_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31979),
            .ce(),
            .sr(N__32377));
    defparam \this_vga_signals.M_this_data_count_q_3_bm_10_LC_21_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_bm_10_LC_21_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_bm_10_LC_21_16_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_bm_10_LC_21_16_0  (
            .in0(N__32616),
            .in1(N__32432),
            .in2(N__33697),
            .in3(N__29163),
            .lcout(\this_vga_signals.M_this_data_count_q_3_bmZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_m_6_LC_21_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_6_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_6_LC_21_16_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_6_LC_21_16_2  (
            .in0(N__28698),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30683),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_tr37_LC_21_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_tr37_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_tr37_LC_21_16_6 .LUT_INIT=16'b1000100010001010;
    LogicCell40 \this_vga_signals.M_this_state_q_tr37_LC_21_16_6  (
            .in0(N__28035),
            .in1(N__27159),
            .in2(N__27098),
            .in3(N__27043),
            .lcout(\this_vga_signals.M_this_map_ram_write_data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_21_16_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_21_16_7 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_21_16_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_21_16_7  (
            .in0(N__27044),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27086),
            .lcout(this_start_data_delay_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31984),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_tr35_LC_21_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_tr35_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_tr35_LC_21_17_2 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_vga_signals.M_this_state_q_tr35_LC_21_17_2  (
            .in0(N__28041),
            .in1(N__27161),
            .in2(N__27127),
            .in3(N__27045),
            .lcout(M_this_map_ram_write_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_1_10_LC_21_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_1_10_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_1_10_LC_21_17_3 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_1_10_LC_21_17_3  (
            .in0(N__26947),
            .in1(N__26882),
            .in2(N__26800),
            .in3(N__26724),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_2_sqmuxa_LC_21_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_2_sqmuxa_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_2_sqmuxa_LC_21_17_7 .LUT_INIT=16'b0101011100000000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_2_sqmuxa_LC_21_17_7  (
            .in0(N__32625),
            .in1(N__33693),
            .in2(N__34063),
            .in3(N__29161),
            .lcout(\this_vga_signals.M_this_external_address_d_2_sqmuxaZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_5_13_LC_21_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_5_13_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_5_13_LC_21_18_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vga_signals.M_this_external_address_d_5_13_LC_21_18_1  (
            .in0(N__28876),
            .in1(N__33614),
            .in2(_gnd_net_),
            .in3(N__32637),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_d_5Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_3_iv_0_13_LC_21_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_3_iv_0_13_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_3_iv_0_13_LC_21_18_2 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \this_vga_signals.M_this_external_address_q_3_iv_0_13_LC_21_18_2  (
            .in0(N__30669),
            .in1(N__30800),
            .in2(N__27337),
            .in3(N__28877),
            .lcout(\this_vga_signals.M_this_external_address_q_3_iv_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_bm_13_LC_21_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_bm_13_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_bm_13_LC_21_19_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_bm_13_LC_21_19_0  (
            .in0(N__32750),
            .in1(N__32433),
            .in2(N__34050),
            .in3(N__29187),
            .lcout(\this_vga_signals.M_this_data_count_q_3_bmZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_13_LC_21_19_2.C_ON=1'b0;
    defparam M_this_state_q_13_LC_21_19_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_13_LC_21_19_2.LUT_INIT=16'b1111111011111010;
    LogicCell40 M_this_state_q_13_LC_21_19_2 (
            .in0(N__27936),
            .in1(N__31150),
            .in2(N__27313),
            .in3(N__31295),
            .lcout(M_this_state_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32005),
            .ce(),
            .sr(N__32378));
    defparam M_this_state_q_11_LC_21_19_4.C_ON=1'b0;
    defparam M_this_state_q_11_LC_21_19_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_11_LC_21_19_4.LUT_INIT=16'b1111111111101010;
    LogicCell40 M_this_state_q_11_LC_21_19_4 (
            .in0(N__27334),
            .in1(N__31149),
            .in2(N__31199),
            .in3(N__32985),
            .lcout(M_this_state_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32005),
            .ce(),
            .sr(N__32378));
    defparam \this_vga_signals.un1_M_this_state_q_21_LC_21_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_21_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_21_LC_21_19_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_21_LC_21_19_5  (
            .in0(N__32984),
            .in1(N__27935),
            .in2(_gnd_net_),
            .in3(N__28785),
            .lcout(\this_vga_signals.un1_M_this_state_q_21_0 ),
            .ltout(\this_vga_signals.un1_M_this_state_q_21_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_13_LC_21_19_6.C_ON=1'b0;
    defparam M_this_external_address_q_13_LC_21_19_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_13_LC_21_19_6.LUT_INIT=16'b1010111011111111;
    LogicCell40 M_this_external_address_q_13_LC_21_19_6 (
            .in0(N__27309),
            .in1(N__28861),
            .in2(N__27301),
            .in3(N__27298),
            .lcout(M_this_external_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32005),
            .ce(),
            .sr(N__32378));
    defparam \this_vga_signals.M_this_external_address_q_m_4_LC_21_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_4_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_4_LC_21_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_4_LC_21_20_1  (
            .in0(_gnd_net_),
            .in1(N__30685),
            .in2(_gnd_net_),
            .in3(N__30237),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_8_m_5_LC_21_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_8_m_5_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_8_m_5_LC_21_20_2 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_8_m_5_LC_21_20_2  (
            .in0(N__30841),
            .in1(N__33630),
            .in2(N__28749),
            .in3(N__32752),
            .lcout(\this_vga_signals.M_this_external_address_d_8_mZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_8_m_4_LC_21_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_8_m_4_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_8_m_4_LC_21_20_3 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_8_m_4_LC_21_20_3  (
            .in0(N__32751),
            .in1(N__30236),
            .in2(N__33328),
            .in3(N__30840),
            .lcout(\this_vga_signals.M_this_external_address_d_8_mZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_8_0_a2_LC_21_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_8_0_a2_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_8_0_a2_LC_21_20_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_8_0_a2_LC_21_20_5  (
            .in0(N__28042),
            .in1(N__27961),
            .in2(N__27944),
            .in3(N__29164),
            .lcout(),
            .ltout(\this_vga_signals.N_293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_16_LC_21_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_16_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_16_LC_21_20_6 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_16_LC_21_20_6  (
            .in0(_gnd_net_),
            .in1(N__27864),
            .in2(N__27847),
            .in3(N__29082),
            .lcout(un1_M_this_state_q_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_13_LC_21_20_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_13_LC_21_20_7 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_13_LC_21_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_sprites_ram.mem_radreg_13_LC_21_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27844),
            .lcout(\this_sprites_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32011),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_5_LC_21_21_1.C_ON=1'b0;
    defparam M_this_external_address_q_5_LC_21_21_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_5_LC_21_21_1.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_external_address_q_5_LC_21_21_1 (
            .in0(N__27703),
            .in1(N__30487),
            .in2(N__27697),
            .in3(N__28717),
            .lcout(M_this_external_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32020),
            .ce(),
            .sr(N__32383));
    defparam \this_vga_signals.M_this_external_address_d_8_m_6_LC_21_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_8_m_6_LC_21_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_8_m_6_LC_21_21_5 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_8_m_6_LC_21_21_5  (
            .in0(N__30842),
            .in1(N__28694),
            .in2(N__33532),
            .in3(N__32753),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_d_8_mZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_6_LC_21_21_6.C_ON=1'b0;
    defparam M_this_external_address_q_6_LC_21_21_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_6_LC_21_21_6.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_external_address_q_6_LC_21_21_6 (
            .in0(N__30488),
            .in1(N__27688),
            .in2(N__27679),
            .in3(N__28669),
            .lcout(M_this_external_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32020),
            .ce(),
            .sr(N__32383));
    defparam \this_vga_signals.M_this_map_address_q_m_8_LC_21_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_m_8_LC_21_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_m_8_LC_21_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_m_8_LC_21_23_3  (
            .in0(_gnd_net_),
            .in1(N__27657),
            .in2(_gnd_net_),
            .in3(N__27631),
            .lcout(\this_vga_signals.M_this_map_address_q_mZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_9_LC_22_13_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_9_LC_22_13_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_9_LC_22_13_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_9_LC_22_13_5  (
            .in0(_gnd_net_),
            .in1(N__28466),
            .in2(_gnd_net_),
            .in3(N__28372),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31969),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_8_LC_22_13_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_8_LC_22_13_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_8_LC_22_13_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_8_LC_22_13_7  (
            .in0(_gnd_net_),
            .in1(N__28465),
            .in2(_gnd_net_),
            .in3(N__28384),
            .lcout(\this_reset_cond.M_stage_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31969),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_22_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_22_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_22_14_3 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_22_14_3  (
            .in0(N__28266),
            .in1(N__28221),
            .in2(N__34363),
            .in3(N__32773),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIV6TA_2_LC_22_15_0.C_ON=1'b0;
    defparam M_this_data_count_q_RNIV6TA_2_LC_22_15_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIV6TA_2_LC_22_15_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 M_this_data_count_q_RNIV6TA_2_LC_22_15_0 (
            .in0(_gnd_net_),
            .in1(N__29537),
            .in2(_gnd_net_),
            .in3(N__29321),
            .lcout(),
            .ltout(M_this_state_d88_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNI44LB1_0_LC_22_15_1.C_ON=1'b0;
    defparam M_this_data_count_q_RNI44LB1_0_LC_22_15_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNI44LB1_0_LC_22_15_1.LUT_INIT=16'b0001000000000000;
    LogicCell40 M_this_data_count_q_RNI44LB1_0_LC_22_15_1 (
            .in0(N__29356),
            .in1(N__29377),
            .in2(N__28081),
            .in3(N__29065),
            .lcout(M_this_state_d88_12),
            .ltout(M_this_state_d88_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d_1_sqmuxa_1_LC_22_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d_1_sqmuxa_1_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d_1_sqmuxa_1_LC_22_15_2 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \this_vga_signals.M_this_state_d_1_sqmuxa_1_LC_22_15_2  (
            .in0(N__28654),
            .in1(N__28074),
            .in2(N__28048),
            .in3(N__31567),
            .lcout(\this_vga_signals.N_387_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_m_7_LC_22_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_7_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_7_LC_22_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_7_LC_22_15_6  (
            .in0(_gnd_net_),
            .in1(N__30978),
            .in2(_gnd_net_),
            .in3(N__30682),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_22_16_0.C_ON=1'b0;
    defparam M_this_data_count_q_0_LC_22_16_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_22_16_0.LUT_INIT=16'b0101000011001100;
    LogicCell40 M_this_data_count_q_0_LC_22_16_0 (
            .in0(N__32252),
            .in1(N__29203),
            .in2(N__29059),
            .in3(N__32154),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31991),
            .ce(N__31676),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_1_LC_22_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_1_LC_22_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_1_LC_22_16_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_1_LC_22_16_3  (
            .in0(N__33989),
            .in1(N__31116),
            .in2(_gnd_net_),
            .in3(N__29355),
            .lcout(),
            .ltout(N_507_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_1_LC_22_16_4.C_ON=1'b0;
    defparam M_this_data_count_q_1_LC_22_16_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_22_16_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 M_this_data_count_q_1_LC_22_16_4 (
            .in0(N__32253),
            .in1(N__29335),
            .in2(N__28045),
            .in3(N__32155),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31991),
            .ce(N__31676),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_2_LC_22_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_2_LC_22_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_2_LC_22_16_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_2_LC_22_16_5  (
            .in0(N__34192),
            .in1(N__31117),
            .in2(_gnd_net_),
            .in3(N__29325),
            .lcout(),
            .ltout(N_508_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_2_LC_22_16_6.C_ON=1'b0;
    defparam M_this_data_count_q_2_LC_22_16_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_22_16_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 M_this_data_count_q_2_LC_22_16_6 (
            .in0(N__32254),
            .in1(N__29548),
            .in2(N__28657),
            .in3(N__32156),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31991),
            .ce(N__31676),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_3_LC_22_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_3_LC_22_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_3_LC_22_16_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_3_LC_22_16_7  (
            .in0(N__34358),
            .in1(N__31115),
            .in2(_gnd_net_),
            .in3(N__29539),
            .lcout(N_509),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_LC_22_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_LC_22_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a2_0_0_LC_22_17_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a2_0_0_LC_22_17_4  (
            .in0(N__33682),
            .in1(N__32789),
            .in2(N__34059),
            .in3(N__29180),
            .lcout(N_436),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNI60TF_15_LC_22_18_0.C_ON=1'b0;
    defparam M_this_data_count_q_RNI60TF_15_LC_22_18_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNI60TF_15_LC_22_18_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNI60TF_15_LC_22_18_0 (
            .in0(N__31404),
            .in1(N__32092),
            .in2(N__31372),
            .in3(N__31437),
            .lcout(M_this_state_d88_11),
            .ltout(M_this_state_d88_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNII1EE2_10_LC_22_18_1.C_ON=1'b0;
    defparam M_this_data_count_q_RNII1EE2_10_LC_22_18_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNII1EE2_10_LC_22_18_1.LUT_INIT=16'b1100000000000000;
    LogicCell40 M_this_data_count_q_RNII1EE2_10_LC_22_18_1 (
            .in0(_gnd_net_),
            .in1(N__31566),
            .in2(N__28645),
            .in3(N__28642),
            .lcout(M_this_state_d88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_0_0_LC_22_18_3.C_ON=1'b0;
    defparam M_this_state_q_RNO_0_0_LC_22_18_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_0_0_LC_22_18_3.LUT_INIT=16'b0100010001010101;
    LogicCell40 M_this_state_q_RNO_0_0_LC_22_18_3 (
            .in0(N__28633),
            .in1(N__31254),
            .in2(_gnd_net_),
            .in3(N__28504),
            .lcout(),
            .ltout(M_this_state_qsr_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_22_18_4.C_ON=1'b0;
    defparam M_this_state_q_0_LC_22_18_4.SEQ_MODE=4'b1001;
    defparam M_this_state_q_0_LC_22_18_4.LUT_INIT=16'b1111111111101111;
    LogicCell40 M_this_state_q_0_LC_22_18_4 (
            .in0(N__28624),
            .in1(N__28609),
            .in2(N__28597),
            .in3(N__28594),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32006),
            .ce(),
            .sr(N__32373));
    defparam \this_vga_signals.N_570_0_i_LC_22_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.N_570_0_i_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_570_0_i_LC_22_19_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \this_vga_signals.N_570_0_i_LC_22_19_3  (
            .in0(N__31253),
            .in1(N__28505),
            .in2(_gnd_net_),
            .in3(N__32434),
            .lcout(N_570_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_5_m_9_LC_22_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_5_m_9_LC_22_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_5_m_9_LC_22_19_5 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_5_m_9_LC_22_19_5  (
            .in0(N__30891),
            .in1(N__30684),
            .in2(N__33966),
            .in3(N__32834),
            .lcout(\this_vga_signals.M_this_external_address_d_5_mZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNIE44V9_0_LC_22_20_0.C_ON=1'b1;
    defparam M_this_external_address_q_RNIE44V9_0_LC_22_20_0.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNIE44V9_0_LC_22_20_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_external_address_q_RNIE44V9_0_LC_22_20_0 (
            .in0(_gnd_net_),
            .in1(N__28971),
            .in2(N__28786),
            .in3(N__28784),
            .lcout(M_this_external_address_q_RNIE44V9Z0Z_0),
            .ltout(),
            .carryin(bfn_22_20_0_),
            .carryout(un1_M_this_external_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_0_c_RNIGGGB_LC_22_20_1.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_0_c_RNIGGGB_LC_22_20_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_0_c_RNIGGGB_LC_22_20_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_0_c_RNIGGGB_LC_22_20_1 (
            .in0(_gnd_net_),
            .in1(N__30361),
            .in2(_gnd_net_),
            .in3(N__28765),
            .lcout(un1_M_this_external_address_q_cry_0_c_RNIGGGBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_0),
            .carryout(un1_M_this_external_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_1_c_RNIIJHB_LC_22_20_2.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_1_c_RNIIJHB_LC_22_20_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_1_c_RNIIJHB_LC_22_20_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_1_c_RNIIJHB_LC_22_20_2 (
            .in0(_gnd_net_),
            .in1(N__30292),
            .in2(_gnd_net_),
            .in3(N__28762),
            .lcout(un1_M_this_external_address_q_cry_1_c_RNIIJHBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_1),
            .carryout(un1_M_this_external_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_2_c_RNIKMIB_LC_22_20_3.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_2_c_RNIKMIB_LC_22_20_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_2_c_RNIKMIB_LC_22_20_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_2_c_RNIKMIB_LC_22_20_3 (
            .in0(_gnd_net_),
            .in1(N__29237),
            .in2(_gnd_net_),
            .in3(N__28759),
            .lcout(un1_M_this_external_address_q_cry_2_c_RNIKMIBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_2),
            .carryout(un1_M_this_external_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_3_c_RNIMPJB_LC_22_20_4.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_3_c_RNIMPJB_LC_22_20_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_3_c_RNIMPJB_LC_22_20_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_3_c_RNIMPJB_LC_22_20_4 (
            .in0(_gnd_net_),
            .in1(N__30227),
            .in2(_gnd_net_),
            .in3(N__28756),
            .lcout(un1_M_this_external_address_q_cry_3_c_RNIMPJBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_3),
            .carryout(un1_M_this_external_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_4_c_RNIOSKB_LC_22_20_5.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_4_c_RNIOSKB_LC_22_20_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_4_c_RNIOSKB_LC_22_20_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_external_address_q_cry_4_c_RNIOSKB_LC_22_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28748),
            .in3(N__28711),
            .lcout(un1_M_this_external_address_q_cry_4_c_RNIOSKBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_4),
            .carryout(un1_M_this_external_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_5_c_RNIQVLB_LC_22_20_6.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_5_c_RNIQVLB_LC_22_20_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_5_c_RNIQVLB_LC_22_20_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_5_c_RNIQVLB_LC_22_20_6 (
            .in0(_gnd_net_),
            .in1(N__28690),
            .in2(_gnd_net_),
            .in3(N__28663),
            .lcout(un1_M_this_external_address_q_cry_5_c_RNIQVLBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_5),
            .carryout(un1_M_this_external_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_6_c_RNIS2NB_LC_22_20_7.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_6_c_RNIS2NB_LC_22_20_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_6_c_RNIS2NB_LC_22_20_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_6_c_RNIS2NB_LC_22_20_7 (
            .in0(_gnd_net_),
            .in1(N__30965),
            .in2(_gnd_net_),
            .in3(N__28660),
            .lcout(un1_M_this_external_address_q_cry_6_c_RNIS2NBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_6),
            .carryout(un1_M_this_external_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_22_21_0.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_22_21_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_22_21_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_22_21_0 (
            .in0(_gnd_net_),
            .in1(N__29020),
            .in2(_gnd_net_),
            .in3(N__28909),
            .lcout(un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0),
            .ltout(),
            .carryin(bfn_22_21_0_),
            .carryout(un1_M_this_external_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_22_21_1.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_22_21_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_22_21_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_22_21_1 (
            .in0(_gnd_net_),
            .in1(N__30883),
            .in2(_gnd_net_),
            .in3(N__28906),
            .lcout(un1_M_this_external_address_q_cry_8_c_RNI09PBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_8),
            .carryout(un1_M_this_external_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_22_21_2.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_22_21_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_22_21_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_22_21_2 (
            .in0(_gnd_net_),
            .in1(N__30928),
            .in2(_gnd_net_),
            .in3(N__28903),
            .lcout(un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_9),
            .carryout(un1_M_this_external_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_22_21_3.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_22_21_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_22_21_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_22_21_3 (
            .in0(_gnd_net_),
            .in1(N__29295),
            .in2(_gnd_net_),
            .in3(N__28900),
            .lcout(un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_10),
            .carryout(un1_M_this_external_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_22_21_4.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_22_21_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_22_21_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_22_21_4 (
            .in0(_gnd_net_),
            .in1(N__30426),
            .in2(_gnd_net_),
            .in3(N__28897),
            .lcout(un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_11),
            .carryout(un1_M_this_external_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_22_21_5.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_22_21_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_22_21_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_22_21_5 (
            .in0(_gnd_net_),
            .in1(N__28884),
            .in2(_gnd_net_),
            .in3(N__28852),
            .lcout(un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_12),
            .carryout(un1_M_this_external_address_q_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_22_21_6.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_22_21_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_22_21_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_22_21_6 (
            .in0(_gnd_net_),
            .in1(N__28842),
            .in2(_gnd_net_),
            .in3(N__28792),
            .lcout(un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_13),
            .carryout(un1_M_this_external_address_q_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_22_21_7.C_ON=1'b0;
    defparam un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_22_21_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_22_21_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_22_21_7 (
            .in0(_gnd_net_),
            .in1(N__30195),
            .in2(_gnd_net_),
            .in3(N__28789),
            .lcout(un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_m_8_LC_22_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_8_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_8_LC_22_22_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_8_LC_22_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29028),
            .in3(N__30859),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_q_mZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_8_LC_22_22_1.C_ON=1'b0;
    defparam M_this_external_address_q_8_LC_22_22_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_8_LC_22_22_1.LUT_INIT=16'b1111111111110100;
    LogicCell40 M_this_external_address_q_8_LC_22_22_1 (
            .in0(N__30522),
            .in1(N__29047),
            .in2(N__29041),
            .in3(N__29002),
            .lcout(M_this_external_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32035),
            .ce(),
            .sr(N__32384));
    defparam \this_vga_signals.M_this_external_address_d_5_m_8_LC_22_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_5_m_8_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_5_m_8_LC_22_22_2 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_5_m_8_LC_22_22_2  (
            .in0(N__29021),
            .in1(N__33828),
            .in2(N__30698),
            .in3(N__32828),
            .lcout(\this_vga_signals.M_this_external_address_d_5_mZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_8_m_0_LC_22_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_8_m_0_LC_22_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_8_m_0_LC_22_22_3 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_8_m_0_LC_22_22_3  (
            .in0(N__32829),
            .in1(N__28967),
            .in2(N__33837),
            .in3(N__30860),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_d_8_mZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_0_LC_22_22_4.C_ON=1'b0;
    defparam M_this_external_address_q_0_LC_22_22_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_0_LC_22_22_4.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_external_address_q_0_LC_22_22_4 (
            .in0(N__28945),
            .in1(N__30521),
            .in2(N__28996),
            .in3(N__28993),
            .lcout(M_this_external_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32035),
            .ce(),
            .sr(N__32384));
    defparam \this_vga_signals.M_this_external_address_q_m_0_LC_22_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_0_LC_22_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_0_LC_22_22_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_0_LC_22_22_5  (
            .in0(N__30671),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28966),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_9_LC_22_22_7.C_ON=1'b0;
    defparam M_this_external_address_q_9_LC_22_22_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_9_LC_22_22_7.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_external_address_q_9_LC_22_22_7 (
            .in0(N__30523),
            .in1(N__30706),
            .in2(N__28939),
            .in3(N__28927),
            .lcout(M_this_external_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32035),
            .ce(),
            .sr(N__32384));
    defparam \this_vga_signals.M_this_external_address_d_5_m_11_LC_22_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_5_m_11_LC_22_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_5_m_11_LC_22_23_0 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_5_m_11_LC_22_23_0  (
            .in0(N__32853),
            .in1(N__29291),
            .in2(N__34331),
            .in3(N__30700),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_d_5_mZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_11_LC_22_23_1.C_ON=1'b0;
    defparam M_this_external_address_q_11_LC_22_23_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_11_LC_22_23_1.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_external_address_q_11_LC_22_23_1 (
            .in0(N__29269),
            .in1(N__30527),
            .in2(N__28921),
            .in3(N__28918),
            .lcout(M_this_external_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32040),
            .ce(),
            .sr(N__32387));
    defparam \this_vga_signals.M_this_external_address_q_m_11_LC_22_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_11_LC_22_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_11_LC_22_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_11_LC_22_23_2  (
            .in0(_gnd_net_),
            .in1(N__30848),
            .in2(_gnd_net_),
            .in3(N__29290),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_m_3_LC_22_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_3_LC_22_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_3_LC_22_23_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_3_LC_22_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29238),
            .in3(N__30699),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_q_mZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_3_LC_22_23_4.C_ON=1'b0;
    defparam M_this_external_address_q_3_LC_22_23_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_3_LC_22_23_4.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_external_address_q_3_LC_22_23_4 (
            .in0(N__30528),
            .in1(N__29209),
            .in2(N__29263),
            .in3(N__29260),
            .lcout(M_this_external_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32040),
            .ce(),
            .sr(N__32387));
    defparam \this_vga_signals.M_this_external_address_d_8_m_3_LC_22_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_8_m_3_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_8_m_3_LC_22_23_5 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_8_m_3_LC_22_23_5  (
            .in0(N__29230),
            .in1(N__34306),
            .in2(N__30861),
            .in3(N__32852),
            .lcout(\this_vga_signals.M_this_external_address_d_8_mZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_0_LC_22_24_0.C_ON=1'b0;
    defparam M_this_data_count_q_RNO_0_0_LC_22_24_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_0_LC_22_24_0.LUT_INIT=16'b1010010101011010;
    LogicCell40 M_this_data_count_q_RNO_0_0_LC_22_24_0 (
            .in0(N__29827),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29389),
            .lcout(M_this_data_count_q_s_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_7_0_a2_LC_23_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_7_0_a2_LC_23_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_7_0_a2_LC_23_15_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_7_0_a2_LC_23_15_0  (
            .in0(N__31231),
            .in1(N__29618),
            .in2(N__32932),
            .in3(N__29189),
            .lcout(),
            .ltout(\this_vga_signals.N_292_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_18_1_LC_23_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_18_1_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_18_1_LC_23_15_1 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_18_1_LC_23_15_1  (
            .in0(N__31128),
            .in1(N__31318),
            .in2(N__29089),
            .in3(N__29086),
            .lcout(\this_vga_signals.un1_M_this_state_q_18Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIAQQL_4_LC_23_15_2.C_ON=1'b0;
    defparam M_this_data_count_q_RNIAQQL_4_LC_23_15_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIAQQL_4_LC_23_15_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNIAQQL_4_LC_23_15_2 (
            .in0(N__29504),
            .in1(N__29447),
            .in2(N__31057),
            .in3(N__29477),
            .lcout(M_this_state_d88_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_0_LC_23_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_0_LC_23_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_0_LC_23_15_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_0_LC_23_15_4  (
            .in0(N__33813),
            .in1(N__31100),
            .in2(_gnd_net_),
            .in3(N__29382),
            .lcout(N_506),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_5_LC_23_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_5_LC_23_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_5_LC_23_15_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_5_LC_23_15_6  (
            .in0(N__33637),
            .in1(N__31101),
            .in2(_gnd_net_),
            .in3(N__29478),
            .lcout(N_511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_6_LC_23_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_6_LC_23_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_6_LC_23_15_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_6_LC_23_15_7  (
            .in0(N__29448),
            .in1(N__33496),
            .in2(_gnd_net_),
            .in3(N__31102),
            .lcout(N_512),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_3_LC_23_16_0.C_ON=1'b0;
    defparam M_this_data_count_q_3_LC_23_16_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_23_16_0.LUT_INIT=16'b0010001011110000;
    LogicCell40 M_this_data_count_q_3_LC_23_16_0 (
            .in0(N__29410),
            .in1(N__32238),
            .in2(N__29521),
            .in3(N__32157),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31998),
            .ce(N__31668),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_4_LC_23_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_4_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_4_LC_23_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_4_LC_23_16_1  (
            .in0(N__31107),
            .in1(N__33327),
            .in2(_gnd_net_),
            .in3(N__29508),
            .lcout(),
            .ltout(N_510_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_4_LC_23_16_2.C_ON=1'b0;
    defparam M_this_data_count_q_4_LC_23_16_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_23_16_2.LUT_INIT=16'b0011000010101010;
    LogicCell40 M_this_data_count_q_4_LC_23_16_2 (
            .in0(N__29488),
            .in1(N__32239),
            .in2(N__29404),
            .in3(N__32158),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31998),
            .ce(N__31668),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_5_LC_23_16_4.C_ON=1'b0;
    defparam M_this_data_count_q_5_LC_23_16_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_23_16_4.LUT_INIT=16'b0100010011110000;
    LogicCell40 M_this_data_count_q_5_LC_23_16_4 (
            .in0(N__32240),
            .in1(N__29401),
            .in2(N__29464),
            .in3(N__32159),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31998),
            .ce(N__31668),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_6_LC_23_16_6.C_ON=1'b0;
    defparam M_this_data_count_q_6_LC_23_16_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_23_16_6.LUT_INIT=16'b0100010011110000;
    LogicCell40 M_this_data_count_q_6_LC_23_16_6 (
            .in0(N__32241),
            .in1(N__29395),
            .in2(N__29434),
            .in3(N__32160),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31998),
            .ce(N__31668),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_c_0_LC_23_17_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_c_0_LC_23_17_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_c_0_LC_23_17_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 M_this_data_count_q_cry_c_0_LC_23_17_0 (
            .in0(_gnd_net_),
            .in1(N__29378),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_23_17_0_),
            .carryout(M_this_data_count_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_1_LC_23_17_1.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_1_LC_23_17_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_1_LC_23_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_1_LC_23_17_1 (
            .in0(_gnd_net_),
            .in1(N__29354),
            .in2(N__30071),
            .in3(N__29329),
            .lcout(M_this_data_count_q_s_1),
            .ltout(),
            .carryin(M_this_data_count_q_cry_0),
            .carryout(M_this_data_count_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_2_LC_23_17_2.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_2_LC_23_17_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_2_LC_23_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_2_LC_23_17_2 (
            .in0(_gnd_net_),
            .in1(N__29997),
            .in2(N__29326),
            .in3(N__29542),
            .lcout(M_this_data_count_q_s_2),
            .ltout(),
            .carryin(M_this_data_count_q_cry_1),
            .carryout(M_this_data_count_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_3_LC_23_17_3.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_3_LC_23_17_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_3_LC_23_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_3_LC_23_17_3 (
            .in0(_gnd_net_),
            .in1(N__29538),
            .in2(N__30072),
            .in3(N__29512),
            .lcout(M_this_data_count_q_s_3),
            .ltout(),
            .carryin(M_this_data_count_q_cry_2),
            .carryout(M_this_data_count_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_4_LC_23_17_4.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_4_LC_23_17_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_4_LC_23_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_4_LC_23_17_4 (
            .in0(_gnd_net_),
            .in1(N__30001),
            .in2(N__29509),
            .in3(N__29482),
            .lcout(M_this_data_count_q_s_4),
            .ltout(),
            .carryin(M_this_data_count_q_cry_3),
            .carryout(M_this_data_count_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_5_LC_23_17_5.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_5_LC_23_17_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_5_LC_23_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_5_LC_23_17_5 (
            .in0(_gnd_net_),
            .in1(N__29479),
            .in2(N__30073),
            .in3(N__29455),
            .lcout(M_this_data_count_q_s_5),
            .ltout(),
            .carryin(M_this_data_count_q_cry_4),
            .carryout(M_this_data_count_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_6_LC_23_17_6.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_6_LC_23_17_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_6_LC_23_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_6_LC_23_17_6 (
            .in0(_gnd_net_),
            .in1(N__30005),
            .in2(N__29452),
            .in3(N__29425),
            .lcout(M_this_data_count_q_s_6),
            .ltout(),
            .carryin(M_this_data_count_q_cry_5),
            .carryout(M_this_data_count_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_7_LC_23_17_7.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_7_LC_23_17_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_7_LC_23_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_7_LC_23_17_7 (
            .in0(_gnd_net_),
            .in1(N__31052),
            .in2(N__30074),
            .in3(N__29422),
            .lcout(M_this_data_count_q_s_7),
            .ltout(),
            .carryin(M_this_data_count_q_cry_6),
            .carryout(M_this_data_count_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_8_LC_23_18_0.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_8_LC_23_18_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_8_LC_23_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_8_LC_23_18_0 (
            .in0(_gnd_net_),
            .in1(N__30014),
            .in2(N__31591),
            .in3(N__29419),
            .lcout(M_this_data_count_q_s_8),
            .ltout(),
            .carryin(bfn_23_18_0_),
            .carryout(M_this_data_count_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_9_LC_23_18_1.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_9_LC_23_18_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_9_LC_23_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_9_LC_23_18_1 (
            .in0(_gnd_net_),
            .in1(N__31634),
            .in2(N__30076),
            .in3(N__29416),
            .lcout(M_this_data_count_q_s_9),
            .ltout(),
            .carryin(M_this_data_count_q_cry_8),
            .carryout(M_this_data_count_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_9_THRU_LUT4_0_LC_23_18_2.C_ON=1'b1;
    defparam M_this_data_count_q_cry_9_THRU_LUT4_0_LC_23_18_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_9_THRU_LUT4_0_LC_23_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_9_THRU_LUT4_0_LC_23_18_2 (
            .in0(_gnd_net_),
            .in1(N__30021),
            .in2(N__31546),
            .in3(N__29413),
            .lcout(M_this_data_count_q_cry_9_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_9),
            .carryout(M_this_data_count_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_11_LC_23_18_3.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_11_LC_23_18_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_11_LC_23_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_11_LC_23_18_3 (
            .in0(_gnd_net_),
            .in1(N__31610),
            .in2(N__30075),
            .in3(N__30169),
            .lcout(M_this_data_count_q_s_11),
            .ltout(),
            .carryin(M_this_data_count_q_cry_10),
            .carryout(M_this_data_count_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_12_LC_23_18_4.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_12_LC_23_18_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_12_LC_23_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_12_LC_23_18_4 (
            .in0(_gnd_net_),
            .in1(N__30012),
            .in2(N__31438),
            .in3(N__30166),
            .lcout(M_this_data_count_q_s_12),
            .ltout(),
            .carryin(M_this_data_count_q_cry_11),
            .carryout(M_this_data_count_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_12_THRU_LUT4_0_LC_23_18_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_12_THRU_LUT4_0_LC_23_18_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_12_THRU_LUT4_0_LC_23_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_12_THRU_LUT4_0_LC_23_18_5 (
            .in0(_gnd_net_),
            .in1(N__32086),
            .in2(N__30077),
            .in3(N__30163),
            .lcout(M_this_data_count_q_cry_12_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_12),
            .carryout(M_this_data_count_q_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_14_LC_23_18_6.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_14_LC_23_18_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_14_LC_23_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_14_LC_23_18_6 (
            .in0(_gnd_net_),
            .in1(N__30013),
            .in2(N__31405),
            .in3(N__29695),
            .lcout(M_this_data_count_q_s_14),
            .ltout(),
            .carryin(M_this_data_count_q_cry_13),
            .carryout(M_this_data_count_q_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_15_LC_23_18_7.C_ON=1'b0;
    defparam M_this_data_count_q_RNO_0_15_LC_23_18_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_15_LC_23_18_7.LUT_INIT=16'b1100110000110011;
    LogicCell40 M_this_data_count_q_RNO_0_15_LC_23_18_7 (
            .in0(_gnd_net_),
            .in1(N__31367),
            .in2(_gnd_net_),
            .in3(N__29692),
            .lcout(M_this_data_count_q_s_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_12_LC_23_19_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_12_LC_23_19_1 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_12_LC_23_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_sprites_ram.mem_radreg_12_LC_23_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29689),
            .lcout(\this_sprites_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32021),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_m_1_LC_23_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_1_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_1_LC_23_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_1_LC_23_19_5  (
            .in0(_gnd_net_),
            .in1(N__30362),
            .in2(_gnd_net_),
            .in3(N__30695),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_sn_m1_LC_23_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_sn_m1_LC_23_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_sn_m1_LC_23_19_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_sn_m1_LC_23_19_6  (
            .in0(N__32929),
            .in1(N__29619),
            .in2(_gnd_net_),
            .in3(N__32430),
            .lcout(M_this_data_count_q_3_sn_N_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_8_m_1_LC_23_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_8_m_1_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_8_m_1_LC_23_20_0 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_8_m_1_LC_23_20_0  (
            .in0(N__32843),
            .in1(N__30363),
            .in2(N__33992),
            .in3(N__30839),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_d_8_mZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_1_LC_23_20_1.C_ON=1'b0;
    defparam M_this_external_address_q_1_LC_23_20_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_1_LC_23_20_1.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_external_address_q_1_LC_23_20_1 (
            .in0(N__30391),
            .in1(N__30518),
            .in2(N__30385),
            .in3(N__30382),
            .lcout(M_this_external_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32026),
            .ce(),
            .sr(N__32374));
    defparam \this_vga_signals.M_this_external_address_d_8_m_2_LC_23_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_8_m_2_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_8_m_2_LC_23_20_3 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_8_m_2_LC_23_20_3  (
            .in0(N__30838),
            .in1(N__30299),
            .in2(N__34202),
            .in3(N__32844),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_d_8_mZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_2_LC_23_20_4.C_ON=1'b0;
    defparam M_this_external_address_q_2_LC_23_20_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_2_LC_23_20_4.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_external_address_q_2_LC_23_20_4 (
            .in0(N__30519),
            .in1(N__30340),
            .in2(N__30325),
            .in3(N__30322),
            .lcout(M_this_external_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32026),
            .ce(),
            .sr(N__32374));
    defparam M_this_external_address_q_4_LC_23_20_7.C_ON=1'b0;
    defparam M_this_external_address_q_4_LC_23_20_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_4_LC_23_20_7.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_external_address_q_4_LC_23_20_7 (
            .in0(N__30274),
            .in1(N__30520),
            .in2(N__30265),
            .in3(N__30253),
            .lcout(M_this_external_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32026),
            .ce(),
            .sr(N__32374));
    defparam \this_vga_signals.M_this_external_address_d_5_i_m_15_LC_23_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_5_i_m_15_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_5_i_m_15_LC_23_21_0 .LUT_INIT=16'b0000100000101010;
    LogicCell40 \this_vga_signals.M_this_external_address_d_5_i_m_15_LC_23_21_0  (
            .in0(N__30696),
            .in1(N__32846),
            .in2(N__33426),
            .in3(N__30194),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_d_5_i_mZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_15_LC_23_21_1.C_ON=1'b0;
    defparam M_this_external_address_q_15_LC_23_21_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_15_LC_23_21_1.LUT_INIT=16'b0000010100000100;
    LogicCell40 M_this_external_address_q_15_LC_23_21_1 (
            .in0(N__30175),
            .in1(N__30525),
            .in2(N__30214),
            .in3(N__30211),
            .lcout(M_this_external_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32036),
            .ce(),
            .sr(N__32379));
    defparam \this_vga_signals.M_this_external_address_q_i_m_15_LC_23_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_i_m_15_LC_23_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_i_m_15_LC_23_21_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_i_m_15_LC_23_21_2  (
            .in0(_gnd_net_),
            .in1(N__30193),
            .in2(_gnd_net_),
            .in3(N__30852),
            .lcout(\this_vga_signals.M_this_external_address_q_i_mZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_8_m_7_LC_23_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_8_m_7_LC_23_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_8_m_7_LC_23_21_3 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_8_m_7_LC_23_21_3  (
            .in0(N__32845),
            .in1(N__33421),
            .in2(N__30862),
            .in3(N__30971),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_d_8_mZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_7_LC_23_21_4.C_ON=1'b0;
    defparam M_this_external_address_q_7_LC_23_21_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_7_LC_23_21_4.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_external_address_q_7_LC_23_21_4 (
            .in0(N__30526),
            .in1(N__31015),
            .in2(N__31003),
            .in3(N__31000),
            .lcout(M_this_external_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32036),
            .ce(),
            .sr(N__32379));
    defparam \this_vga_signals.M_this_external_address_d_5_m_10_LC_23_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_5_m_10_LC_23_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_5_m_10_LC_23_21_6 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_5_m_10_LC_23_21_6  (
            .in0(N__30697),
            .in1(N__32847),
            .in2(N__34150),
            .in3(N__30932),
            .lcout(),
            .ltout(\this_vga_signals.M_this_external_address_d_5_mZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_10_LC_23_21_7.C_ON=1'b0;
    defparam M_this_external_address_q_10_LC_23_21_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_10_LC_23_21_7.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_external_address_q_10_LC_23_21_7 (
            .in0(N__30907),
            .in1(N__30524),
            .in2(N__30949),
            .in3(N__30946),
            .lcout(M_this_external_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32036),
            .ce(),
            .sr(N__32379));
    defparam \this_vga_signals.M_this_external_address_q_m_10_LC_23_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_10_LC_23_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_10_LC_23_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_10_LC_23_22_0  (
            .in0(_gnd_net_),
            .in1(N__30936),
            .in2(_gnd_net_),
            .in3(N__30856),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_m_12_LC_23_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_12_LC_23_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_12_LC_23_22_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_12_LC_23_22_1  (
            .in0(N__30857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30422),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_m_9_LC_23_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_m_9_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_m_9_LC_23_22_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_m_9_LC_23_22_2  (
            .in0(N__30887),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30858),
            .lcout(\this_vga_signals.M_this_external_address_q_mZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_5_m_12_LC_23_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_5_m_12_LC_23_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_5_m_12_LC_23_22_6 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_5_m_12_LC_23_22_6  (
            .in0(N__30421),
            .in1(N__30670),
            .in2(N__33326),
            .in3(N__32827),
            .lcout(\this_vga_signals.M_this_external_address_d_5_mZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_12_LC_23_23_3.C_ON=1'b0;
    defparam M_this_external_address_q_12_LC_23_23_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_12_LC_23_23_3.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_external_address_q_12_LC_23_23_3 (
            .in0(N__30535),
            .in1(N__30529),
            .in2(N__30454),
            .in3(N__30445),
            .lcout(M_this_external_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32044),
            .ce(),
            .sr(N__32385));
    defparam \this_vga_signals.M_this_map_ram_write_data_3_LC_23_29_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_3_LC_23_29_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_3_LC_23_29_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_3_LC_23_29_6  (
            .in0(N__34318),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33022),
            .lcout(M_this_map_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_e_0_LC_24_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_e_0_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_e_0_LC_24_15_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_e_0_LC_24_15_2  (
            .in0(N__32931),
            .in1(N__32723),
            .in2(_gnd_net_),
            .in3(N__32429),
            .lcout(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_7_0_LC_24_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_7_0_LC_24_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_7_0_LC_24_16_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o3_7_0_LC_24_16_1  (
            .in0(_gnd_net_),
            .in1(N__31317),
            .in2(_gnd_net_),
            .in3(N__31203),
            .lcout(N_391_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qe_0_i_LC_24_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qe_0_i_LC_24_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qe_0_i_LC_24_16_5 .LUT_INIT=16'b1111111100101010;
    LogicCell40 \this_vga_signals.M_this_data_count_qe_0_i_LC_24_16_5  (
            .in0(N__31210),
            .in1(N__31204),
            .in2(N__31148),
            .in3(N__32435),
            .lcout(M_this_data_count_qe_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_7_LC_24_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_7_LC_24_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_7_LC_24_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_7_LC_24_16_7  (
            .in0(N__33390),
            .in1(N__31053),
            .in2(_gnd_net_),
            .in3(N__31103),
            .lcout(N_513),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_7_LC_24_17_0.C_ON=1'b0;
    defparam M_this_data_count_q_7_LC_24_17_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_24_17_0.LUT_INIT=16'b0100010011110000;
    LogicCell40 M_this_data_count_q_7_LC_24_17_0 (
            .in0(N__32249),
            .in1(N__31072),
            .in2(N__31066),
            .in3(N__32165),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32012),
            .ce(N__31677),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_8_LC_24_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_8_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_8_LC_24_17_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_8_LC_24_17_1  (
            .in0(N__33835),
            .in1(N__31589),
            .in2(_gnd_net_),
            .in3(N__31515),
            .lcout(),
            .ltout(N_514_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_8_LC_24_17_2.C_ON=1'b0;
    defparam M_this_data_count_q_8_LC_24_17_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_24_17_2.LUT_INIT=16'b0101000011001100;
    LogicCell40 M_this_data_count_q_8_LC_24_17_2 (
            .in0(N__32250),
            .in1(N__31033),
            .in2(N__31027),
            .in3(N__32166),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32012),
            .ce(N__31677),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_9_LC_24_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_9_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_9_LC_24_17_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_9_LC_24_17_3  (
            .in0(N__34000),
            .in1(N__31635),
            .in2(_gnd_net_),
            .in3(N__31516),
            .lcout(),
            .ltout(N_515_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_9_LC_24_17_4.C_ON=1'b0;
    defparam M_this_data_count_q_9_LC_24_17_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_24_17_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 M_this_data_count_q_9_LC_24_17_4 (
            .in0(N__32251),
            .in1(N__31024),
            .in2(N__31018),
            .in3(N__32167),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32012),
            .ce(N__31677),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_11_LC_24_18_0.C_ON=1'b0;
    defparam M_this_data_count_q_11_LC_24_18_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_24_18_0.LUT_INIT=16'b0100010011110000;
    LogicCell40 M_this_data_count_q_11_LC_24_18_0 (
            .in0(N__32234),
            .in1(N__31348),
            .in2(N__31456),
            .in3(N__32161),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32022),
            .ce(N__31669),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_12_LC_24_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_12_LC_24_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_12_LC_24_18_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_12_LC_24_18_1  (
            .in0(N__33312),
            .in1(N__31436),
            .in2(_gnd_net_),
            .in3(N__31506),
            .lcout(),
            .ltout(N_518_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_12_LC_24_18_2.C_ON=1'b0;
    defparam M_this_data_count_q_12_LC_24_18_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_24_18_2.LUT_INIT=16'b0101000011001100;
    LogicCell40 M_this_data_count_q_12_LC_24_18_2 (
            .in0(N__32235),
            .in1(N__31447),
            .in2(N__31441),
            .in3(N__32162),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32022),
            .ce(N__31669),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_14_LC_24_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_14_LC_24_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_14_LC_24_18_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_14_LC_24_18_3  (
            .in0(N__33480),
            .in1(N__31403),
            .in2(_gnd_net_),
            .in3(N__31507),
            .lcout(),
            .ltout(N_520_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_14_LC_24_18_4.C_ON=1'b0;
    defparam M_this_data_count_q_14_LC_24_18_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_14_LC_24_18_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 M_this_data_count_q_14_LC_24_18_4 (
            .in0(N__32236),
            .in1(N__31414),
            .in2(N__31408),
            .in3(N__32163),
            .lcout(M_this_data_count_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32022),
            .ce(N__31669),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_15_LC_24_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_15_LC_24_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_15_LC_24_18_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_15_LC_24_18_5  (
            .in0(N__33406),
            .in1(N__31368),
            .in2(_gnd_net_),
            .in3(N__31508),
            .lcout(),
            .ltout(N_521_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_15_LC_24_18_6.C_ON=1'b0;
    defparam M_this_data_count_q_15_LC_24_18_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_15_LC_24_18_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 M_this_data_count_q_15_LC_24_18_6 (
            .in0(N__32237),
            .in1(N__31381),
            .in2(N__31375),
            .in3(N__32164),
            .lcout(M_this_data_count_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32022),
            .ce(N__31669),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_11_LC_24_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_11_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_11_LC_24_18_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_11_LC_24_18_7  (
            .in0(N__34357),
            .in1(N__31611),
            .in2(_gnd_net_),
            .in3(N__31505),
            .lcout(N_517),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_ns_10_LC_24_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_ns_10_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_ns_10_LC_24_19_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_ns_10_LC_24_19_0  (
            .in0(N__31342),
            .in1(N__32203),
            .in2(_gnd_net_),
            .in3(N__31480),
            .lcout(),
            .ltout(M_this_data_count_q_3_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_10_LC_24_19_1.C_ON=1'b0;
    defparam M_this_data_count_q_10_LC_24_19_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_24_19_1.LUT_INIT=16'b1111000010011001;
    LogicCell40 M_this_data_count_q_10_LC_24_19_1 (
            .in0(N__31544),
            .in1(N__32941),
            .in2(N__32935),
            .in3(N__32136),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32027),
            .ce(N__31678),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_e_8_LC_24_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_e_8_LC_24_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_e_8_LC_24_19_4 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_e_8_LC_24_19_4  (
            .in0(N__32930),
            .in1(N__32791),
            .in2(_gnd_net_),
            .in3(N__32428),
            .lcout(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8 ),
            .ltout(\this_vga_signals.M_this_data_count_q_3_0_eZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_am_13_LC_24_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_am_13_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_am_13_LC_24_19_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_am_13_LC_24_19_5  (
            .in0(N__33578),
            .in1(_gnd_net_),
            .in2(N__32269),
            .in3(N__32087),
            .lcout(),
            .ltout(\this_vga_signals.M_this_data_count_q_3_amZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_ns_13_LC_24_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_ns_13_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_ns_13_LC_24_19_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_ns_13_LC_24_19_6  (
            .in0(_gnd_net_),
            .in1(N__32266),
            .in2(N__32257),
            .in3(N__32204),
            .lcout(),
            .ltout(M_this_data_count_q_3_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_24_19_7.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_24_19_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_24_19_7.LUT_INIT=16'b1111000010011001;
    LogicCell40 M_this_data_count_q_13_LC_24_19_7 (
            .in0(N__32088),
            .in1(N__32176),
            .in2(N__32170),
            .in3(N__32137),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32027),
            .ce(N__31678),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNI8TRI_10_LC_24_20_1.C_ON=1'b0;
    defparam M_this_data_count_q_RNI8TRI_10_LC_24_20_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNI8TRI_10_LC_24_20_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNI8TRI_10_LC_24_20_1 (
            .in0(N__31537),
            .in1(N__31636),
            .in2(N__31615),
            .in3(N__31590),
            .lcout(M_this_state_d88_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_am_10_LC_24_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_am_10_LC_24_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_am_10_LC_24_21_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_am_10_LC_24_21_1  (
            .in0(N__34129),
            .in1(N__31545),
            .in2(_gnd_net_),
            .in3(N__31514),
            .lcout(\this_vga_signals.M_this_data_count_q_3_amZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_6_LC_24_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_6_LC_24_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_6_LC_24_24_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_6_LC_24_24_1  (
            .in0(N__33508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33005),
            .lcout(M_this_map_ram_write_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_7_LC_24_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_7_LC_24_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_7_LC_24_24_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_7_LC_24_24_2  (
            .in0(N__33006),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33422),
            .lcout(M_this_map_ram_write_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI5S7_7_LC_24_26_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI5S7_7_LC_24_26_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI5S7_7_LC_24_26_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_haddress_q_RNI5S7_7_LC_24_26_3  (
            .in0(_gnd_net_),
            .in1(N__33175),
            .in2(_gnd_net_),
            .in3(N__33125),
            .lcout(M_this_ppu_map_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIIT3_6_LC_24_26_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIIT3_6_LC_24_26_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIIT3_6_LC_24_26_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_ppu.M_haddress_q_RNIIT3_6_LC_24_26_4  (
            .in0(N__33126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_ppu_vram_addr_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_2_LC_24_28_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_2_LC_24_28_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_2_LC_24_28_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_2_LC_24_28_5  (
            .in0(N__33024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34144),
            .lcout(M_this_map_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_1_LC_24_28_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_1_LC_24_28_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_1_LC_24_28_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_1_LC_24_28_6  (
            .in0(N__33945),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33023),
            .lcout(M_this_map_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_LC_24_29_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_LC_24_29_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_LC_24_29_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_LC_24_29_2  (
            .in0(N__33043),
            .in1(N__33814),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_map_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_5_LC_24_31_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_5_LC_24_31_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_5_LC_24_31_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_5_LC_24_31_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33046),
            .in3(N__33613),
            .lcout(M_this_map_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_4_LC_24_31_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_4_LC_24_31_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_4_LC_24_31_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_4_LC_24_31_5  (
            .in0(_gnd_net_),
            .in1(N__33039),
            .in2(_gnd_net_),
            .in3(N__33266),
            .lcout(M_this_map_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d21_2_LC_26_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d21_2_LC_26_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d21_2_LC_26_19_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_external_address_d21_2_LC_26_19_0  (
            .in0(N__34343),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34151),
            .lcout(\this_vga_signals.M_this_external_address_d21Z0Z_2 ),
            .ltout(\this_vga_signals.M_this_external_address_d21Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d21_LC_26_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d21_LC_26_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d21_LC_26_19_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_vga_signals.M_this_external_address_d21_LC_26_19_1  (
            .in0(N__33198),
            .in1(N__33970),
            .in2(N__34066),
            .in3(N__33822),
            .lcout(\this_vga_signals.M_this_external_address_dZ0Z21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d22_LC_26_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d22_LC_26_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d22_LC_26_19_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_d22_LC_26_19_5  (
            .in0(N__33199),
            .in1(N__33971),
            .in2(N__33850),
            .in3(N__33823),
            .lcout(\this_vga_signals.M_this_external_address_dZ0Z22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d21_6_LC_26_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d21_6_LC_26_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d21_6_LC_26_21_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_external_address_d21_6_LC_26_21_2  (
            .in0(N__33595),
            .in1(N__33519),
            .in2(N__33389),
            .in3(N__33248),
            .lcout(\this_vga_signals.M_this_external_address_d21Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
