// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 9 2022 09:54:28

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    rgb,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    debug,
    clk);

    input [15:0] port_address;
    input [7:0] port_data;
    output [5:0] rgb;
    output vsync;
    output vblank;
    input rst_n;
    input port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    output debug;
    input clk;

    wire N__20798;
    wire N__20797;
    wire N__20796;
    wire N__20787;
    wire N__20786;
    wire N__20785;
    wire N__20778;
    wire N__20777;
    wire N__20776;
    wire N__20769;
    wire N__20768;
    wire N__20767;
    wire N__20760;
    wire N__20759;
    wire N__20758;
    wire N__20751;
    wire N__20750;
    wire N__20749;
    wire N__20742;
    wire N__20741;
    wire N__20740;
    wire N__20733;
    wire N__20732;
    wire N__20731;
    wire N__20724;
    wire N__20723;
    wire N__20722;
    wire N__20715;
    wire N__20714;
    wire N__20713;
    wire N__20706;
    wire N__20705;
    wire N__20704;
    wire N__20697;
    wire N__20696;
    wire N__20695;
    wire N__20688;
    wire N__20687;
    wire N__20686;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20670;
    wire N__20669;
    wire N__20668;
    wire N__20661;
    wire N__20660;
    wire N__20659;
    wire N__20652;
    wire N__20651;
    wire N__20650;
    wire N__20643;
    wire N__20642;
    wire N__20641;
    wire N__20634;
    wire N__20633;
    wire N__20632;
    wire N__20625;
    wire N__20624;
    wire N__20623;
    wire N__20616;
    wire N__20615;
    wire N__20614;
    wire N__20607;
    wire N__20606;
    wire N__20605;
    wire N__20598;
    wire N__20597;
    wire N__20596;
    wire N__20589;
    wire N__20588;
    wire N__20587;
    wire N__20580;
    wire N__20579;
    wire N__20578;
    wire N__20571;
    wire N__20570;
    wire N__20569;
    wire N__20562;
    wire N__20561;
    wire N__20560;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20544;
    wire N__20543;
    wire N__20542;
    wire N__20535;
    wire N__20534;
    wire N__20533;
    wire N__20526;
    wire N__20525;
    wire N__20524;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20508;
    wire N__20507;
    wire N__20506;
    wire N__20499;
    wire N__20498;
    wire N__20497;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20338;
    wire N__20335;
    wire N__20334;
    wire N__20333;
    wire N__20332;
    wire N__20331;
    wire N__20330;
    wire N__20329;
    wire N__20326;
    wire N__20325;
    wire N__20324;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20310;
    wire N__20309;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20291;
    wire N__20290;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20266;
    wire N__20263;
    wire N__20262;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20232;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20201;
    wire N__20198;
    wire N__20191;
    wire N__20182;
    wire N__20177;
    wire N__20168;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20150;
    wire N__20149;
    wire N__20148;
    wire N__20145;
    wire N__20140;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19879;
    wire N__19878;
    wire N__19877;
    wire N__19876;
    wire N__19873;
    wire N__19872;
    wire N__19871;
    wire N__19870;
    wire N__19869;
    wire N__19868;
    wire N__19863;
    wire N__19854;
    wire N__19851;
    wire N__19844;
    wire N__19843;
    wire N__19842;
    wire N__19841;
    wire N__19834;
    wire N__19831;
    wire N__19824;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19814;
    wire N__19809;
    wire N__19806;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19772;
    wire N__19771;
    wire N__19768;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19727;
    wire N__19724;
    wire N__19723;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19715;
    wire N__19712;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19694;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19678;
    wire N__19675;
    wire N__19670;
    wire N__19667;
    wire N__19662;
    wire N__19661;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19643;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19597;
    wire N__19596;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19582;
    wire N__19581;
    wire N__19580;
    wire N__19579;
    wire N__19576;
    wire N__19571;
    wire N__19568;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19545;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19502;
    wire N__19501;
    wire N__19500;
    wire N__19499;
    wire N__19498;
    wire N__19497;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19480;
    wire N__19477;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19462;
    wire N__19459;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19443;
    wire N__19440;
    wire N__19433;
    wire N__19432;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19410;
    wire N__19403;
    wire N__19402;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19394;
    wire N__19393;
    wire N__19392;
    wire N__19391;
    wire N__19390;
    wire N__19387;
    wire N__19386;
    wire N__19383;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19341;
    wire N__19336;
    wire N__19333;
    wire N__19328;
    wire N__19325;
    wire N__19316;
    wire N__19315;
    wire N__19314;
    wire N__19313;
    wire N__19312;
    wire N__19311;
    wire N__19310;
    wire N__19309;
    wire N__19306;
    wire N__19301;
    wire N__19298;
    wire N__19297;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19278;
    wire N__19277;
    wire N__19276;
    wire N__19273;
    wire N__19266;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19251;
    wire N__19248;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19226;
    wire N__19223;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18943;
    wire N__18940;
    wire N__18937;
    wire N__18936;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18877;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18866;
    wire N__18865;
    wire N__18864;
    wire N__18863;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18851;
    wire N__18844;
    wire N__18837;
    wire N__18834;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18820;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18437;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18397;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18382;
    wire N__18379;
    wire N__18374;
    wire N__18371;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18363;
    wire N__18360;
    wire N__18359;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18342;
    wire N__18341;
    wire N__18340;
    wire N__18339;
    wire N__18338;
    wire N__18337;
    wire N__18336;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18322;
    wire N__18319;
    wire N__18316;
    wire N__18309;
    wire N__18304;
    wire N__18303;
    wire N__18298;
    wire N__18297;
    wire N__18296;
    wire N__18291;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18260;
    wire N__18239;
    wire N__18238;
    wire N__18237;
    wire N__18236;
    wire N__18235;
    wire N__18234;
    wire N__18233;
    wire N__18232;
    wire N__18231;
    wire N__18230;
    wire N__18229;
    wire N__18228;
    wire N__18227;
    wire N__18226;
    wire N__18225;
    wire N__18224;
    wire N__18223;
    wire N__18222;
    wire N__18221;
    wire N__18220;
    wire N__18219;
    wire N__18218;
    wire N__18217;
    wire N__18216;
    wire N__18215;
    wire N__18214;
    wire N__18213;
    wire N__18212;
    wire N__18211;
    wire N__18210;
    wire N__18209;
    wire N__18208;
    wire N__18207;
    wire N__18206;
    wire N__18205;
    wire N__18204;
    wire N__18203;
    wire N__18202;
    wire N__18201;
    wire N__18200;
    wire N__18199;
    wire N__18198;
    wire N__18197;
    wire N__18196;
    wire N__18195;
    wire N__18194;
    wire N__18193;
    wire N__18192;
    wire N__18191;
    wire N__18190;
    wire N__18189;
    wire N__18188;
    wire N__18187;
    wire N__18186;
    wire N__18185;
    wire N__18184;
    wire N__18183;
    wire N__18182;
    wire N__18181;
    wire N__18180;
    wire N__18179;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18049;
    wire N__18046;
    wire N__18045;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18008;
    wire N__18005;
    wire N__18004;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17996;
    wire N__17993;
    wire N__17992;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17964;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17943;
    wire N__17938;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17878;
    wire N__17875;
    wire N__17874;
    wire N__17873;
    wire N__17870;
    wire N__17869;
    wire N__17866;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17854;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17833;
    wire N__17832;
    wire N__17831;
    wire N__17828;
    wire N__17823;
    wire N__17816;
    wire N__17809;
    wire N__17806;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17779;
    wire N__17776;
    wire N__17775;
    wire N__17774;
    wire N__17771;
    wire N__17770;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17754;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17627;
    wire N__17624;
    wire N__17623;
    wire N__17622;
    wire N__17619;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17590;
    wire N__17587;
    wire N__17582;
    wire N__17581;
    wire N__17578;
    wire N__17577;
    wire N__17574;
    wire N__17573;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17556;
    wire N__17555;
    wire N__17550;
    wire N__17547;
    wire N__17544;
    wire N__17541;
    wire N__17538;
    wire N__17535;
    wire N__17530;
    wire N__17525;
    wire N__17520;
    wire N__17519;
    wire N__17516;
    wire N__17511;
    wire N__17508;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17350;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17339;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17323;
    wire N__17322;
    wire N__17321;
    wire N__17320;
    wire N__17319;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17311;
    wire N__17310;
    wire N__17305;
    wire N__17302;
    wire N__17301;
    wire N__17300;
    wire N__17299;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17243;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17200;
    wire N__17199;
    wire N__17198;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17187;
    wire N__17182;
    wire N__17181;
    wire N__17180;
    wire N__17179;
    wire N__17178;
    wire N__17171;
    wire N__17170;
    wire N__17169;
    wire N__17168;
    wire N__17165;
    wire N__17164;
    wire N__17163;
    wire N__17162;
    wire N__17161;
    wire N__17160;
    wire N__17159;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17145;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17119;
    wire N__17118;
    wire N__17117;
    wire N__17116;
    wire N__17115;
    wire N__17112;
    wire N__17111;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17103;
    wire N__17102;
    wire N__17101;
    wire N__17094;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17074;
    wire N__17071;
    wire N__17064;
    wire N__17059;
    wire N__17050;
    wire N__17045;
    wire N__17042;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17002;
    wire N__17001;
    wire N__17000;
    wire N__16999;
    wire N__16994;
    wire N__16987;
    wire N__16986;
    wire N__16985;
    wire N__16984;
    wire N__16979;
    wire N__16972;
    wire N__16971;
    wire N__16970;
    wire N__16969;
    wire N__16968;
    wire N__16967;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16934;
    wire N__16933;
    wire N__16932;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16924;
    wire N__16921;
    wire N__16916;
    wire N__16909;
    wire N__16908;
    wire N__16907;
    wire N__16906;
    wire N__16905;
    wire N__16904;
    wire N__16903;
    wire N__16898;
    wire N__16891;
    wire N__16888;
    wire N__16887;
    wire N__16884;
    wire N__16881;
    wire N__16880;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16864;
    wire N__16861;
    wire N__16858;
    wire N__16847;
    wire N__16846;
    wire N__16845;
    wire N__16844;
    wire N__16843;
    wire N__16842;
    wire N__16837;
    wire N__16830;
    wire N__16827;
    wire N__16826;
    wire N__16825;
    wire N__16824;
    wire N__16823;
    wire N__16818;
    wire N__16811;
    wire N__16810;
    wire N__16809;
    wire N__16808;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16786;
    wire N__16783;
    wire N__16780;
    wire N__16769;
    wire N__16768;
    wire N__16767;
    wire N__16766;
    wire N__16763;
    wire N__16762;
    wire N__16761;
    wire N__16760;
    wire N__16755;
    wire N__16748;
    wire N__16747;
    wire N__16744;
    wire N__16741;
    wire N__16740;
    wire N__16735;
    wire N__16728;
    wire N__16727;
    wire N__16724;
    wire N__16723;
    wire N__16722;
    wire N__16721;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16688;
    wire N__16687;
    wire N__16682;
    wire N__16679;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16636;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16574;
    wire N__16571;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16557;
    wire N__16556;
    wire N__16551;
    wire N__16548;
    wire N__16547;
    wire N__16546;
    wire N__16543;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16508;
    wire N__16507;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16483;
    wire N__16478;
    wire N__16477;
    wire N__16474;
    wire N__16473;
    wire N__16472;
    wire N__16471;
    wire N__16466;
    wire N__16463;
    wire N__16462;
    wire N__16461;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16453;
    wire N__16452;
    wire N__16451;
    wire N__16450;
    wire N__16449;
    wire N__16444;
    wire N__16439;
    wire N__16438;
    wire N__16437;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16422;
    wire N__16419;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16401;
    wire N__16396;
    wire N__16391;
    wire N__16376;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16328;
    wire N__16327;
    wire N__16326;
    wire N__16325;
    wire N__16322;
    wire N__16321;
    wire N__16320;
    wire N__16319;
    wire N__16318;
    wire N__16317;
    wire N__16316;
    wire N__16315;
    wire N__16314;
    wire N__16313;
    wire N__16312;
    wire N__16311;
    wire N__16310;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16302;
    wire N__16301;
    wire N__16300;
    wire N__16299;
    wire N__16298;
    wire N__16297;
    wire N__16296;
    wire N__16295;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16287;
    wire N__16286;
    wire N__16285;
    wire N__16284;
    wire N__16281;
    wire N__16270;
    wire N__16267;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16247;
    wire N__16242;
    wire N__16241;
    wire N__16240;
    wire N__16235;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16215;
    wire N__16208;
    wire N__16199;
    wire N__16196;
    wire N__16193;
    wire N__16188;
    wire N__16183;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16147;
    wire N__16146;
    wire N__16143;
    wire N__16142;
    wire N__16141;
    wire N__16140;
    wire N__16137;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16125;
    wire N__16122;
    wire N__16121;
    wire N__16114;
    wire N__16107;
    wire N__16104;
    wire N__16101;
    wire N__16094;
    wire N__16093;
    wire N__16090;
    wire N__16089;
    wire N__16088;
    wire N__16087;
    wire N__16086;
    wire N__16085;
    wire N__16084;
    wire N__16083;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16069;
    wire N__16062;
    wire N__16061;
    wire N__16060;
    wire N__16059;
    wire N__16058;
    wire N__16057;
    wire N__16056;
    wire N__16051;
    wire N__16042;
    wire N__16033;
    wire N__16028;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15905;
    wire N__15904;
    wire N__15903;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15882;
    wire N__15881;
    wire N__15880;
    wire N__15879;
    wire N__15876;
    wire N__15871;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15855;
    wire N__15852;
    wire N__15845;
    wire N__15842;
    wire N__15841;
    wire N__15840;
    wire N__15839;
    wire N__15838;
    wire N__15837;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15825;
    wire N__15820;
    wire N__15817;
    wire N__15816;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15783;
    wire N__15778;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15731;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15597;
    wire N__15594;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15577;
    wire N__15576;
    wire N__15575;
    wire N__15574;
    wire N__15573;
    wire N__15570;
    wire N__15569;
    wire N__15566;
    wire N__15565;
    wire N__15564;
    wire N__15563;
    wire N__15562;
    wire N__15559;
    wire N__15558;
    wire N__15557;
    wire N__15556;
    wire N__15555;
    wire N__15548;
    wire N__15541;
    wire N__15538;
    wire N__15531;
    wire N__15530;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15522;
    wire N__15517;
    wire N__15514;
    wire N__15511;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15493;
    wire N__15490;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15326;
    wire N__15325;
    wire N__15324;
    wire N__15323;
    wire N__15322;
    wire N__15321;
    wire N__15316;
    wire N__15313;
    wire N__15312;
    wire N__15309;
    wire N__15308;
    wire N__15307;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15274;
    wire N__15271;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15257;
    wire N__15256;
    wire N__15249;
    wire N__15244;
    wire N__15241;
    wire N__15236;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15127;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14962;
    wire N__14959;
    wire N__14956;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14948;
    wire N__14947;
    wire N__14944;
    wire N__14939;
    wire N__14938;
    wire N__14937;
    wire N__14936;
    wire N__14931;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14906;
    wire N__14905;
    wire N__14904;
    wire N__14901;
    wire N__14898;
    wire N__14895;
    wire N__14892;
    wire N__14891;
    wire N__14890;
    wire N__14889;
    wire N__14884;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14716;
    wire N__14713;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14698;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14568;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14556;
    wire N__14549;
    wire N__14546;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14491;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14479;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14440;
    wire N__14437;
    wire N__14436;
    wire N__14435;
    wire N__14434;
    wire N__14431;
    wire N__14430;
    wire N__14427;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14419;
    wire N__14418;
    wire N__14415;
    wire N__14414;
    wire N__14413;
    wire N__14412;
    wire N__14409;
    wire N__14406;
    wire N__14403;
    wire N__14400;
    wire N__14399;
    wire N__14398;
    wire N__14393;
    wire N__14390;
    wire N__14389;
    wire N__14388;
    wire N__14387;
    wire N__14386;
    wire N__14385;
    wire N__14382;
    wire N__14379;
    wire N__14376;
    wire N__14373;
    wire N__14370;
    wire N__14369;
    wire N__14368;
    wire N__14363;
    wire N__14358;
    wire N__14355;
    wire N__14352;
    wire N__14351;
    wire N__14346;
    wire N__14343;
    wire N__14340;
    wire N__14339;
    wire N__14338;
    wire N__14337;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14327;
    wire N__14320;
    wire N__14315;
    wire N__14312;
    wire N__14311;
    wire N__14308;
    wire N__14307;
    wire N__14306;
    wire N__14305;
    wire N__14298;
    wire N__14295;
    wire N__14292;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14271;
    wire N__14266;
    wire N__14263;
    wire N__14256;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14234;
    wire N__14227;
    wire N__14224;
    wire N__14223;
    wire N__14220;
    wire N__14217;
    wire N__14214;
    wire N__14209;
    wire N__14204;
    wire N__14199;
    wire N__14194;
    wire N__14187;
    wire N__14184;
    wire N__14183;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14172;
    wire N__14169;
    wire N__14164;
    wire N__14157;
    wire N__14154;
    wire N__14151;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14131;
    wire N__14128;
    wire N__14123;
    wire N__14120;
    wire N__14113;
    wire N__14110;
    wire N__14105;
    wire N__14096;
    wire N__14093;
    wire N__14092;
    wire N__14091;
    wire N__14090;
    wire N__14085;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14057;
    wire N__14054;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13870;
    wire N__13867;
    wire N__13866;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13828;
    wire N__13825;
    wire N__13822;
    wire N__13819;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13802;
    wire N__13799;
    wire N__13796;
    wire N__13793;
    wire N__13792;
    wire N__13789;
    wire N__13788;
    wire N__13787;
    wire N__13784;
    wire N__13779;
    wire N__13776;
    wire N__13775;
    wire N__13774;
    wire N__13771;
    wire N__13770;
    wire N__13769;
    wire N__13766;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13751;
    wire N__13750;
    wire N__13747;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13731;
    wire N__13726;
    wire N__13721;
    wire N__13714;
    wire N__13711;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13697;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13681;
    wire N__13678;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13543;
    wire N__13542;
    wire N__13539;
    wire N__13536;
    wire N__13533;
    wire N__13530;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13408;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13398;
    wire N__13395;
    wire N__13392;
    wire N__13387;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13270;
    wire N__13269;
    wire N__13266;
    wire N__13263;
    wire N__13260;
    wire N__13257;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13135;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13099;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13087;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13067;
    wire N__13066;
    wire N__13063;
    wire N__13060;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13039;
    wire N__13038;
    wire N__13033;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13010;
    wire N__13009;
    wire N__13008;
    wire N__13007;
    wire N__13006;
    wire N__13003;
    wire N__12998;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12988;
    wire N__12987;
    wire N__12986;
    wire N__12981;
    wire N__12976;
    wire N__12973;
    wire N__12968;
    wire N__12963;
    wire N__12960;
    wire N__12959;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12931;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12890;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12856;
    wire N__12855;
    wire N__12852;
    wire N__12847;
    wire N__12842;
    wire N__12841;
    wire N__12838;
    wire N__12835;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12823;
    wire N__12822;
    wire N__12821;
    wire N__12818;
    wire N__12811;
    wire N__12808;
    wire N__12805;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12781;
    wire N__12778;
    wire N__12775;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12745;
    wire N__12744;
    wire N__12741;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12628;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12608;
    wire N__12607;
    wire N__12604;
    wire N__12601;
    wire N__12598;
    wire N__12593;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12552;
    wire N__12549;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12527;
    wire N__12524;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12509;
    wire N__12508;
    wire N__12505;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12475;
    wire N__12474;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12460;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12441;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12429;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12415;
    wire N__12410;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12394;
    wire N__12391;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12364;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12356;
    wire N__12355;
    wire N__12354;
    wire N__12353;
    wire N__12352;
    wire N__12351;
    wire N__12350;
    wire N__12349;
    wire N__12348;
    wire N__12347;
    wire N__12344;
    wire N__12337;
    wire N__12336;
    wire N__12335;
    wire N__12334;
    wire N__12333;
    wire N__12332;
    wire N__12331;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12316;
    wire N__12313;
    wire N__12306;
    wire N__12305;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12286;
    wire N__12281;
    wire N__12278;
    wire N__12273;
    wire N__12264;
    wire N__12259;
    wire N__12258;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12247;
    wire N__12242;
    wire N__12237;
    wire N__12234;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12204;
    wire N__12199;
    wire N__12182;
    wire N__12181;
    wire N__12180;
    wire N__12179;
    wire N__12178;
    wire N__12175;
    wire N__12174;
    wire N__12173;
    wire N__12172;
    wire N__12171;
    wire N__12170;
    wire N__12169;
    wire N__12168;
    wire N__12165;
    wire N__12162;
    wire N__12157;
    wire N__12152;
    wire N__12149;
    wire N__12144;
    wire N__12141;
    wire N__12140;
    wire N__12139;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12127;
    wire N__12124;
    wire N__12117;
    wire N__12114;
    wire N__12109;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12095;
    wire N__12092;
    wire N__12087;
    wire N__12084;
    wire N__12081;
    wire N__12076;
    wire N__12073;
    wire N__12070;
    wire N__12059;
    wire N__12058;
    wire N__12057;
    wire N__12056;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12046;
    wire N__12041;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11902;
    wire N__11901;
    wire N__11898;
    wire N__11897;
    wire N__11896;
    wire N__11893;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11873;
    wire N__11872;
    wire N__11871;
    wire N__11870;
    wire N__11867;
    wire N__11864;
    wire N__11859;
    wire N__11852;
    wire N__11849;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11746;
    wire N__11745;
    wire N__11742;
    wire N__11737;
    wire N__11736;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11715;
    wire N__11708;
    wire N__11707;
    wire N__11706;
    wire N__11705;
    wire N__11704;
    wire N__11703;
    wire N__11702;
    wire N__11701;
    wire N__11700;
    wire N__11699;
    wire N__11694;
    wire N__11693;
    wire N__11690;
    wire N__11689;
    wire N__11688;
    wire N__11687;
    wire N__11686;
    wire N__11677;
    wire N__11670;
    wire N__11667;
    wire N__11664;
    wire N__11661;
    wire N__11660;
    wire N__11655;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11618;
    wire N__11615;
    wire N__11614;
    wire N__11611;
    wire N__11610;
    wire N__11607;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11582;
    wire N__11579;
    wire N__11578;
    wire N__11577;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11567;
    wire N__11562;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11505;
    wire N__11504;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11496;
    wire N__11493;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11474;
    wire N__11465;
    wire N__11464;
    wire N__11463;
    wire N__11462;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11458;
    wire N__11457;
    wire N__11456;
    wire N__11455;
    wire N__11452;
    wire N__11451;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11443;
    wire N__11442;
    wire N__11439;
    wire N__11438;
    wire N__11437;
    wire N__11436;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11428;
    wire N__11427;
    wire N__11426;
    wire N__11423;
    wire N__11422;
    wire N__11419;
    wire N__11418;
    wire N__11417;
    wire N__11414;
    wire N__11413;
    wire N__11410;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11406;
    wire N__11403;
    wire N__11396;
    wire N__11395;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11368;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11349;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11337;
    wire N__11332;
    wire N__11331;
    wire N__11328;
    wire N__11323;
    wire N__11318;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11298;
    wire N__11295;
    wire N__11290;
    wire N__11289;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11271;
    wire N__11270;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11254;
    wire N__11245;
    wire N__11242;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11219;
    wire N__11216;
    wire N__11209;
    wire N__11198;
    wire N__11195;
    wire N__11194;
    wire N__11193;
    wire N__11192;
    wire N__11191;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11183;
    wire N__11180;
    wire N__11175;
    wire N__11174;
    wire N__11173;
    wire N__11170;
    wire N__11169;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11155;
    wire N__11150;
    wire N__11149;
    wire N__11148;
    wire N__11147;
    wire N__11146;
    wire N__11145;
    wire N__11144;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11126;
    wire N__11119;
    wire N__11114;
    wire N__11109;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11077;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11044;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11006;
    wire N__11005;
    wire N__11002;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10988;
    wire N__10987;
    wire N__10982;
    wire N__10981;
    wire N__10980;
    wire N__10977;
    wire N__10972;
    wire N__10971;
    wire N__10970;
    wire N__10969;
    wire N__10968;
    wire N__10967;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10950;
    wire N__10949;
    wire N__10944;
    wire N__10937;
    wire N__10934;
    wire N__10925;
    wire N__10916;
    wire N__10915;
    wire N__10914;
    wire N__10913;
    wire N__10912;
    wire N__10907;
    wire N__10906;
    wire N__10903;
    wire N__10902;
    wire N__10901;
    wire N__10900;
    wire N__10899;
    wire N__10894;
    wire N__10891;
    wire N__10884;
    wire N__10883;
    wire N__10882;
    wire N__10881;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10853;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10774;
    wire N__10773;
    wire N__10772;
    wire N__10771;
    wire N__10770;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10758;
    wire N__10751;
    wire N__10742;
    wire N__10741;
    wire N__10740;
    wire N__10739;
    wire N__10738;
    wire N__10737;
    wire N__10734;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10722;
    wire N__10715;
    wire N__10706;
    wire N__10705;
    wire N__10704;
    wire N__10703;
    wire N__10702;
    wire N__10701;
    wire N__10696;
    wire N__10693;
    wire N__10690;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10673;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10654;
    wire N__10653;
    wire N__10650;
    wire N__10645;
    wire N__10640;
    wire N__10639;
    wire N__10638;
    wire N__10637;
    wire N__10636;
    wire N__10633;
    wire N__10632;
    wire N__10631;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10616;
    wire N__10609;
    wire N__10598;
    wire N__10595;
    wire N__10594;
    wire N__10593;
    wire N__10592;
    wire N__10591;
    wire N__10590;
    wire N__10589;
    wire N__10588;
    wire N__10587;
    wire N__10584;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10564;
    wire N__10553;
    wire N__10552;
    wire N__10551;
    wire N__10550;
    wire N__10549;
    wire N__10548;
    wire N__10545;
    wire N__10536;
    wire N__10535;
    wire N__10534;
    wire N__10531;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10511;
    wire N__10510;
    wire N__10509;
    wire N__10508;
    wire N__10507;
    wire N__10506;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10494;
    wire N__10487;
    wire N__10478;
    wire N__10475;
    wire N__10474;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10420;
    wire N__10417;
    wire N__10414;
    wire N__10413;
    wire N__10412;
    wire N__10411;
    wire N__10410;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10392;
    wire N__10387;
    wire N__10382;
    wire N__10377;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10354;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10333;
    wire N__10332;
    wire N__10331;
    wire N__10330;
    wire N__10327;
    wire N__10326;
    wire N__10325;
    wire N__10318;
    wire N__10313;
    wire N__10310;
    wire N__10309;
    wire N__10308;
    wire N__10305;
    wire N__10300;
    wire N__10293;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10274;
    wire N__10269;
    wire N__10264;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9901;
    wire N__9898;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9874;
    wire N__9873;
    wire N__9868;
    wire N__9867;
    wire N__9864;
    wire N__9863;
    wire N__9862;
    wire N__9861;
    wire N__9860;
    wire N__9859;
    wire N__9856;
    wire N__9853;
    wire N__9852;
    wire N__9849;
    wire N__9844;
    wire N__9841;
    wire N__9836;
    wire N__9835;
    wire N__9834;
    wire N__9833;
    wire N__9832;
    wire N__9831;
    wire N__9830;
    wire N__9825;
    wire N__9822;
    wire N__9821;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9801;
    wire N__9796;
    wire N__9795;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9791;
    wire N__9790;
    wire N__9785;
    wire N__9782;
    wire N__9775;
    wire N__9770;
    wire N__9763;
    wire N__9756;
    wire N__9743;
    wire N__9742;
    wire N__9741;
    wire N__9740;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9732;
    wire N__9729;
    wire N__9728;
    wire N__9727;
    wire N__9722;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9711;
    wire N__9710;
    wire N__9709;
    wire N__9706;
    wire N__9701;
    wire N__9698;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9680;
    wire N__9677;
    wire N__9670;
    wire N__9667;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9578;
    wire N__9575;
    wire N__9574;
    wire N__9571;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9554;
    wire N__9551;
    wire N__9550;
    wire N__9549;
    wire N__9546;
    wire N__9541;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9496;
    wire N__9495;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9485;
    wire N__9484;
    wire N__9481;
    wire N__9476;
    wire N__9475;
    wire N__9474;
    wire N__9473;
    wire N__9472;
    wire N__9471;
    wire N__9470;
    wire N__9469;
    wire N__9466;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9448;
    wire N__9445;
    wire N__9440;
    wire N__9435;
    wire N__9430;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9406;
    wire N__9405;
    wire N__9404;
    wire N__9403;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9392;
    wire N__9391;
    wire N__9390;
    wire N__9385;
    wire N__9382;
    wire N__9381;
    wire N__9380;
    wire N__9379;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9365;
    wire N__9364;
    wire N__9361;
    wire N__9360;
    wire N__9359;
    wire N__9358;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9344;
    wire N__9339;
    wire N__9336;
    wire N__9331;
    wire N__9324;
    wire N__9321;
    wire N__9312;
    wire N__9309;
    wire N__9302;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9262;
    wire N__9261;
    wire N__9260;
    wire N__9259;
    wire N__9258;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9229;
    wire N__9228;
    wire N__9227;
    wire N__9224;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9212;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9200;
    wire N__9197;
    wire N__9192;
    wire N__9185;
    wire N__9182;
    wire N__9167;
    wire N__9164;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9142;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9136;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9122;
    wire N__9119;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9091;
    wire N__9090;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9017;
    wire N__9016;
    wire N__9015;
    wire N__9014;
    wire N__9013;
    wire N__9012;
    wire N__9011;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8990;
    wire N__8987;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8962;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8944;
    wire N__8943;
    wire N__8936;
    wire N__8929;
    wire N__8926;
    wire N__8919;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8897;
    wire N__8894;
    wire N__8893;
    wire N__8892;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8880;
    wire N__8877;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8745;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8701;
    wire N__8700;
    wire N__8697;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8681;
    wire N__8680;
    wire N__8679;
    wire N__8678;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8647;
    wire N__8646;
    wire N__8645;
    wire N__8644;
    wire N__8643;
    wire N__8642;
    wire N__8641;
    wire N__8640;
    wire N__8639;
    wire N__8636;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8574;
    wire N__8569;
    wire N__8566;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8551;
    wire N__8550;
    wire N__8547;
    wire N__8542;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8530;
    wire N__8529;
    wire N__8526;
    wire N__8521;
    wire N__8516;
    wire N__8513;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8462;
    wire N__8461;
    wire N__8460;
    wire N__8455;
    wire N__8454;
    wire N__8453;
    wire N__8452;
    wire N__8449;
    wire N__8448;
    wire N__8447;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8435;
    wire N__8432;
    wire N__8425;
    wire N__8414;
    wire N__8413;
    wire N__8412;
    wire N__8411;
    wire N__8410;
    wire N__8409;
    wire N__8406;
    wire N__8401;
    wire N__8396;
    wire N__8391;
    wire N__8384;
    wire N__8381;
    wire N__8380;
    wire N__8379;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8371;
    wire N__8368;
    wire N__8367;
    wire N__8364;
    wire N__8363;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8327;
    wire N__8326;
    wire N__8325;
    wire N__8324;
    wire N__8323;
    wire N__8322;
    wire N__8321;
    wire N__8320;
    wire N__8315;
    wire N__8312;
    wire N__8305;
    wire N__8300;
    wire N__8291;
    wire N__8290;
    wire N__8289;
    wire N__8288;
    wire N__8285;
    wire N__8284;
    wire N__8283;
    wire N__8282;
    wire N__8281;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8263;
    wire N__8258;
    wire N__8253;
    wire N__8240;
    wire N__8239;
    wire N__8238;
    wire N__8237;
    wire N__8230;
    wire N__8229;
    wire N__8228;
    wire N__8225;
    wire N__8224;
    wire N__8223;
    wire N__8222;
    wire N__8221;
    wire N__8220;
    wire N__8219;
    wire N__8218;
    wire N__8215;
    wire N__8210;
    wire N__8207;
    wire N__8198;
    wire N__8193;
    wire N__8190;
    wire N__8185;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8125;
    wire N__8120;
    wire N__8119;
    wire N__8116;
    wire N__8113;
    wire N__8108;
    wire N__8105;
    wire N__8104;
    wire N__8103;
    wire N__8102;
    wire N__8095;
    wire N__8092;
    wire N__8091;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8066;
    wire N__8065;
    wire N__8064;
    wire N__8063;
    wire N__8058;
    wire N__8053;
    wire N__8048;
    wire N__8047;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8029;
    wire N__8026;
    wire N__8021;
    wire N__8020;
    wire N__8019;
    wire N__8016;
    wire N__8011;
    wire N__8008;
    wire N__8003;
    wire N__8002;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7985;
    wire N__7984;
    wire N__7981;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7963;
    wire N__7962;
    wire N__7961;
    wire N__7958;
    wire N__7953;
    wire N__7950;
    wire N__7943;
    wire N__7942;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7899;
    wire N__7898;
    wire N__7895;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7887;
    wire N__7884;
    wire N__7883;
    wire N__7882;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7859;
    wire N__7844;
    wire N__7843;
    wire N__7842;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7834;
    wire N__7833;
    wire N__7832;
    wire N__7831;
    wire N__7830;
    wire N__7827;
    wire N__7824;
    wire N__7821;
    wire N__7818;
    wire N__7815;
    wire N__7810;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7798;
    wire N__7791;
    wire N__7788;
    wire N__7781;
    wire N__7778;
    wire N__7769;
    wire N__7766;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7754;
    wire N__7751;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7739;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7729;
    wire N__7724;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7673;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7661;
    wire N__7660;
    wire N__7655;
    wire N__7654;
    wire N__7651;
    wire N__7648;
    wire N__7645;
    wire N__7642;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7603;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7548;
    wire N__7545;
    wire N__7540;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7519;
    wire N__7516;
    wire N__7513;
    wire N__7512;
    wire N__7509;
    wire N__7504;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7388;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7291;
    wire N__7290;
    wire N__7289;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire VCCG0;
    wire GNDG0;
    wire port_clk_c;
    wire \this_vga_signals.N_469_0 ;
    wire port_rw_c_i;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire N_33;
    wire N_11;
    wire rgb_c_0;
    wire \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1Z0Z_9 ;
    wire \this_vga_signals.rgb_cnst_i_1Z0Z_3_cascade_ ;
    wire \this_vga_signals.rgb_cnst_i_1Z0Z_5 ;
    wire rgb_c_5;
    wire \this_vga_signals.M_vcounter_q_esr_RNIAV48E1Z0Z_9 ;
    wire rgb_c_3;
    wire \this_vga_signals.N_379_0 ;
    wire \this_vga_signals.M_vcounter_q_esr_RNIA99QRZ0Z_9_cascade_ ;
    wire rgb_c_1;
    wire \this_vga_signals.rgb_cnst_i_0_5 ;
    wire N_11_0;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire \this_vga_signals.if_i3_mux_2_0_cascade_ ;
    wire \this_vga_signals.if_m2_8_0_cascade_ ;
    wire \this_vga_signals.if_m8_0_ns_1 ;
    wire \this_vga_signals.if_m8_0_ns_1_cascade_ ;
    wire \this_vga_signals.g1_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ;
    wire \this_vga_signals.g1_cascade_ ;
    wire \this_vga_signals.if_m1_3_cascade_ ;
    wire \this_vga_signals.if_m1_3 ;
    wire \this_vga_signals.if_N_4_2 ;
    wire \this_vga_signals.if_i4_mux_0_1_cascade_ ;
    wire \this_vga_signals.vsync_1_0_a3_5_cascade_ ;
    wire this_vga_signals_vsync_1_i;
    wire \this_vga_signals.if_m13_0_ns_1_cascade_ ;
    wire \this_vga_signals.if_i3_mux_0_0_cascade_ ;
    wire \this_vga_signals.if_m13_0_ns_1 ;
    wire \this_vga_signals.if_i3_mux_0_0_0 ;
    wire \this_vga_signals.g2_1_cascade_ ;
    wire \this_vga_signals.g2_1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_1_1_0 ;
    wire \this_vga_signals.g0_5_0_1 ;
    wire \this_vga_signals.g3_0_2_0 ;
    wire \this_vga_signals.g2_cascade_ ;
    wire \this_vga_signals.g0_3_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_2_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_1_cascade_ ;
    wire \this_vga_signals.rgb_1_2_cascade_ ;
    wire \this_vga_signals.if_i3_mux_0_0 ;
    wire \this_vga_signals.if_i3_mux_2 ;
    wire \this_vga_signals.g1 ;
    wire \this_vga_signals.g3_0_2_cascade_ ;
    wire \this_vga_signals.if_N_3_0_i_1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_c_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_1 ;
    wire \this_vga_signals.if_N_15_mux ;
    wire \this_vga_signals.if_m13_ns_1_cascade_ ;
    wire \this_vga_signals.if_m13_ns ;
    wire \this_vga_signals.if_N_7 ;
    wire \this_vga_signals.d_N_9_0 ;
    wire \this_vga_signals.rgb_1_4_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIETZ0Z844 ;
    wire \this_vga_signals.d_N_5_0 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_i_x1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_2_N_2L1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.un11_address_0_5 ;
    wire \this_vga_signals.vsync_1_0_a3_4 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_9 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.d_N_8_0 ;
    wire \this_vga_signals.un11_address_1_5_cascade_ ;
    wire \this_vga_signals.g0_11_1 ;
    wire \this_vga_signals.g0_6_0 ;
    wire \this_vga_signals.g2_1_0_cascade_ ;
    wire \this_vga_signals.g3_cascade_ ;
    wire \this_vga_signals.g2_4_0 ;
    wire \this_vga_signals.mult1_un54_sum_c2_0 ;
    wire \this_vga_signals.mult1_un54_sum_i_1_cascade_ ;
    wire \this_vga_signals.un11_address_2_5_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_i_x0_3_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3 ;
    wire \this_vga_signals.if_N_3_0_i ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_c_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_c ;
    wire \this_vga_signals.mult1_un54_sum_ac0_1_0 ;
    wire \this_vga_signals.if_N_3_0_i_0 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_2 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_0 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_0 ;
    wire \this_vga_signals.g0_5_1 ;
    wire \this_vga_signals.mult1_un47_sum_c2_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_x1 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_x0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ;
    wire \this_vga_signals.g0_1 ;
    wire \this_vga_signals.un11_address_c4_i_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1_5_4_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABCZ0Z21 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_5_4_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.un11_address_c4_i ;
    wire \this_vga_signals.SUM_2_i_a4_1_0_3_cascade_ ;
    wire \this_vga_signals.un11_address_c5_a0_0_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPMZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_9_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_8_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_7_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.SUM_2_i_a4_0_a0_2_3_cascade_ ;
    wire \this_vga_signals.SUM_2_i_a4_a0_2_3 ;
    wire \this_vga_signals.SUM_2_i_1_0_3 ;
    wire \this_vga_signals.SUM_2_i_0_1_3 ;
    wire \this_vga_signals.SUM_2_i_0_3 ;
    wire bfn_11_23_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire bfn_11_24_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ;
    wire N_18;
    wire \this_vga_signals.hsync_1_i_0_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.N_469_0_g ;
    wire \this_vga_signals.N_608_g ;
    wire \this_vga_signals.N_381_0 ;
    wire \this_vga_signals.N_390_cascade_ ;
    wire \this_vga_signals.rgb_cnst_i_0_2_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_esr_RNIO6OD01Z0Z_9_cascade_ ;
    wire rgb_c_2;
    wire \this_vga_signals.g0_i_x2_1_0 ;
    wire \this_vga_signals.N_10_i ;
    wire \this_vga_signals.N_10_i_cascade_ ;
    wire \this_vga_signals.g0_i_x2_5_1 ;
    wire \this_vga_signals.if_N_13_i_i_1 ;
    wire \this_vga_signals.g4_0_0_cascade_ ;
    wire \this_vga_signals.g0_i_0_N_3L3 ;
    wire \this_vga_signals.N_3_1_0_1 ;
    wire \this_vga_signals.g0_i_x2_1_1_cascade_ ;
    wire this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_cascade_;
    wire \this_vga_signals.g0_i_x2_1_1 ;
    wire \this_vga_signals.g0_i_x1 ;
    wire \this_vga_signals.g0_i_x0_cascade_ ;
    wire this_vga_signals_un16_address_if_i1_mux_0_cascade_;
    wire \this_vga_signals.N_6_i_cascade_ ;
    wire \this_vga_signals.g1_1_0 ;
    wire \this_vga_signals.N_11_i ;
    wire \this_vga_signals.mult1_un40_sum_axb1 ;
    wire \this_vga_signals.g0_5_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_5_4 ;
    wire \this_vga_signals.g0_25_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_c ;
    wire \this_vga_signals.if_N_13_i_i_1_0_0_cascade_ ;
    wire \this_vga_signals.g2_0_0_0 ;
    wire \this_vga_signals.N_371_0 ;
    wire rgb_c_4;
    wire \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0 ;
    wire \this_vga_signals.un11_address_0_7_cascade_ ;
    wire \this_vga_signals.SUM_2 ;
    wire \this_vga_signals.g0_3_0 ;
    wire \this_vga_signals.N_28_0_cascade_ ;
    wire \this_vga_signals.N_42_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_esr_RNIVV6F6Z0Z_9 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.rgb297_i_a3_0_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.SUM_2_i_a4_0_a0_2_3 ;
    wire \this_vga_signals.N_33_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire \this_vga_signals.N_49 ;
    wire \this_vga_signals.N_33_0_cascade_ ;
    wire \this_vga_signals.CO0_i_i ;
    wire \this_vga_signals.N_45_cascade_ ;
    wire N_23_0;
    wire N_23_0_cascade_;
    wire \this_pixel_clock.M_counter_q_i_1 ;
    wire bfn_12_24_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_12_25_0_;
    wire \this_vga_signals.N_22 ;
    wire \this_vga_signals.g1_0_0_2_cascade_ ;
    wire \this_vga_signals.N_21 ;
    wire \this_vga_signals.g0_i_x2_1 ;
    wire \this_vga_signals.g4_1 ;
    wire \this_vga_signals.g0_1_0_cascade_ ;
    wire \this_vga_signals.g0_i_x2_5 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_cascade_ ;
    wire \this_vga_signals.N_9_1_0 ;
    wire \this_vga_signals.g1_5 ;
    wire \this_vga_signals.N_6 ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_0_0_1_cascade_ ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.g2_0_1_0 ;
    wire \this_vga_signals.g0_i_x2_2 ;
    wire \this_vga_signals.g0_i_0_N_4L5_cascade_ ;
    wire \this_vga_signals.g0_i_0_N_5L7 ;
    wire \this_vga_signals.if_i4_mux_0_0_0_1 ;
    wire \this_vga_signals.N_6_i ;
    wire \this_vga_signals.g1_1_2 ;
    wire \this_vga_signals.g1_4_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.g0_i_0_N_2L1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_vcounter_d_1_sqmuxa_i_a3_1 ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.if_N_8_i_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axb1 ;
    wire \this_vga_signals.mult1_un89_sum_c3 ;
    wire \this_vga_signals.mult1_un82_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_2 ;
    wire \this_vga_signals.mult1_un82_sum_c2_0 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0_0_cascade_ ;
    wire \this_vga_signals.if_N_9_0_0 ;
    wire \this_vga_signals.mult1_un68_sum_axb1 ;
    wire \this_vga_signals.SUM_3_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.N_34 ;
    wire \this_vga_signals.N_34_cascade_ ;
    wire \this_vga_signals.SUM_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c2_0 ;
    wire \this_vga_signals.N_469_1 ;
    wire debug_0_i;
    wire \this_vga_signals.rgb_cnst_i_a5_0_0Z0Z_3 ;
    wire M_this_vram_read_data_0;
    wire \this_vga_signals.mult1_un61_sum_axb1 ;
    wire \this_vga_signals.if_m3_5_cascade_ ;
    wire \this_vga_signals.if_N_3_i ;
    wire \this_vga_signals.if_m5_4_cascade_ ;
    wire \this_vga_signals.g1_1_4 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_1 ;
    wire \this_vga_signals.mult1_un68_sum_axb2_0_1_cascade_ ;
    wire \this_vga_signals.g1_1_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0 ;
    wire \this_vga_signals.g0_1_0_0_cascade_ ;
    wire \this_vga_signals.g4_0 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_d_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_ac0_4 ;
    wire \this_vga_signals.g0_i_o2_0_0_x2_0_cascade_ ;
    wire \this_vga_signals.N_16 ;
    wire \this_vga_signals.mult1_un54_sum_i_1 ;
    wire \this_vga_signals.if_N_1_i_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_0 ;
    wire N_401;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_2 ;
    wire M_this_vga_signals_address_4;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire M_counter_q_RNIJR071_1;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire M_counter_q_RNIQR4I2_1;
    wire \this_vga_signals.rgb_bmZ0Z_1 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_5 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.if_N_13_i_i_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_0 ;
    wire \this_vga_signals.if_N_16_i_0 ;
    wire \this_vga_signals.g0_1_N_5L8 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_0 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_d ;
    wire \this_vga_signals.g0_1_N_3L3 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.g0_1_N_6L11_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c2_0 ;
    wire \this_vga_signals.g0_1_N_7L13 ;
    wire \this_vga_signals.g0_1_N_8L15_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.mult1_un68_sum_axb2_0 ;
    wire \this_vga_signals.mult1_un68_sum_c2_0_0_cascade_ ;
    wire \this_vga_signals.if_N_6_3_0 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0_cascade_ ;
    wire M_this_vga_signals_address_8;
    wire N_349_0_cascade_;
    wire port_enb_c;
    wire \this_delay_clk.M_this_delay_clk_out_0 ;
    wire debug_0;
    wire port_rw_c;
    wire port_address_c_7;
    wire debug_0_cascade_;
    wire this_start_data_delay_M_last_q;
    wire M_current_address_qZ0Z_0;
    wire N_312_0;
    wire M_current_address_q_RNO_1Z0Z_0;
    wire bfn_15_21_0_;
    wire un1_M_current_address_q_cry_0;
    wire un1_M_current_address_q_cry_1;
    wire un1_M_current_address_q_cry_2;
    wire un1_M_current_address_q_cry_3;
    wire un1_M_current_address_q_cry_4;
    wire un1_M_current_address_q_cry_5;
    wire un1_M_current_address_q_cry_6;
    wire un1_M_current_address_q_cry_7;
    wire bfn_15_22_0_;
    wire un1_M_current_address_q_cry_8;
    wire un1_M_current_address_q_cry_9;
    wire un1_M_current_address_q_cry_10;
    wire un1_M_current_address_q_cry_11;
    wire un1_M_current_address_q_cry_12;
    wire \this_pixel_clock.M_counter_qZ0Z_0 ;
    wire M_this_vram_read_data_3;
    wire \this_vga_signals.rgb_bmZ0Z_0 ;
    wire \this_vga_signals.rgb_bmZ0Z_2 ;
    wire m7_am_cascade_;
    wire m7_ns;
    wire m28_cascade_;
    wire m32_am_cascade_;
    wire m7_bm;
    wire m32_bm;
    wire m32_ns;
    wire rgb_2_4;
    wire m29;
    wire \this_vga_signals.rgb_bmZ0Z_3 ;
    wire port_data_c_5;
    wire N_413_cascade_;
    wire M_current_address_q_RNO_1Z0Z_12;
    wire N_411;
    wire M_current_address_q_RNO_1Z0Z_10;
    wire M_current_address_qZ0Z_10;
    wire N_404;
    wire M_current_address_q_RNO_1Z0Z_3;
    wire M_current_address_qZ0Z_3;
    wire M_current_address_q_RNO_1Z0Z_5;
    wire N_406;
    wire M_current_address_qZ0Z_5;
    wire N_402_cascade_;
    wire M_current_address_q_RNO_1Z0Z_1;
    wire M_current_address_qZ0Z_1;
    wire M_current_address_q_RNO_1Z0Z_8;
    wire N_409;
    wire M_current_address_qZ0Z_8;
    wire N_412;
    wire M_current_address_q_RNO_1Z0Z_11;
    wire port_data_c_4;
    wire M_current_address_q_RNO_1Z0Z_9;
    wire M_this_vram_read_data_1;
    wire bfn_17_16_0_;
    wire rgb291_cry_0;
    wire rgb291_cry_1;
    wire CONSTANT_ONE_NET;
    wire rgb291_cry_2;
    wire rgb291;
    wire \this_vga_signals.rgb_1_sqmuxa ;
    wire mem_radreg_RNIMTEJ4_0_11;
    wire mem_radreg_RNIETEJ4_0_11;
    wire m44_cascade_;
    wire m22_am_cascade_;
    wire m22_ns;
    wire m22_bm;
    wire m24;
    wire m40_cascade_;
    wire m41;
    wire m10;
    wire rgb_1_axb_0_cascade_;
    wire m15;
    wire rgb_1_0;
    wire m37;
    wire m19;
    wire rgb_1_axb_0;
    wire a0_b_0;
    wire m46_am_cascade_;
    wire m46_bm;
    wire rgb_2_5;
    wire N_352;
    wire N_408_cascade_;
    wire M_current_address_q_RNO_1Z0Z_7;
    wire M_current_address_qZ0Z_7;
    wire N_405;
    wire M_current_address_q_RNO_1Z0Z_4;
    wire M_current_address_qZ0Z_4;
    wire M_state_q_ns_0_a3_0_2_0;
    wire N_351;
    wire N_403_cascade_;
    wire M_current_address_q_RNO_1Z0Z_2;
    wire M_current_address_qZ0Z_2;
    wire M_current_address_q_RNO_1Z0Z_13;
    wire M_state_qZ0Z_1;
    wire N_407_cascade_;
    wire M_current_address_q_RNO_1Z0Z_6;
    wire M_current_address_qZ0Z_6;
    wire M_this_reset_cond_out_0;
    wire M_current_address_qZ0Z_9;
    wire N_410;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0 ;
    wire M_this_vga_signals_address_5;
    wire mem_radreg_RNIETEJ4_11;
    wire M_this_vram_read_data_2;
    wire this_vram_mem_radreg_11;
    wire mem_radreg_RNIMTEJ4_11;
    wire m14;
    wire rgb_1_cry_0_0_c_RNOZ0;
    wire bfn_18_20_0_;
    wire M_vcounter_q_esr_RNIB9J4TN_9;
    wire M_vcounter_q_esr_RNICJRF0D_9;
    wire rgb_1_cry_0;
    wire rgb_1_cry_1;
    wire rgb_1_cry_2;
    wire rgb_1_6;
    wire this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3;
    wire rgb_1_cry_0_0_c_RNOZ0Z_0;
    wire M_vcounter_q_esr_RNI1H9RHL_9;
    wire rgb_1_3;
    wire rgb_1_4;
    wire rgb_1_5;
    wire rgb_1_6_THRU_CO;
    wire m36;
    wire port_address_c_0;
    wire port_address_c_1;
    wire M_state_q_ns_0_a3_0_1_1;
    wire port_data_c_1;
    wire M_this_vram_write_data_1;
    wire N_349_0;
    wire port_data_c_6;
    wire M_state_qZ0Z_0;
    wire N_414;
    wire this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1;
    wire this_vga_signals_un16_address_if_i1_mux_0;
    wire M_this_vga_signals_address_10;
    wire rgbZ0Z_1_cascade_;
    wire M_vcounter_q_esr_RNI2RH6LA_9;
    wire rgbZ0Z_1;
    wire M_vcounter_q_esr_RNIVLNKSA_9;
    wire \this_vga_signals.mult1_un68_sum_axbxc3 ;
    wire M_this_vga_signals_address_3;
    wire port_data_c_0;
    wire M_this_vram_write_data_0;
    wire \this_vga_signals.SUM_3_1 ;
    wire M_this_vga_signals_address_6;
    wire \this_vram.mem_WE_12 ;
    wire \this_vga_signals.rgb_1_2 ;
    wire \this_vram.mem_WE_8 ;
    wire \this_vram.mem_out_bus0_3 ;
    wire \this_vram.mem_out_bus4_3 ;
    wire \this_vram.mem_N_88 ;
    wire \this_vram.mem_mem_0_1_RNISOI11Z0Z_0 ;
    wire \this_vram.mem_N_105 ;
    wire \this_vram.mem_WE_10 ;
    wire \this_vram.mem_WE_14 ;
    wire this_vram_mem_N_112;
    wire \this_vga_signals.rgb_1_4 ;
    wire clk_0_c_g;
    wire port_data_c_3;
    wire M_this_vram_write_data_3;
    wire \this_vram.mem_out_bus4_1 ;
    wire \this_vram.mem_out_bus0_1 ;
    wire \this_vram.mem_out_bus2_1 ;
    wire \this_vram.mem_out_bus6_1 ;
    wire \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0 ;
    wire \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_91 ;
    wire \this_vram.mem_out_bus5_1 ;
    wire \this_vram.mem_out_bus1_1 ;
    wire \this_vram.mem_mem_1_0_RNISSK11Z0Z_0 ;
    wire \this_vram.mem_out_bus3_1 ;
    wire \this_vram.mem_out_bus7_1 ;
    wire \this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ;
    wire \this_vram.mem_out_bus1_0 ;
    wire \this_vram.mem_out_bus5_0 ;
    wire \this_vram.mem_out_bus2_3 ;
    wire \this_vram.mem_out_bus6_3 ;
    wire \this_vram.mem_mem_2_1_RNI01N11Z0Z_0 ;
    wire \this_vram.mem_out_bus0_2 ;
    wire \this_vram.mem_out_bus4_2 ;
    wire \this_vram.mem_out_bus1_2 ;
    wire \this_vram.mem_out_bus5_2 ;
    wire \this_vram.mem_out_bus2_2 ;
    wire \this_vram.mem_out_bus6_2 ;
    wire \this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_ ;
    wire \this_vram.mem_mem_0_1_RNISOIZ0Z11 ;
    wire \this_vram.mem_N_98 ;
    wire \this_vram.mem_out_bus1_3 ;
    wire \this_vram.mem_out_bus5_3 ;
    wire \this_vram.mem_out_bus3_3 ;
    wire \this_vram.mem_out_bus7_3 ;
    wire \this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_ ;
    wire \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0 ;
    wire \this_vram.mem_N_102 ;
    wire \this_vram.mem_mem_1_0_RNISSKZ0Z11 ;
    wire this_vram_mem_N_109;
    wire \this_vram.mem_out_bus3_2 ;
    wire \this_vram.mem_out_bus7_2 ;
    wire \this_vram.mem_mem_1_1_RNIUSKZ0Z11 ;
    wire \this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_ ;
    wire \this_vram.mem_radregZ0Z_12 ;
    wire \this_vram.mem_N_95 ;
    wire \this_vram.mem_out_bus6_0 ;
    wire \this_vram.mem_out_bus2_0 ;
    wire \this_vram.mem_mem_2_0_RNIU0NZ0Z11 ;
    wire \this_vram.mem_out_bus7_0 ;
    wire \this_vram.mem_out_bus3_0 ;
    wire \this_vram.mem_mem_3_0_RNI05PZ0Z11 ;
    wire \this_vram.mem_out_bus0_0 ;
    wire \this_vram.mem_out_bus4_0 ;
    wire \this_vram.mem_radregZ0Z_13 ;
    wire \this_vram.mem_mem_0_0_RNIQOIZ0Z11 ;
    wire \this_vram.mem_WE_6 ;
    wire port_data_c_2;
    wire M_this_vram_write_data_2;
    wire \this_vram.mem_WE_4 ;
    wire \this_vram.mem_WE_0 ;
    wire M_current_address_qZ0Z_12;
    wire M_current_address_qZ0Z_13;
    wire M_current_address_qZ0Z_11;
    wire M_this_vram_write_en_0_sqmuxa;
    wire \this_vram.mem_WE_2 ;
    wire M_this_vga_signals_address_2;
    wire \this_vga_signals.if_m2_5_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0 ;
    wire M_this_vga_signals_address_9;
    wire \this_vga_signals.N_9_0 ;
    wire \this_vga_signals.mult1_un75_sum_c3_0 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_1 ;
    wire M_this_vga_signals_address_1;
    wire port_address_c_5;
    wire port_address_c_6;
    wire port_address_c_2;
    wire port_address_c_3;
    wire port_address_c_4;
    wire M_state_q_ns_0_a3_0_0_1_0;
    wire M_state_q_ns_0_a3_0_0_0;
    wire _gnd_net_;

    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,\this_vram.mem_out_bus0_1 ,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,\this_vram.mem_out_bus0_0 ,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__16019,N__20438,N__12020,N__10076,N__17483,N__15089,N__11852,N__17747,N__19205,N__20123,N__10259}),
            .WADDR({N__13640,N__15224,N__13973,N__14816,N__15458,N__13367,N__14675,N__13508,N__15710,N__13241,N__12731}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,N__16574,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__17582,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .RCLKE(),
            .RCLK(N__18179),
            .RE(N__14434),
            .WCLKE(N__18436),
            .WCLK(N__18180),
            .WE(N__14418));
    defparam \this_vram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,\this_vram.mem_out_bus0_3 ,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,\this_vram.mem_out_bus0_2 ,dangling_wire_55,dangling_wire_56,dangling_wire_57}),
            .RADDR({N__16013,N__20432,N__12014,N__10070,N__17477,N__15083,N__11846,N__17741,N__19199,N__20117,N__10253}),
            .WADDR({N__13634,N__15218,N__13967,N__14810,N__15452,N__13361,N__14669,N__13502,N__15704,N__13235,N__12725}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,N__18008,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,N__19727,dangling_wire_85,dangling_wire_86,dangling_wire_87}),
            .RCLKE(),
            .RCLK(N__18181),
            .RE(N__14413),
            .WCLKE(N__18437),
            .WCLK(N__18182),
            .WE(N__14414));
    defparam \this_vram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,\this_vram.mem_out_bus1_1 ,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,\this_vram.mem_out_bus1_0 ,dangling_wire_99,dangling_wire_100,dangling_wire_101}),
            .RADDR({N__16007,N__20426,N__12008,N__10064,N__17471,N__15077,N__11840,N__17735,N__19193,N__20111,N__10247}),
            .WADDR({N__13628,N__15212,N__13961,N__14804,N__15446,N__13355,N__14663,N__13496,N__15698,N__13229,N__12719}),
            .MASK({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .WDATA({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__16570,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__17577,dangling_wire_129,dangling_wire_130,dangling_wire_131}),
            .RCLKE(),
            .RCLK(N__18183),
            .RE(N__14412),
            .WCLKE(N__17375),
            .WCLK(N__18184),
            .WE(N__14386));
    defparam \this_vram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,\this_vram.mem_out_bus1_3 ,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,\this_vram.mem_out_bus1_2 ,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .RADDR({N__16001,N__20420,N__12002,N__10058,N__17465,N__15071,N__11834,N__17729,N__19187,N__20105,N__10241}),
            .WADDR({N__13622,N__15206,N__13955,N__14798,N__15440,N__13349,N__14657,N__13490,N__15692,N__13223,N__12713}),
            .MASK({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161}),
            .WDATA({dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__18004,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,N__19723,dangling_wire_173,dangling_wire_174,dangling_wire_175}),
            .RCLKE(),
            .RCLK(N__18185),
            .RE(N__14369),
            .WCLKE(N__17371),
            .WCLK(N__18186),
            .WE(N__14385));
    defparam \this_vram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,\this_vram.mem_out_bus2_1 ,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,\this_vram.mem_out_bus2_0 ,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .RADDR({N__15995,N__20414,N__11996,N__10052,N__17459,N__15065,N__11828,N__17723,N__19181,N__20099,N__10235}),
            .WADDR({N__13616,N__15200,N__13949,N__14792,N__15434,N__13343,N__14651,N__13484,N__15686,N__13217,N__12707}),
            .MASK({dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205}),
            .WDATA({dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,N__16546,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,N__17565,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .RCLKE(),
            .RCLK(N__18188),
            .RE(N__14327),
            .WCLKE(N__18464),
            .WCLK(N__18187),
            .WE(N__14306));
    defparam \this_vram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,\this_vram.mem_out_bus2_3 ,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,\this_vram.mem_out_bus2_2 ,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .RADDR({N__15989,N__20408,N__11990,N__10046,N__17453,N__15059,N__11822,N__17717,N__19175,N__20093,N__10229}),
            .WADDR({N__13610,N__15194,N__13943,N__14786,N__15428,N__13337,N__14645,N__13478,N__15680,N__13211,N__12701}),
            .MASK({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .WDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,N__17996,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,N__19715,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RCLKE(),
            .RCLK(N__18190),
            .RE(N__14311),
            .WCLKE(N__18460),
            .WCLK(N__18191),
            .WE(N__14305));
    defparam \this_vram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,\this_vram.mem_out_bus3_1 ,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,\this_vram.mem_out_bus3_0 ,dangling_wire_275,dangling_wire_276,dangling_wire_277}),
            .RADDR({N__15983,N__20402,N__11984,N__10040,N__17447,N__15053,N__11816,N__17711,N__19169,N__20087,N__10223}),
            .WADDR({N__13604,N__15188,N__13937,N__14780,N__15422,N__13331,N__14639,N__13472,N__15674,N__13205,N__12695}),
            .MASK({dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293}),
            .WDATA({dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,N__16557,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,N__17581,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .RCLKE(),
            .RCLK(N__18198),
            .RE(N__14223),
            .WCLKE(N__17243),
            .WCLK(N__18199),
            .WE(N__14172));
    defparam \this_vram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,\this_vram.mem_out_bus3_3 ,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,\this_vram.mem_out_bus3_2 ,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .RADDR({N__15977,N__20396,N__11978,N__10034,N__17441,N__15047,N__11810,N__17705,N__19163,N__20081,N__10217}),
            .WADDR({N__13598,N__15182,N__13931,N__14774,N__15416,N__13325,N__14633,N__13466,N__15668,N__13199,N__12689}),
            .MASK({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .WDATA({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,N__17982,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,N__19701,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .RCLKE(),
            .RCLK(N__18206),
            .RE(N__14307),
            .WCLKE(N__17242),
            .WCLK(N__18207),
            .WE(N__14278));
    defparam \this_vram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,\this_vram.mem_out_bus4_1 ,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,\this_vram.mem_out_bus4_0 ,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .RADDR({N__15971,N__20390,N__11972,N__10028,N__17435,N__15041,N__11804,N__17699,N__19157,N__20075,N__10211}),
            .WADDR({N__13592,N__15176,N__13925,N__14768,N__15410,N__13319,N__14627,N__13460,N__15662,N__13193,N__12683}),
            .MASK({dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381}),
            .WDATA({dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,N__16547,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,N__17573,dangling_wire_393,dangling_wire_394,dangling_wire_395}),
            .RCLKE(),
            .RCLK(N__18210),
            .RE(N__14368),
            .WCLKE(N__19789),
            .WCLK(N__18211),
            .WE(N__14338));
    defparam \this_vram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,\this_vram.mem_out_bus4_3 ,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,\this_vram.mem_out_bus4_2 ,dangling_wire_407,dangling_wire_408,dangling_wire_409}),
            .RADDR({N__15965,N__20384,N__11966,N__10022,N__17429,N__15035,N__11798,N__17693,N__19151,N__20069,N__10205}),
            .WADDR({N__13586,N__15170,N__13919,N__14762,N__15404,N__13313,N__14621,N__13454,N__15656,N__13187,N__12677}),
            .MASK({dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425}),
            .WDATA({dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,N__17963,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,N__19661,dangling_wire_437,dangling_wire_438,dangling_wire_439}),
            .RCLKE(),
            .RCLK(N__18218),
            .RE(N__14351),
            .WCLKE(N__19793),
            .WCLK(N__18219),
            .WE(N__14339));
    defparam \this_vram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,\this_vram.mem_out_bus5_1 ,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,\this_vram.mem_out_bus5_0 ,dangling_wire_451,dangling_wire_452,dangling_wire_453}),
            .RADDR({N__15959,N__20378,N__11960,N__10016,N__17423,N__15029,N__11792,N__17687,N__19145,N__20063,N__10199}),
            .WADDR({N__13580,N__15164,N__13913,N__14756,N__15398,N__13307,N__14615,N__13448,N__15650,N__13181,N__12671}),
            .MASK({dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469}),
            .WDATA({dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,N__16507,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,N__17519,dangling_wire_481,dangling_wire_482,dangling_wire_483}),
            .RCLKE(),
            .RCLK(N__18224),
            .RE(N__14398),
            .WCLKE(N__19642),
            .WCLK(N__18225),
            .WE(N__14388));
    defparam \this_vram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,\this_vram.mem_out_bus5_3 ,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,\this_vram.mem_out_bus5_2 ,dangling_wire_495,dangling_wire_496,dangling_wire_497}),
            .RADDR({N__15953,N__20372,N__11954,N__10010,N__17417,N__15023,N__11786,N__17681,N__19139,N__20057,N__10193}),
            .WADDR({N__13574,N__15158,N__13907,N__14750,N__15392,N__13301,N__14609,N__13442,N__15644,N__13175,N__12665}),
            .MASK({dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513}),
            .WDATA({dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,N__17964,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,N__19694,dangling_wire_525,dangling_wire_526,dangling_wire_527}),
            .RCLKE(),
            .RCLK(N__18228),
            .RE(N__14399),
            .WCLKE(N__19643),
            .WCLK(N__18229),
            .WE(N__14389));
    defparam \this_vram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,\this_vram.mem_out_bus6_1 ,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,\this_vram.mem_out_bus6_0 ,dangling_wire_539,dangling_wire_540,dangling_wire_541}),
            .RADDR({N__15947,N__20366,N__11948,N__10004,N__17411,N__15017,N__11780,N__17675,N__19133,N__20051,N__10187}),
            .WADDR({N__13568,N__15152,N__13901,N__14744,N__15386,N__13295,N__14603,N__13436,N__15638,N__13169,N__12659}),
            .MASK({dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557}),
            .WDATA({dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,N__16542,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,N__17555,dangling_wire_569,dangling_wire_570,dangling_wire_571}),
            .RCLKE(),
            .RCLK(N__18232),
            .RE(N__14426),
            .WCLKE(N__19222),
            .WCLK(N__18233),
            .WE(N__14271));
    defparam \this_vram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,\this_vram.mem_out_bus6_3 ,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,\this_vram.mem_out_bus6_2 ,dangling_wire_583,dangling_wire_584,dangling_wire_585}),
            .RADDR({N__15941,N__20360,N__11942,N__9998,N__17405,N__15011,N__11774,N__17669,N__19127,N__20045,N__10181}),
            .WADDR({N__13562,N__15146,N__13895,N__14738,N__15380,N__13289,N__14597,N__13430,N__15632,N__13163,N__12653}),
            .MASK({dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601}),
            .WDATA({dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,N__17992,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,N__19711,dangling_wire_613,dangling_wire_614,dangling_wire_615}),
            .RCLKE(),
            .RCLK(N__18234),
            .RE(N__14430),
            .WCLKE(N__19226),
            .WCLK(N__18235),
            .WE(N__14419));
    defparam \this_vram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,\this_vram.mem_out_bus7_1 ,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,\this_vram.mem_out_bus7_0 ,dangling_wire_627,dangling_wire_628,dangling_wire_629}),
            .RADDR({N__15935,N__20354,N__11936,N__9992,N__17399,N__15005,N__11768,N__17663,N__19121,N__20039,N__10175}),
            .WADDR({N__13556,N__15140,N__13889,N__14732,N__15374,N__13283,N__14591,N__13424,N__15626,N__13157,N__12647}),
            .MASK({dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645}),
            .WDATA({dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,N__16556,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,N__17572,dangling_wire_657,dangling_wire_658,dangling_wire_659}),
            .RCLKE(),
            .RCLK(N__18236),
            .RE(N__14440),
            .WCLKE(N__19621),
            .WCLK(N__18237),
            .WE(N__14435));
    defparam \this_vram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,\this_vram.mem_out_bus7_3 ,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,\this_vram.mem_out_bus7_2 ,dangling_wire_671,dangling_wire_672,dangling_wire_673}),
            .RADDR({N__15929,N__20348,N__11930,N__9986,N__17393,N__14999,N__11762,N__17657,N__19115,N__20033,N__10169}),
            .WADDR({N__13550,N__15134,N__13883,N__14726,N__15368,N__13277,N__14585,N__13418,N__15620,N__13151,N__12641}),
            .MASK({dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689}),
            .WDATA({dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,N__18003,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,N__19722,dangling_wire_701,dangling_wire_702,dangling_wire_703}),
            .RCLKE(),
            .RCLK(N__18238),
            .RE(N__14441),
            .WCLKE(N__19625),
            .WCLK(N__18239),
            .WE(N__14436));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__20796),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__20798),
            .DIN(N__20797),
            .DOUT(N__20796),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__20798),
            .PADOUT(N__20797),
            .PADIN(N__20796),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_iopad (
            .OE(N__20787),
            .DIN(N__20786),
            .DOUT(N__20785),
            .PACKAGEPIN(debug));
    defparam debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_preio (
            .PADOEN(N__20787),
            .PADOUT(N__20786),
            .PADIN(N__20785),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10457),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__20778),
            .DIN(N__20777),
            .DOUT(N__20776),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__20778),
            .PADOUT(N__20777),
            .PADIN(N__20776),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7100),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__20769),
            .DIN(N__20768),
            .DOUT(N__20767),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__20769),
            .PADOUT(N__20768),
            .PADIN(N__20767),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8726),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_0_iopad (
            .OE(N__20760),
            .DIN(N__20759),
            .DOUT(N__20758),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_0_preio (
            .PADOEN(N__20760),
            .PADOUT(N__20759),
            .PADIN(N__20758),
            .CLOCKENABLE(),
            .DIN0(port_address_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_1_iopad (
            .OE(N__20751),
            .DIN(N__20750),
            .DOUT(N__20749),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_1_preio (
            .PADOEN(N__20751),
            .PADOUT(N__20750),
            .PADIN(N__20749),
            .CLOCKENABLE(),
            .DIN0(port_address_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_2_iopad (
            .OE(N__20742),
            .DIN(N__20741),
            .DOUT(N__20740),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_2_preio (
            .PADOEN(N__20742),
            .PADOUT(N__20741),
            .PADIN(N__20740),
            .CLOCKENABLE(),
            .DIN0(port_address_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_3_iopad (
            .OE(N__20733),
            .DIN(N__20732),
            .DOUT(N__20731),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_3_preio (
            .PADOEN(N__20733),
            .PADOUT(N__20732),
            .PADIN(N__20731),
            .CLOCKENABLE(),
            .DIN0(port_address_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_4_iopad (
            .OE(N__20724),
            .DIN(N__20723),
            .DOUT(N__20722),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_4_preio (
            .PADOEN(N__20724),
            .PADOUT(N__20723),
            .PADIN(N__20722),
            .CLOCKENABLE(),
            .DIN0(port_address_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_5_iopad (
            .OE(N__20715),
            .DIN(N__20714),
            .DOUT(N__20713),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_5_preio (
            .PADOEN(N__20715),
            .PADOUT(N__20714),
            .PADIN(N__20713),
            .CLOCKENABLE(),
            .DIN0(port_address_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_6_iopad (
            .OE(N__20706),
            .DIN(N__20705),
            .DOUT(N__20704),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_6_preio (
            .PADOEN(N__20706),
            .PADOUT(N__20705),
            .PADIN(N__20704),
            .CLOCKENABLE(),
            .DIN0(port_address_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_7_iopad (
            .OE(N__20697),
            .DIN(N__20696),
            .DOUT(N__20695),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_7_preio (
            .PADOEN(N__20697),
            .PADOUT(N__20696),
            .PADIN(N__20695),
            .CLOCKENABLE(),
            .DIN0(port_address_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__20688),
            .DIN(N__20687),
            .DOUT(N__20686),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__20688),
            .PADOUT(N__20687),
            .PADIN(N__20686),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__20679),
            .DIN(N__20678),
            .DOUT(N__20677),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__20679),
            .PADOUT(N__20678),
            .PADIN(N__20677),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__20670),
            .DIN(N__20669),
            .DOUT(N__20668),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__20670),
            .PADOUT(N__20669),
            .PADIN(N__20668),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__20661),
            .DIN(N__20660),
            .DOUT(N__20659),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__20661),
            .PADOUT(N__20660),
            .PADIN(N__20659),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__20652),
            .DIN(N__20651),
            .DOUT(N__20650),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__20652),
            .PADOUT(N__20651),
            .PADIN(N__20650),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__20643),
            .DIN(N__20642),
            .DOUT(N__20641),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__20643),
            .PADOUT(N__20642),
            .PADIN(N__20641),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__20634),
            .DIN(N__20633),
            .DOUT(N__20632),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__20634),
            .PADOUT(N__20633),
            .PADIN(N__20632),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__20625),
            .DIN(N__20624),
            .DOUT(N__20623),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__20625),
            .PADOUT(N__20624),
            .PADIN(N__20623),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__20616),
            .DIN(N__20615),
            .DOUT(N__20614),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__20616),
            .PADOUT(N__20615),
            .PADIN(N__20614),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7034),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__20607),
            .DIN(N__20606),
            .DOUT(N__20605),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__20607),
            .PADOUT(N__20606),
            .PADIN(N__20605),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14387),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__20598),
            .DIN(N__20597),
            .DOUT(N__20596),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__20598),
            .PADOUT(N__20597),
            .PADIN(N__20596),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__20589),
            .DIN(N__20588),
            .DOUT(N__20587),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__20589),
            .PADOUT(N__20588),
            .PADIN(N__20587),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7160),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_ibuf_iopad (
            .OE(N__20580),
            .DIN(N__20579),
            .DOUT(N__20578),
            .PACKAGEPIN(port_rw));
    defparam port_rw_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_rw_ibuf_preio (
            .PADOEN(N__20580),
            .PADOUT(N__20579),
            .PADIN(N__20578),
            .CLOCKENABLE(),
            .DIN0(port_rw_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__20571),
            .DIN(N__20570),
            .DOUT(N__20569),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__20571),
            .PADOUT(N__20570),
            .PADIN(N__20569),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7082),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__20562),
            .DIN(N__20561),
            .DOUT(N__20560),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__20562),
            .PADOUT(N__20561),
            .PADIN(N__20560),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7178),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__20553),
            .DIN(N__20552),
            .DOUT(N__20551),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__20553),
            .PADOUT(N__20552),
            .PADIN(N__20551),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8828),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__20544),
            .DIN(N__20543),
            .DOUT(N__20542),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__20544),
            .PADOUT(N__20543),
            .PADIN(N__20542),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7211),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__20535),
            .DIN(N__20534),
            .DOUT(N__20533),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__20535),
            .PADOUT(N__20534),
            .PADIN(N__20533),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__9032),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__20526),
            .DIN(N__20525),
            .DOUT(N__20524),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__20526),
            .PADOUT(N__20525),
            .PADIN(N__20524),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7238),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__20517),
            .DIN(N__20516),
            .DOUT(N__20515),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__20517),
            .PADOUT(N__20516),
            .PADIN(N__20515),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__20508),
            .DIN(N__20507),
            .DOUT(N__20506),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__20508),
            .PADOUT(N__20507),
            .PADIN(N__20506),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7091),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__20499),
            .DIN(N__20498),
            .DOUT(N__20497),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__20499),
            .PADOUT(N__20498),
            .PADIN(N__20497),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7343),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__4987 (
            .O(N__20480),
            .I(N__20477));
    LocalMux I__4986 (
            .O(N__20477),
            .I(N__20474));
    Span12Mux_s10_h I__4985 (
            .O(N__20474),
            .I(N__20470));
    InMux I__4984 (
            .O(N__20473),
            .I(N__20467));
    Span12Mux_v I__4983 (
            .O(N__20470),
            .I(N__20464));
    LocalMux I__4982 (
            .O(N__20467),
            .I(\this_vga_signals.if_m2_5_0 ));
    Odrv12 I__4981 (
            .O(N__20464),
            .I(\this_vga_signals.if_m2_5_0 ));
    InMux I__4980 (
            .O(N__20459),
            .I(N__20456));
    LocalMux I__4979 (
            .O(N__20456),
            .I(N__20453));
    Span12Mux_h I__4978 (
            .O(N__20453),
            .I(N__20450));
    Span12Mux_v I__4977 (
            .O(N__20450),
            .I(N__20446));
    InMux I__4976 (
            .O(N__20449),
            .I(N__20443));
    Odrv12 I__4975 (
            .O(N__20446),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__4974 (
            .O(N__20443),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    CascadeMux I__4973 (
            .O(N__20438),
            .I(N__20435));
    CascadeBuf I__4972 (
            .O(N__20435),
            .I(N__20432));
    CascadeMux I__4971 (
            .O(N__20432),
            .I(N__20429));
    CascadeBuf I__4970 (
            .O(N__20429),
            .I(N__20426));
    CascadeMux I__4969 (
            .O(N__20426),
            .I(N__20423));
    CascadeBuf I__4968 (
            .O(N__20423),
            .I(N__20420));
    CascadeMux I__4967 (
            .O(N__20420),
            .I(N__20417));
    CascadeBuf I__4966 (
            .O(N__20417),
            .I(N__20414));
    CascadeMux I__4965 (
            .O(N__20414),
            .I(N__20411));
    CascadeBuf I__4964 (
            .O(N__20411),
            .I(N__20408));
    CascadeMux I__4963 (
            .O(N__20408),
            .I(N__20405));
    CascadeBuf I__4962 (
            .O(N__20405),
            .I(N__20402));
    CascadeMux I__4961 (
            .O(N__20402),
            .I(N__20399));
    CascadeBuf I__4960 (
            .O(N__20399),
            .I(N__20396));
    CascadeMux I__4959 (
            .O(N__20396),
            .I(N__20393));
    CascadeBuf I__4958 (
            .O(N__20393),
            .I(N__20390));
    CascadeMux I__4957 (
            .O(N__20390),
            .I(N__20387));
    CascadeBuf I__4956 (
            .O(N__20387),
            .I(N__20384));
    CascadeMux I__4955 (
            .O(N__20384),
            .I(N__20381));
    CascadeBuf I__4954 (
            .O(N__20381),
            .I(N__20378));
    CascadeMux I__4953 (
            .O(N__20378),
            .I(N__20375));
    CascadeBuf I__4952 (
            .O(N__20375),
            .I(N__20372));
    CascadeMux I__4951 (
            .O(N__20372),
            .I(N__20369));
    CascadeBuf I__4950 (
            .O(N__20369),
            .I(N__20366));
    CascadeMux I__4949 (
            .O(N__20366),
            .I(N__20363));
    CascadeBuf I__4948 (
            .O(N__20363),
            .I(N__20360));
    CascadeMux I__4947 (
            .O(N__20360),
            .I(N__20357));
    CascadeBuf I__4946 (
            .O(N__20357),
            .I(N__20354));
    CascadeMux I__4945 (
            .O(N__20354),
            .I(N__20351));
    CascadeBuf I__4944 (
            .O(N__20351),
            .I(N__20348));
    CascadeMux I__4943 (
            .O(N__20348),
            .I(N__20345));
    InMux I__4942 (
            .O(N__20345),
            .I(N__20342));
    LocalMux I__4941 (
            .O(N__20342),
            .I(M_this_vga_signals_address_9));
    InMux I__4940 (
            .O(N__20339),
            .I(N__20335));
    InMux I__4939 (
            .O(N__20338),
            .I(N__20326));
    LocalMux I__4938 (
            .O(N__20335),
            .I(N__20320));
    InMux I__4937 (
            .O(N__20334),
            .I(N__20317));
    InMux I__4936 (
            .O(N__20333),
            .I(N__20314));
    InMux I__4935 (
            .O(N__20332),
            .I(N__20311));
    InMux I__4934 (
            .O(N__20331),
            .I(N__20305));
    InMux I__4933 (
            .O(N__20330),
            .I(N__20302));
    InMux I__4932 (
            .O(N__20329),
            .I(N__20299));
    LocalMux I__4931 (
            .O(N__20326),
            .I(N__20295));
    InMux I__4930 (
            .O(N__20325),
            .I(N__20292));
    InMux I__4929 (
            .O(N__20324),
            .I(N__20286));
    InMux I__4928 (
            .O(N__20323),
            .I(N__20283));
    Sp12to4 I__4927 (
            .O(N__20320),
            .I(N__20280));
    LocalMux I__4926 (
            .O(N__20317),
            .I(N__20273));
    LocalMux I__4925 (
            .O(N__20314),
            .I(N__20273));
    LocalMux I__4924 (
            .O(N__20311),
            .I(N__20273));
    InMux I__4923 (
            .O(N__20310),
            .I(N__20270));
    InMux I__4922 (
            .O(N__20309),
            .I(N__20267));
    InMux I__4921 (
            .O(N__20308),
            .I(N__20263));
    LocalMux I__4920 (
            .O(N__20305),
            .I(N__20257));
    LocalMux I__4919 (
            .O(N__20302),
            .I(N__20257));
    LocalMux I__4918 (
            .O(N__20299),
            .I(N__20254));
    InMux I__4917 (
            .O(N__20298),
            .I(N__20251));
    Span4Mux_v I__4916 (
            .O(N__20295),
            .I(N__20246));
    LocalMux I__4915 (
            .O(N__20292),
            .I(N__20246));
    InMux I__4914 (
            .O(N__20291),
            .I(N__20243));
    CascadeMux I__4913 (
            .O(N__20290),
            .I(N__20240));
    InMux I__4912 (
            .O(N__20289),
            .I(N__20237));
    LocalMux I__4911 (
            .O(N__20286),
            .I(N__20232));
    LocalMux I__4910 (
            .O(N__20283),
            .I(N__20232));
    Span12Mux_v I__4909 (
            .O(N__20280),
            .I(N__20225));
    Span12Mux_s7_v I__4908 (
            .O(N__20273),
            .I(N__20225));
    LocalMux I__4907 (
            .O(N__20270),
            .I(N__20225));
    LocalMux I__4906 (
            .O(N__20267),
            .I(N__20222));
    InMux I__4905 (
            .O(N__20266),
            .I(N__20219));
    LocalMux I__4904 (
            .O(N__20263),
            .I(N__20216));
    InMux I__4903 (
            .O(N__20262),
            .I(N__20213));
    Span4Mux_h I__4902 (
            .O(N__20257),
            .I(N__20210));
    Span4Mux_v I__4901 (
            .O(N__20254),
            .I(N__20201));
    LocalMux I__4900 (
            .O(N__20251),
            .I(N__20201));
    Span4Mux_h I__4899 (
            .O(N__20246),
            .I(N__20201));
    LocalMux I__4898 (
            .O(N__20243),
            .I(N__20201));
    InMux I__4897 (
            .O(N__20240),
            .I(N__20198));
    LocalMux I__4896 (
            .O(N__20237),
            .I(N__20191));
    Sp12to4 I__4895 (
            .O(N__20232),
            .I(N__20191));
    Span12Mux_h I__4894 (
            .O(N__20225),
            .I(N__20191));
    Span12Mux_v I__4893 (
            .O(N__20222),
            .I(N__20182));
    LocalMux I__4892 (
            .O(N__20219),
            .I(N__20182));
    Span12Mux_h I__4891 (
            .O(N__20216),
            .I(N__20182));
    LocalMux I__4890 (
            .O(N__20213),
            .I(N__20182));
    Span4Mux_h I__4889 (
            .O(N__20210),
            .I(N__20177));
    Span4Mux_h I__4888 (
            .O(N__20201),
            .I(N__20177));
    LocalMux I__4887 (
            .O(N__20198),
            .I(\this_vga_signals.N_9_0 ));
    Odrv12 I__4886 (
            .O(N__20191),
            .I(\this_vga_signals.N_9_0 ));
    Odrv12 I__4885 (
            .O(N__20182),
            .I(\this_vga_signals.N_9_0 ));
    Odrv4 I__4884 (
            .O(N__20177),
            .I(\this_vga_signals.N_9_0 ));
    InMux I__4883 (
            .O(N__20168),
            .I(N__20164));
    InMux I__4882 (
            .O(N__20167),
            .I(N__20161));
    LocalMux I__4881 (
            .O(N__20164),
            .I(N__20158));
    LocalMux I__4880 (
            .O(N__20161),
            .I(N__20155));
    Sp12to4 I__4879 (
            .O(N__20158),
            .I(N__20150));
    Sp12to4 I__4878 (
            .O(N__20155),
            .I(N__20150));
    Span12Mux_s9_v I__4877 (
            .O(N__20150),
            .I(N__20145));
    InMux I__4876 (
            .O(N__20149),
            .I(N__20140));
    InMux I__4875 (
            .O(N__20148),
            .I(N__20140));
    Odrv12 I__4874 (
            .O(N__20145),
            .I(\this_vga_signals.mult1_un75_sum_c3_0 ));
    LocalMux I__4873 (
            .O(N__20140),
            .I(\this_vga_signals.mult1_un75_sum_c3_0 ));
    InMux I__4872 (
            .O(N__20135),
            .I(N__20132));
    LocalMux I__4871 (
            .O(N__20132),
            .I(N__20129));
    Span12Mux_h I__4870 (
            .O(N__20129),
            .I(N__20126));
    Odrv12 I__4869 (
            .O(N__20126),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1 ));
    CascadeMux I__4868 (
            .O(N__20123),
            .I(N__20120));
    CascadeBuf I__4867 (
            .O(N__20120),
            .I(N__20117));
    CascadeMux I__4866 (
            .O(N__20117),
            .I(N__20114));
    CascadeBuf I__4865 (
            .O(N__20114),
            .I(N__20111));
    CascadeMux I__4864 (
            .O(N__20111),
            .I(N__20108));
    CascadeBuf I__4863 (
            .O(N__20108),
            .I(N__20105));
    CascadeMux I__4862 (
            .O(N__20105),
            .I(N__20102));
    CascadeBuf I__4861 (
            .O(N__20102),
            .I(N__20099));
    CascadeMux I__4860 (
            .O(N__20099),
            .I(N__20096));
    CascadeBuf I__4859 (
            .O(N__20096),
            .I(N__20093));
    CascadeMux I__4858 (
            .O(N__20093),
            .I(N__20090));
    CascadeBuf I__4857 (
            .O(N__20090),
            .I(N__20087));
    CascadeMux I__4856 (
            .O(N__20087),
            .I(N__20084));
    CascadeBuf I__4855 (
            .O(N__20084),
            .I(N__20081));
    CascadeMux I__4854 (
            .O(N__20081),
            .I(N__20078));
    CascadeBuf I__4853 (
            .O(N__20078),
            .I(N__20075));
    CascadeMux I__4852 (
            .O(N__20075),
            .I(N__20072));
    CascadeBuf I__4851 (
            .O(N__20072),
            .I(N__20069));
    CascadeMux I__4850 (
            .O(N__20069),
            .I(N__20066));
    CascadeBuf I__4849 (
            .O(N__20066),
            .I(N__20063));
    CascadeMux I__4848 (
            .O(N__20063),
            .I(N__20060));
    CascadeBuf I__4847 (
            .O(N__20060),
            .I(N__20057));
    CascadeMux I__4846 (
            .O(N__20057),
            .I(N__20054));
    CascadeBuf I__4845 (
            .O(N__20054),
            .I(N__20051));
    CascadeMux I__4844 (
            .O(N__20051),
            .I(N__20048));
    CascadeBuf I__4843 (
            .O(N__20048),
            .I(N__20045));
    CascadeMux I__4842 (
            .O(N__20045),
            .I(N__20042));
    CascadeBuf I__4841 (
            .O(N__20042),
            .I(N__20039));
    CascadeMux I__4840 (
            .O(N__20039),
            .I(N__20036));
    CascadeBuf I__4839 (
            .O(N__20036),
            .I(N__20033));
    CascadeMux I__4838 (
            .O(N__20033),
            .I(N__20030));
    InMux I__4837 (
            .O(N__20030),
            .I(N__20027));
    LocalMux I__4836 (
            .O(N__20027),
            .I(M_this_vga_signals_address_1));
    InMux I__4835 (
            .O(N__20024),
            .I(N__20021));
    LocalMux I__4834 (
            .O(N__20021),
            .I(port_address_c_5));
    InMux I__4833 (
            .O(N__20018),
            .I(N__20015));
    LocalMux I__4832 (
            .O(N__20015),
            .I(N__20012));
    Span4Mux_v I__4831 (
            .O(N__20012),
            .I(N__20009));
    Odrv4 I__4830 (
            .O(N__20009),
            .I(port_address_c_6));
    InMux I__4829 (
            .O(N__20006),
            .I(N__20003));
    LocalMux I__4828 (
            .O(N__20003),
            .I(N__20000));
    Span12Mux_s10_h I__4827 (
            .O(N__20000),
            .I(N__19997));
    Odrv12 I__4826 (
            .O(N__19997),
            .I(port_address_c_2));
    InMux I__4825 (
            .O(N__19994),
            .I(N__19991));
    LocalMux I__4824 (
            .O(N__19991),
            .I(N__19988));
    Span12Mux_v I__4823 (
            .O(N__19988),
            .I(N__19985));
    Odrv12 I__4822 (
            .O(N__19985),
            .I(port_address_c_3));
    CascadeMux I__4821 (
            .O(N__19982),
            .I(N__19979));
    InMux I__4820 (
            .O(N__19979),
            .I(N__19976));
    LocalMux I__4819 (
            .O(N__19976),
            .I(port_address_c_4));
    InMux I__4818 (
            .O(N__19973),
            .I(N__19970));
    LocalMux I__4817 (
            .O(N__19970),
            .I(N__19967));
    Odrv4 I__4816 (
            .O(N__19967),
            .I(M_state_q_ns_0_a3_0_0_1_0));
    CascadeMux I__4815 (
            .O(N__19964),
            .I(N__19960));
    CascadeMux I__4814 (
            .O(N__19963),
            .I(N__19957));
    InMux I__4813 (
            .O(N__19960),
            .I(N__19954));
    InMux I__4812 (
            .O(N__19957),
            .I(N__19951));
    LocalMux I__4811 (
            .O(N__19954),
            .I(N__19946));
    LocalMux I__4810 (
            .O(N__19951),
            .I(N__19946));
    Span12Mux_h I__4809 (
            .O(N__19946),
            .I(N__19943));
    Span12Mux_h I__4808 (
            .O(N__19943),
            .I(N__19940));
    Odrv12 I__4807 (
            .O(N__19940),
            .I(M_state_q_ns_0_a3_0_0_0));
    InMux I__4806 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__4805 (
            .O(N__19934),
            .I(\this_vram.mem_mem_2_0_RNIU0NZ0Z11 ));
    InMux I__4804 (
            .O(N__19931),
            .I(N__19928));
    LocalMux I__4803 (
            .O(N__19928),
            .I(N__19925));
    Sp12to4 I__4802 (
            .O(N__19925),
            .I(N__19922));
    Span12Mux_v I__4801 (
            .O(N__19922),
            .I(N__19919));
    Odrv12 I__4800 (
            .O(N__19919),
            .I(\this_vram.mem_out_bus7_0 ));
    InMux I__4799 (
            .O(N__19916),
            .I(N__19913));
    LocalMux I__4798 (
            .O(N__19913),
            .I(N__19910));
    Odrv4 I__4797 (
            .O(N__19910),
            .I(\this_vram.mem_out_bus3_0 ));
    InMux I__4796 (
            .O(N__19907),
            .I(N__19904));
    LocalMux I__4795 (
            .O(N__19904),
            .I(\this_vram.mem_mem_3_0_RNI05PZ0Z11 ));
    InMux I__4794 (
            .O(N__19901),
            .I(N__19898));
    LocalMux I__4793 (
            .O(N__19898),
            .I(N__19895));
    Sp12to4 I__4792 (
            .O(N__19895),
            .I(N__19892));
    Span12Mux_v I__4791 (
            .O(N__19892),
            .I(N__19889));
    Odrv12 I__4790 (
            .O(N__19889),
            .I(\this_vram.mem_out_bus0_0 ));
    InMux I__4789 (
            .O(N__19886),
            .I(N__19883));
    LocalMux I__4788 (
            .O(N__19883),
            .I(\this_vram.mem_out_bus4_0 ));
    CascadeMux I__4787 (
            .O(N__19880),
            .I(N__19873));
    InMux I__4786 (
            .O(N__19879),
            .I(N__19863));
    InMux I__4785 (
            .O(N__19878),
            .I(N__19863));
    InMux I__4784 (
            .O(N__19877),
            .I(N__19854));
    InMux I__4783 (
            .O(N__19876),
            .I(N__19854));
    InMux I__4782 (
            .O(N__19873),
            .I(N__19854));
    InMux I__4781 (
            .O(N__19872),
            .I(N__19854));
    InMux I__4780 (
            .O(N__19871),
            .I(N__19851));
    InMux I__4779 (
            .O(N__19870),
            .I(N__19844));
    InMux I__4778 (
            .O(N__19869),
            .I(N__19844));
    InMux I__4777 (
            .O(N__19868),
            .I(N__19844));
    LocalMux I__4776 (
            .O(N__19863),
            .I(N__19834));
    LocalMux I__4775 (
            .O(N__19854),
            .I(N__19834));
    LocalMux I__4774 (
            .O(N__19851),
            .I(N__19834));
    LocalMux I__4773 (
            .O(N__19844),
            .I(N__19831));
    InMux I__4772 (
            .O(N__19843),
            .I(N__19824));
    InMux I__4771 (
            .O(N__19842),
            .I(N__19824));
    InMux I__4770 (
            .O(N__19841),
            .I(N__19824));
    Span4Mux_v I__4769 (
            .O(N__19834),
            .I(N__19814));
    Span4Mux_h I__4768 (
            .O(N__19831),
            .I(N__19814));
    LocalMux I__4767 (
            .O(N__19824),
            .I(N__19814));
    InMux I__4766 (
            .O(N__19823),
            .I(N__19809));
    InMux I__4765 (
            .O(N__19822),
            .I(N__19809));
    InMux I__4764 (
            .O(N__19821),
            .I(N__19806));
    Odrv4 I__4763 (
            .O(N__19814),
            .I(\this_vram.mem_radregZ0Z_13 ));
    LocalMux I__4762 (
            .O(N__19809),
            .I(\this_vram.mem_radregZ0Z_13 ));
    LocalMux I__4761 (
            .O(N__19806),
            .I(\this_vram.mem_radregZ0Z_13 ));
    InMux I__4760 (
            .O(N__19799),
            .I(N__19796));
    LocalMux I__4759 (
            .O(N__19796),
            .I(\this_vram.mem_mem_0_0_RNIQOIZ0Z11 ));
    CEMux I__4758 (
            .O(N__19793),
            .I(N__19790));
    LocalMux I__4757 (
            .O(N__19790),
            .I(N__19786));
    CEMux I__4756 (
            .O(N__19789),
            .I(N__19783));
    Span4Mux_v I__4755 (
            .O(N__19786),
            .I(N__19780));
    LocalMux I__4754 (
            .O(N__19783),
            .I(N__19777));
    Odrv4 I__4753 (
            .O(N__19780),
            .I(\this_vram.mem_WE_6 ));
    Odrv4 I__4752 (
            .O(N__19777),
            .I(\this_vram.mem_WE_6 ));
    CascadeMux I__4751 (
            .O(N__19772),
            .I(N__19768));
    InMux I__4750 (
            .O(N__19771),
            .I(N__19764));
    InMux I__4749 (
            .O(N__19768),
            .I(N__19761));
    InMux I__4748 (
            .O(N__19767),
            .I(N__19758));
    LocalMux I__4747 (
            .O(N__19764),
            .I(N__19753));
    LocalMux I__4746 (
            .O(N__19761),
            .I(N__19753));
    LocalMux I__4745 (
            .O(N__19758),
            .I(N__19750));
    Span4Mux_v I__4744 (
            .O(N__19753),
            .I(N__19747));
    Span4Mux_v I__4743 (
            .O(N__19750),
            .I(N__19744));
    Sp12to4 I__4742 (
            .O(N__19747),
            .I(N__19741));
    Sp12to4 I__4741 (
            .O(N__19744),
            .I(N__19738));
    Span12Mux_h I__4740 (
            .O(N__19741),
            .I(N__19735));
    Span12Mux_h I__4739 (
            .O(N__19738),
            .I(N__19732));
    Odrv12 I__4738 (
            .O(N__19735),
            .I(port_data_c_2));
    Odrv12 I__4737 (
            .O(N__19732),
            .I(port_data_c_2));
    InMux I__4736 (
            .O(N__19727),
            .I(N__19724));
    LocalMux I__4735 (
            .O(N__19724),
            .I(N__19719));
    InMux I__4734 (
            .O(N__19723),
            .I(N__19716));
    InMux I__4733 (
            .O(N__19722),
            .I(N__19712));
    Span4Mux_h I__4732 (
            .O(N__19719),
            .I(N__19708));
    LocalMux I__4731 (
            .O(N__19716),
            .I(N__19705));
    InMux I__4730 (
            .O(N__19715),
            .I(N__19702));
    LocalMux I__4729 (
            .O(N__19712),
            .I(N__19698));
    InMux I__4728 (
            .O(N__19711),
            .I(N__19695));
    Span4Mux_v I__4727 (
            .O(N__19708),
            .I(N__19689));
    Span4Mux_h I__4726 (
            .O(N__19705),
            .I(N__19689));
    LocalMux I__4725 (
            .O(N__19702),
            .I(N__19686));
    InMux I__4724 (
            .O(N__19701),
            .I(N__19683));
    Span4Mux_v I__4723 (
            .O(N__19698),
            .I(N__19678));
    LocalMux I__4722 (
            .O(N__19695),
            .I(N__19678));
    InMux I__4721 (
            .O(N__19694),
            .I(N__19675));
    Span4Mux_v I__4720 (
            .O(N__19689),
            .I(N__19670));
    Span4Mux_h I__4719 (
            .O(N__19686),
            .I(N__19670));
    LocalMux I__4718 (
            .O(N__19683),
            .I(N__19667));
    Span4Mux_v I__4717 (
            .O(N__19678),
            .I(N__19662));
    LocalMux I__4716 (
            .O(N__19675),
            .I(N__19662));
    Span4Mux_v I__4715 (
            .O(N__19670),
            .I(N__19656));
    Span4Mux_h I__4714 (
            .O(N__19667),
            .I(N__19656));
    Span4Mux_v I__4713 (
            .O(N__19662),
            .I(N__19653));
    InMux I__4712 (
            .O(N__19661),
            .I(N__19650));
    Odrv4 I__4711 (
            .O(N__19656),
            .I(M_this_vram_write_data_2));
    Odrv4 I__4710 (
            .O(N__19653),
            .I(M_this_vram_write_data_2));
    LocalMux I__4709 (
            .O(N__19650),
            .I(M_this_vram_write_data_2));
    CEMux I__4708 (
            .O(N__19643),
            .I(N__19639));
    CEMux I__4707 (
            .O(N__19642),
            .I(N__19636));
    LocalMux I__4706 (
            .O(N__19639),
            .I(N__19631));
    LocalMux I__4705 (
            .O(N__19636),
            .I(N__19631));
    Span4Mux_v I__4704 (
            .O(N__19631),
            .I(N__19628));
    Odrv4 I__4703 (
            .O(N__19628),
            .I(\this_vram.mem_WE_4 ));
    CEMux I__4702 (
            .O(N__19625),
            .I(N__19622));
    LocalMux I__4701 (
            .O(N__19622),
            .I(N__19618));
    CEMux I__4700 (
            .O(N__19621),
            .I(N__19615));
    Span4Mux_s2_v I__4699 (
            .O(N__19618),
            .I(N__19610));
    LocalMux I__4698 (
            .O(N__19615),
            .I(N__19610));
    Span4Mux_v I__4697 (
            .O(N__19610),
            .I(N__19607));
    Span4Mux_v I__4696 (
            .O(N__19607),
            .I(N__19604));
    Odrv4 I__4695 (
            .O(N__19604),
            .I(\this_vram.mem_WE_0 ));
    CascadeMux I__4694 (
            .O(N__19601),
            .I(N__19598));
    InMux I__4693 (
            .O(N__19598),
            .I(N__19592));
    InMux I__4692 (
            .O(N__19597),
            .I(N__19589));
    InMux I__4691 (
            .O(N__19596),
            .I(N__19586));
    InMux I__4690 (
            .O(N__19595),
            .I(N__19583));
    LocalMux I__4689 (
            .O(N__19592),
            .I(N__19576));
    LocalMux I__4688 (
            .O(N__19589),
            .I(N__19571));
    LocalMux I__4687 (
            .O(N__19586),
            .I(N__19571));
    LocalMux I__4686 (
            .O(N__19583),
            .I(N__19568));
    InMux I__4685 (
            .O(N__19582),
            .I(N__19563));
    InMux I__4684 (
            .O(N__19581),
            .I(N__19563));
    InMux I__4683 (
            .O(N__19580),
            .I(N__19560));
    InMux I__4682 (
            .O(N__19579),
            .I(N__19557));
    Span4Mux_v I__4681 (
            .O(N__19576),
            .I(N__19552));
    Span4Mux_v I__4680 (
            .O(N__19571),
            .I(N__19552));
    Span4Mux_v I__4679 (
            .O(N__19568),
            .I(N__19549));
    LocalMux I__4678 (
            .O(N__19563),
            .I(N__19546));
    LocalMux I__4677 (
            .O(N__19560),
            .I(N__19541));
    LocalMux I__4676 (
            .O(N__19557),
            .I(N__19538));
    Span4Mux_h I__4675 (
            .O(N__19552),
            .I(N__19535));
    Span4Mux_v I__4674 (
            .O(N__19549),
            .I(N__19530));
    Span4Mux_h I__4673 (
            .O(N__19546),
            .I(N__19530));
    InMux I__4672 (
            .O(N__19545),
            .I(N__19527));
    InMux I__4671 (
            .O(N__19544),
            .I(N__19524));
    Span12Mux_s10_h I__4670 (
            .O(N__19541),
            .I(N__19519));
    Span12Mux_v I__4669 (
            .O(N__19538),
            .I(N__19519));
    Span4Mux_h I__4668 (
            .O(N__19535),
            .I(N__19516));
    Span4Mux_h I__4667 (
            .O(N__19530),
            .I(N__19513));
    LocalMux I__4666 (
            .O(N__19527),
            .I(M_current_address_qZ0Z_12));
    LocalMux I__4665 (
            .O(N__19524),
            .I(M_current_address_qZ0Z_12));
    Odrv12 I__4664 (
            .O(N__19519),
            .I(M_current_address_qZ0Z_12));
    Odrv4 I__4663 (
            .O(N__19516),
            .I(M_current_address_qZ0Z_12));
    Odrv4 I__4662 (
            .O(N__19513),
            .I(M_current_address_qZ0Z_12));
    CascadeMux I__4661 (
            .O(N__19502),
            .I(N__19493));
    CascadeMux I__4660 (
            .O(N__19501),
            .I(N__19490));
    CascadeMux I__4659 (
            .O(N__19500),
            .I(N__19487));
    CascadeMux I__4658 (
            .O(N__19499),
            .I(N__19484));
    CascadeMux I__4657 (
            .O(N__19498),
            .I(N__19481));
    CascadeMux I__4656 (
            .O(N__19497),
            .I(N__19477));
    InMux I__4655 (
            .O(N__19496),
            .I(N__19472));
    InMux I__4654 (
            .O(N__19493),
            .I(N__19472));
    InMux I__4653 (
            .O(N__19490),
            .I(N__19469));
    InMux I__4652 (
            .O(N__19487),
            .I(N__19466));
    InMux I__4651 (
            .O(N__19484),
            .I(N__19463));
    InMux I__4650 (
            .O(N__19481),
            .I(N__19459));
    InMux I__4649 (
            .O(N__19480),
            .I(N__19454));
    InMux I__4648 (
            .O(N__19477),
            .I(N__19454));
    LocalMux I__4647 (
            .O(N__19472),
            .I(N__19451));
    LocalMux I__4646 (
            .O(N__19469),
            .I(N__19448));
    LocalMux I__4645 (
            .O(N__19466),
            .I(N__19443));
    LocalMux I__4644 (
            .O(N__19463),
            .I(N__19443));
    InMux I__4643 (
            .O(N__19462),
            .I(N__19440));
    LocalMux I__4642 (
            .O(N__19459),
            .I(N__19433));
    LocalMux I__4641 (
            .O(N__19454),
            .I(N__19433));
    Span4Mux_v I__4640 (
            .O(N__19451),
            .I(N__19433));
    Span4Mux_h I__4639 (
            .O(N__19448),
            .I(N__19427));
    Span4Mux_v I__4638 (
            .O(N__19443),
            .I(N__19427));
    LocalMux I__4637 (
            .O(N__19440),
            .I(N__19424));
    Span4Mux_v I__4636 (
            .O(N__19433),
            .I(N__19421));
    InMux I__4635 (
            .O(N__19432),
            .I(N__19418));
    Span4Mux_h I__4634 (
            .O(N__19427),
            .I(N__19415));
    Span4Mux_h I__4633 (
            .O(N__19424),
            .I(N__19410));
    Span4Mux_h I__4632 (
            .O(N__19421),
            .I(N__19410));
    LocalMux I__4631 (
            .O(N__19418),
            .I(M_current_address_qZ0Z_13));
    Odrv4 I__4630 (
            .O(N__19415),
            .I(M_current_address_qZ0Z_13));
    Odrv4 I__4629 (
            .O(N__19410),
            .I(M_current_address_qZ0Z_13));
    InMux I__4628 (
            .O(N__19403),
            .I(N__19398));
    InMux I__4627 (
            .O(N__19402),
            .I(N__19395));
    CascadeMux I__4626 (
            .O(N__19401),
            .I(N__19387));
    LocalMux I__4625 (
            .O(N__19398),
            .I(N__19383));
    LocalMux I__4624 (
            .O(N__19395),
            .I(N__19379));
    InMux I__4623 (
            .O(N__19394),
            .I(N__19376));
    InMux I__4622 (
            .O(N__19393),
            .I(N__19373));
    InMux I__4621 (
            .O(N__19392),
            .I(N__19370));
    InMux I__4620 (
            .O(N__19391),
            .I(N__19367));
    InMux I__4619 (
            .O(N__19390),
            .I(N__19364));
    InMux I__4618 (
            .O(N__19387),
            .I(N__19359));
    InMux I__4617 (
            .O(N__19386),
            .I(N__19359));
    Span4Mux_h I__4616 (
            .O(N__19383),
            .I(N__19356));
    InMux I__4615 (
            .O(N__19382),
            .I(N__19353));
    Span4Mux_h I__4614 (
            .O(N__19379),
            .I(N__19350));
    LocalMux I__4613 (
            .O(N__19376),
            .I(N__19341));
    LocalMux I__4612 (
            .O(N__19373),
            .I(N__19341));
    LocalMux I__4611 (
            .O(N__19370),
            .I(N__19341));
    LocalMux I__4610 (
            .O(N__19367),
            .I(N__19341));
    LocalMux I__4609 (
            .O(N__19364),
            .I(N__19336));
    LocalMux I__4608 (
            .O(N__19359),
            .I(N__19336));
    Span4Mux_h I__4607 (
            .O(N__19356),
            .I(N__19333));
    LocalMux I__4606 (
            .O(N__19353),
            .I(N__19328));
    Span4Mux_h I__4605 (
            .O(N__19350),
            .I(N__19328));
    Span12Mux_h I__4604 (
            .O(N__19341),
            .I(N__19325));
    Odrv12 I__4603 (
            .O(N__19336),
            .I(M_current_address_qZ0Z_11));
    Odrv4 I__4602 (
            .O(N__19333),
            .I(M_current_address_qZ0Z_11));
    Odrv4 I__4601 (
            .O(N__19328),
            .I(M_current_address_qZ0Z_11));
    Odrv12 I__4600 (
            .O(N__19325),
            .I(M_current_address_qZ0Z_11));
    InMux I__4599 (
            .O(N__19316),
            .I(N__19306));
    InMux I__4598 (
            .O(N__19315),
            .I(N__19301));
    InMux I__4597 (
            .O(N__19314),
            .I(N__19301));
    InMux I__4596 (
            .O(N__19313),
            .I(N__19298));
    InMux I__4595 (
            .O(N__19312),
            .I(N__19292));
    InMux I__4594 (
            .O(N__19311),
            .I(N__19292));
    InMux I__4593 (
            .O(N__19310),
            .I(N__19289));
    InMux I__4592 (
            .O(N__19309),
            .I(N__19286));
    LocalMux I__4591 (
            .O(N__19306),
            .I(N__19283));
    LocalMux I__4590 (
            .O(N__19301),
            .I(N__19278));
    LocalMux I__4589 (
            .O(N__19298),
            .I(N__19278));
    InMux I__4588 (
            .O(N__19297),
            .I(N__19273));
    LocalMux I__4587 (
            .O(N__19292),
            .I(N__19266));
    LocalMux I__4586 (
            .O(N__19289),
            .I(N__19266));
    LocalMux I__4585 (
            .O(N__19286),
            .I(N__19266));
    Span4Mux_v I__4584 (
            .O(N__19283),
            .I(N__19261));
    Span4Mux_v I__4583 (
            .O(N__19278),
            .I(N__19261));
    InMux I__4582 (
            .O(N__19277),
            .I(N__19258));
    InMux I__4581 (
            .O(N__19276),
            .I(N__19255));
    LocalMux I__4580 (
            .O(N__19273),
            .I(N__19252));
    Span12Mux_h I__4579 (
            .O(N__19266),
            .I(N__19248));
    Sp12to4 I__4578 (
            .O(N__19261),
            .I(N__19241));
    LocalMux I__4577 (
            .O(N__19258),
            .I(N__19241));
    LocalMux I__4576 (
            .O(N__19255),
            .I(N__19241));
    Span4Mux_h I__4575 (
            .O(N__19252),
            .I(N__19238));
    InMux I__4574 (
            .O(N__19251),
            .I(N__19235));
    Odrv12 I__4573 (
            .O(N__19248),
            .I(M_this_vram_write_en_0_sqmuxa));
    Odrv12 I__4572 (
            .O(N__19241),
            .I(M_this_vram_write_en_0_sqmuxa));
    Odrv4 I__4571 (
            .O(N__19238),
            .I(M_this_vram_write_en_0_sqmuxa));
    LocalMux I__4570 (
            .O(N__19235),
            .I(M_this_vram_write_en_0_sqmuxa));
    CEMux I__4569 (
            .O(N__19226),
            .I(N__19223));
    LocalMux I__4568 (
            .O(N__19223),
            .I(N__19219));
    CEMux I__4567 (
            .O(N__19222),
            .I(N__19216));
    Span4Mux_v I__4566 (
            .O(N__19219),
            .I(N__19211));
    LocalMux I__4565 (
            .O(N__19216),
            .I(N__19211));
    Span4Mux_v I__4564 (
            .O(N__19211),
            .I(N__19208));
    Odrv4 I__4563 (
            .O(N__19208),
            .I(\this_vram.mem_WE_2 ));
    CascadeMux I__4562 (
            .O(N__19205),
            .I(N__19202));
    CascadeBuf I__4561 (
            .O(N__19202),
            .I(N__19199));
    CascadeMux I__4560 (
            .O(N__19199),
            .I(N__19196));
    CascadeBuf I__4559 (
            .O(N__19196),
            .I(N__19193));
    CascadeMux I__4558 (
            .O(N__19193),
            .I(N__19190));
    CascadeBuf I__4557 (
            .O(N__19190),
            .I(N__19187));
    CascadeMux I__4556 (
            .O(N__19187),
            .I(N__19184));
    CascadeBuf I__4555 (
            .O(N__19184),
            .I(N__19181));
    CascadeMux I__4554 (
            .O(N__19181),
            .I(N__19178));
    CascadeBuf I__4553 (
            .O(N__19178),
            .I(N__19175));
    CascadeMux I__4552 (
            .O(N__19175),
            .I(N__19172));
    CascadeBuf I__4551 (
            .O(N__19172),
            .I(N__19169));
    CascadeMux I__4550 (
            .O(N__19169),
            .I(N__19166));
    CascadeBuf I__4549 (
            .O(N__19166),
            .I(N__19163));
    CascadeMux I__4548 (
            .O(N__19163),
            .I(N__19160));
    CascadeBuf I__4547 (
            .O(N__19160),
            .I(N__19157));
    CascadeMux I__4546 (
            .O(N__19157),
            .I(N__19154));
    CascadeBuf I__4545 (
            .O(N__19154),
            .I(N__19151));
    CascadeMux I__4544 (
            .O(N__19151),
            .I(N__19148));
    CascadeBuf I__4543 (
            .O(N__19148),
            .I(N__19145));
    CascadeMux I__4542 (
            .O(N__19145),
            .I(N__19142));
    CascadeBuf I__4541 (
            .O(N__19142),
            .I(N__19139));
    CascadeMux I__4540 (
            .O(N__19139),
            .I(N__19136));
    CascadeBuf I__4539 (
            .O(N__19136),
            .I(N__19133));
    CascadeMux I__4538 (
            .O(N__19133),
            .I(N__19130));
    CascadeBuf I__4537 (
            .O(N__19130),
            .I(N__19127));
    CascadeMux I__4536 (
            .O(N__19127),
            .I(N__19124));
    CascadeBuf I__4535 (
            .O(N__19124),
            .I(N__19121));
    CascadeMux I__4534 (
            .O(N__19121),
            .I(N__19118));
    CascadeBuf I__4533 (
            .O(N__19118),
            .I(N__19115));
    CascadeMux I__4532 (
            .O(N__19115),
            .I(N__19112));
    InMux I__4531 (
            .O(N__19112),
            .I(N__19109));
    LocalMux I__4530 (
            .O(N__19109),
            .I(N__19106));
    Odrv4 I__4529 (
            .O(N__19106),
            .I(M_this_vga_signals_address_2));
    InMux I__4528 (
            .O(N__19103),
            .I(N__19100));
    LocalMux I__4527 (
            .O(N__19100),
            .I(N__19097));
    Odrv4 I__4526 (
            .O(N__19097),
            .I(\this_vram.mem_out_bus2_2 ));
    InMux I__4525 (
            .O(N__19094),
            .I(N__19091));
    LocalMux I__4524 (
            .O(N__19091),
            .I(N__19088));
    Span4Mux_h I__4523 (
            .O(N__19088),
            .I(N__19085));
    Sp12to4 I__4522 (
            .O(N__19085),
            .I(N__19082));
    Span12Mux_v I__4521 (
            .O(N__19082),
            .I(N__19079));
    Odrv12 I__4520 (
            .O(N__19079),
            .I(\this_vram.mem_out_bus6_2 ));
    CascadeMux I__4519 (
            .O(N__19076),
            .I(\this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_ ));
    InMux I__4518 (
            .O(N__19073),
            .I(N__19070));
    LocalMux I__4517 (
            .O(N__19070),
            .I(\this_vram.mem_mem_0_1_RNISOIZ0Z11 ));
    InMux I__4516 (
            .O(N__19067),
            .I(N__19063));
    InMux I__4515 (
            .O(N__19066),
            .I(N__19060));
    LocalMux I__4514 (
            .O(N__19063),
            .I(N__19055));
    LocalMux I__4513 (
            .O(N__19060),
            .I(N__19055));
    Span4Mux_v I__4512 (
            .O(N__19055),
            .I(N__19052));
    Span4Mux_h I__4511 (
            .O(N__19052),
            .I(N__19049));
    Odrv4 I__4510 (
            .O(N__19049),
            .I(\this_vram.mem_N_98 ));
    InMux I__4509 (
            .O(N__19046),
            .I(N__19043));
    LocalMux I__4508 (
            .O(N__19043),
            .I(N__19040));
    Sp12to4 I__4507 (
            .O(N__19040),
            .I(N__19037));
    Span12Mux_v I__4506 (
            .O(N__19037),
            .I(N__19034));
    Odrv12 I__4505 (
            .O(N__19034),
            .I(\this_vram.mem_out_bus1_3 ));
    InMux I__4504 (
            .O(N__19031),
            .I(N__19028));
    LocalMux I__4503 (
            .O(N__19028),
            .I(N__19025));
    Span4Mux_v I__4502 (
            .O(N__19025),
            .I(N__19022));
    Span4Mux_v I__4501 (
            .O(N__19022),
            .I(N__19019));
    Odrv4 I__4500 (
            .O(N__19019),
            .I(\this_vram.mem_out_bus5_3 ));
    CascadeMux I__4499 (
            .O(N__19016),
            .I(N__19013));
    InMux I__4498 (
            .O(N__19013),
            .I(N__19010));
    LocalMux I__4497 (
            .O(N__19010),
            .I(\this_vram.mem_out_bus3_3 ));
    InMux I__4496 (
            .O(N__19007),
            .I(N__19004));
    LocalMux I__4495 (
            .O(N__19004),
            .I(N__19001));
    Span4Mux_v I__4494 (
            .O(N__19001),
            .I(N__18998));
    Span4Mux_v I__4493 (
            .O(N__18998),
            .I(N__18995));
    Span4Mux_v I__4492 (
            .O(N__18995),
            .I(N__18992));
    Span4Mux_v I__4491 (
            .O(N__18992),
            .I(N__18989));
    Odrv4 I__4490 (
            .O(N__18989),
            .I(\this_vram.mem_out_bus7_3 ));
    CascadeMux I__4489 (
            .O(N__18986),
            .I(\this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_ ));
    InMux I__4488 (
            .O(N__18983),
            .I(N__18980));
    LocalMux I__4487 (
            .O(N__18980),
            .I(N__18977));
    Odrv4 I__4486 (
            .O(N__18977),
            .I(\this_vram.mem_mem_1_1_RNIUSK11Z0Z_0 ));
    InMux I__4485 (
            .O(N__18974),
            .I(N__18970));
    InMux I__4484 (
            .O(N__18973),
            .I(N__18967));
    LocalMux I__4483 (
            .O(N__18970),
            .I(N__18962));
    LocalMux I__4482 (
            .O(N__18967),
            .I(N__18962));
    Span4Mux_v I__4481 (
            .O(N__18962),
            .I(N__18959));
    Span4Mux_h I__4480 (
            .O(N__18959),
            .I(N__18956));
    Odrv4 I__4479 (
            .O(N__18956),
            .I(\this_vram.mem_N_102 ));
    InMux I__4478 (
            .O(N__18953),
            .I(N__18950));
    LocalMux I__4477 (
            .O(N__18950),
            .I(N__18947));
    Odrv4 I__4476 (
            .O(N__18947),
            .I(\this_vram.mem_mem_1_0_RNISSKZ0Z11 ));
    InMux I__4475 (
            .O(N__18944),
            .I(N__18940));
    InMux I__4474 (
            .O(N__18943),
            .I(N__18937));
    LocalMux I__4473 (
            .O(N__18940),
            .I(N__18931));
    LocalMux I__4472 (
            .O(N__18937),
            .I(N__18931));
    InMux I__4471 (
            .O(N__18936),
            .I(N__18928));
    Span4Mux_v I__4470 (
            .O(N__18931),
            .I(N__18925));
    LocalMux I__4469 (
            .O(N__18928),
            .I(N__18922));
    Span4Mux_h I__4468 (
            .O(N__18925),
            .I(N__18917));
    Span4Mux_v I__4467 (
            .O(N__18922),
            .I(N__18917));
    Span4Mux_h I__4466 (
            .O(N__18917),
            .I(N__18914));
    Odrv4 I__4465 (
            .O(N__18914),
            .I(this_vram_mem_N_109));
    InMux I__4464 (
            .O(N__18911),
            .I(N__18908));
    LocalMux I__4463 (
            .O(N__18908),
            .I(\this_vram.mem_out_bus3_2 ));
    InMux I__4462 (
            .O(N__18905),
            .I(N__18902));
    LocalMux I__4461 (
            .O(N__18902),
            .I(N__18899));
    Span4Mux_v I__4460 (
            .O(N__18899),
            .I(N__18896));
    Sp12to4 I__4459 (
            .O(N__18896),
            .I(N__18893));
    Span12Mux_v I__4458 (
            .O(N__18893),
            .I(N__18890));
    Odrv12 I__4457 (
            .O(N__18890),
            .I(\this_vram.mem_out_bus7_2 ));
    InMux I__4456 (
            .O(N__18887),
            .I(N__18884));
    LocalMux I__4455 (
            .O(N__18884),
            .I(\this_vram.mem_mem_1_1_RNIUSKZ0Z11 ));
    CascadeMux I__4454 (
            .O(N__18881),
            .I(\this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_ ));
    InMux I__4453 (
            .O(N__18878),
            .I(N__18873));
    InMux I__4452 (
            .O(N__18877),
            .I(N__18870));
    InMux I__4451 (
            .O(N__18876),
            .I(N__18867));
    LocalMux I__4450 (
            .O(N__18873),
            .I(N__18858));
    LocalMux I__4449 (
            .O(N__18870),
            .I(N__18858));
    LocalMux I__4448 (
            .O(N__18867),
            .I(N__18855));
    InMux I__4447 (
            .O(N__18866),
            .I(N__18852));
    InMux I__4446 (
            .O(N__18865),
            .I(N__18844));
    InMux I__4445 (
            .O(N__18864),
            .I(N__18844));
    InMux I__4444 (
            .O(N__18863),
            .I(N__18844));
    Span4Mux_v I__4443 (
            .O(N__18858),
            .I(N__18837));
    Span4Mux_h I__4442 (
            .O(N__18855),
            .I(N__18837));
    LocalMux I__4441 (
            .O(N__18852),
            .I(N__18837));
    InMux I__4440 (
            .O(N__18851),
            .I(N__18834));
    LocalMux I__4439 (
            .O(N__18844),
            .I(N__18827));
    Span4Mux_h I__4438 (
            .O(N__18837),
            .I(N__18827));
    LocalMux I__4437 (
            .O(N__18834),
            .I(N__18827));
    Span4Mux_v I__4436 (
            .O(N__18827),
            .I(N__18824));
    Odrv4 I__4435 (
            .O(N__18824),
            .I(\this_vram.mem_radregZ0Z_12 ));
    InMux I__4434 (
            .O(N__18821),
            .I(N__18815));
    InMux I__4433 (
            .O(N__18820),
            .I(N__18815));
    LocalMux I__4432 (
            .O(N__18815),
            .I(N__18812));
    Span4Mux_v I__4431 (
            .O(N__18812),
            .I(N__18809));
    Span4Mux_h I__4430 (
            .O(N__18809),
            .I(N__18806));
    Odrv4 I__4429 (
            .O(N__18806),
            .I(\this_vram.mem_N_95 ));
    InMux I__4428 (
            .O(N__18803),
            .I(N__18800));
    LocalMux I__4427 (
            .O(N__18800),
            .I(N__18797));
    Span4Mux_h I__4426 (
            .O(N__18797),
            .I(N__18794));
    Sp12to4 I__4425 (
            .O(N__18794),
            .I(N__18791));
    Odrv12 I__4424 (
            .O(N__18791),
            .I(\this_vram.mem_out_bus6_0 ));
    InMux I__4423 (
            .O(N__18788),
            .I(N__18785));
    LocalMux I__4422 (
            .O(N__18785),
            .I(N__18782));
    Span4Mux_v I__4421 (
            .O(N__18782),
            .I(N__18779));
    Odrv4 I__4420 (
            .O(N__18779),
            .I(\this_vram.mem_out_bus2_0 ));
    InMux I__4419 (
            .O(N__18776),
            .I(N__18773));
    LocalMux I__4418 (
            .O(N__18773),
            .I(N__18770));
    Span4Mux_v I__4417 (
            .O(N__18770),
            .I(N__18767));
    Odrv4 I__4416 (
            .O(N__18767),
            .I(\this_vram.mem_out_bus2_1 ));
    InMux I__4415 (
            .O(N__18764),
            .I(N__18761));
    LocalMux I__4414 (
            .O(N__18761),
            .I(N__18758));
    Span4Mux_v I__4413 (
            .O(N__18758),
            .I(N__18755));
    Span4Mux_v I__4412 (
            .O(N__18755),
            .I(N__18752));
    Span4Mux_v I__4411 (
            .O(N__18752),
            .I(N__18749));
    Odrv4 I__4410 (
            .O(N__18749),
            .I(\this_vram.mem_out_bus6_1 ));
    InMux I__4409 (
            .O(N__18746),
            .I(N__18743));
    LocalMux I__4408 (
            .O(N__18743),
            .I(\this_vram.mem_mem_0_0_RNIQOI11Z0Z_0 ));
    CascadeMux I__4407 (
            .O(N__18740),
            .I(\this_vram.mem_mem_2_0_RNIU0N11Z0Z_0_cascade_ ));
    InMux I__4406 (
            .O(N__18737),
            .I(N__18733));
    InMux I__4405 (
            .O(N__18736),
            .I(N__18730));
    LocalMux I__4404 (
            .O(N__18733),
            .I(N__18727));
    LocalMux I__4403 (
            .O(N__18730),
            .I(N__18724));
    Span4Mux_v I__4402 (
            .O(N__18727),
            .I(N__18721));
    Span4Mux_v I__4401 (
            .O(N__18724),
            .I(N__18718));
    Span4Mux_h I__4400 (
            .O(N__18721),
            .I(N__18715));
    Span4Mux_h I__4399 (
            .O(N__18718),
            .I(N__18712));
    Odrv4 I__4398 (
            .O(N__18715),
            .I(\this_vram.mem_N_91 ));
    Odrv4 I__4397 (
            .O(N__18712),
            .I(\this_vram.mem_N_91 ));
    InMux I__4396 (
            .O(N__18707),
            .I(N__18704));
    LocalMux I__4395 (
            .O(N__18704),
            .I(N__18701));
    Sp12to4 I__4394 (
            .O(N__18701),
            .I(N__18698));
    Odrv12 I__4393 (
            .O(N__18698),
            .I(\this_vram.mem_out_bus5_1 ));
    InMux I__4392 (
            .O(N__18695),
            .I(N__18692));
    LocalMux I__4391 (
            .O(N__18692),
            .I(N__18689));
    Sp12to4 I__4390 (
            .O(N__18689),
            .I(N__18686));
    Span12Mux_v I__4389 (
            .O(N__18686),
            .I(N__18683));
    Odrv12 I__4388 (
            .O(N__18683),
            .I(\this_vram.mem_out_bus1_1 ));
    InMux I__4387 (
            .O(N__18680),
            .I(N__18677));
    LocalMux I__4386 (
            .O(N__18677),
            .I(\this_vram.mem_mem_1_0_RNISSK11Z0Z_0 ));
    InMux I__4385 (
            .O(N__18674),
            .I(N__18671));
    LocalMux I__4384 (
            .O(N__18671),
            .I(\this_vram.mem_out_bus3_1 ));
    InMux I__4383 (
            .O(N__18668),
            .I(N__18665));
    LocalMux I__4382 (
            .O(N__18665),
            .I(N__18662));
    Sp12to4 I__4381 (
            .O(N__18662),
            .I(N__18659));
    Span12Mux_v I__4380 (
            .O(N__18659),
            .I(N__18656));
    Odrv12 I__4379 (
            .O(N__18656),
            .I(\this_vram.mem_out_bus7_1 ));
    InMux I__4378 (
            .O(N__18653),
            .I(N__18650));
    LocalMux I__4377 (
            .O(N__18650),
            .I(\this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ));
    InMux I__4376 (
            .O(N__18647),
            .I(N__18644));
    LocalMux I__4375 (
            .O(N__18644),
            .I(N__18641));
    Span4Mux_v I__4374 (
            .O(N__18641),
            .I(N__18638));
    Odrv4 I__4373 (
            .O(N__18638),
            .I(\this_vram.mem_out_bus1_0 ));
    InMux I__4372 (
            .O(N__18635),
            .I(N__18632));
    LocalMux I__4371 (
            .O(N__18632),
            .I(N__18629));
    Span4Mux_v I__4370 (
            .O(N__18629),
            .I(N__18626));
    Span4Mux_v I__4369 (
            .O(N__18626),
            .I(N__18623));
    Odrv4 I__4368 (
            .O(N__18623),
            .I(\this_vram.mem_out_bus5_0 ));
    InMux I__4367 (
            .O(N__18620),
            .I(N__18617));
    LocalMux I__4366 (
            .O(N__18617),
            .I(N__18614));
    Odrv4 I__4365 (
            .O(N__18614),
            .I(\this_vram.mem_out_bus2_3 ));
    InMux I__4364 (
            .O(N__18611),
            .I(N__18608));
    LocalMux I__4363 (
            .O(N__18608),
            .I(N__18605));
    Span4Mux_h I__4362 (
            .O(N__18605),
            .I(N__18602));
    Sp12to4 I__4361 (
            .O(N__18602),
            .I(N__18599));
    Span12Mux_v I__4360 (
            .O(N__18599),
            .I(N__18596));
    Odrv12 I__4359 (
            .O(N__18596),
            .I(\this_vram.mem_out_bus6_3 ));
    InMux I__4358 (
            .O(N__18593),
            .I(N__18590));
    LocalMux I__4357 (
            .O(N__18590),
            .I(\this_vram.mem_mem_2_1_RNI01N11Z0Z_0 ));
    InMux I__4356 (
            .O(N__18587),
            .I(N__18584));
    LocalMux I__4355 (
            .O(N__18584),
            .I(N__18581));
    Span4Mux_v I__4354 (
            .O(N__18581),
            .I(N__18578));
    Span4Mux_v I__4353 (
            .O(N__18578),
            .I(N__18575));
    Odrv4 I__4352 (
            .O(N__18575),
            .I(\this_vram.mem_out_bus0_2 ));
    InMux I__4351 (
            .O(N__18572),
            .I(N__18569));
    LocalMux I__4350 (
            .O(N__18569),
            .I(N__18566));
    Span4Mux_v I__4349 (
            .O(N__18566),
            .I(N__18563));
    Odrv4 I__4348 (
            .O(N__18563),
            .I(\this_vram.mem_out_bus4_2 ));
    InMux I__4347 (
            .O(N__18560),
            .I(N__18557));
    LocalMux I__4346 (
            .O(N__18557),
            .I(N__18554));
    Span4Mux_v I__4345 (
            .O(N__18554),
            .I(N__18551));
    Odrv4 I__4344 (
            .O(N__18551),
            .I(\this_vram.mem_out_bus1_2 ));
    InMux I__4343 (
            .O(N__18548),
            .I(N__18545));
    LocalMux I__4342 (
            .O(N__18545),
            .I(N__18542));
    Span4Mux_v I__4341 (
            .O(N__18542),
            .I(N__18539));
    Span4Mux_v I__4340 (
            .O(N__18539),
            .I(N__18536));
    Odrv4 I__4339 (
            .O(N__18536),
            .I(\this_vram.mem_out_bus5_2 ));
    InMux I__4338 (
            .O(N__18533),
            .I(N__18530));
    LocalMux I__4337 (
            .O(N__18530),
            .I(N__18527));
    Span4Mux_v I__4336 (
            .O(N__18527),
            .I(N__18524));
    Span4Mux_v I__4335 (
            .O(N__18524),
            .I(N__18521));
    Odrv4 I__4334 (
            .O(N__18521),
            .I(\this_vram.mem_out_bus4_3 ));
    CascadeMux I__4333 (
            .O(N__18518),
            .I(N__18515));
    InMux I__4332 (
            .O(N__18515),
            .I(N__18511));
    InMux I__4331 (
            .O(N__18514),
            .I(N__18508));
    LocalMux I__4330 (
            .O(N__18511),
            .I(N__18503));
    LocalMux I__4329 (
            .O(N__18508),
            .I(N__18503));
    Span4Mux_v I__4328 (
            .O(N__18503),
            .I(N__18500));
    Span4Mux_h I__4327 (
            .O(N__18500),
            .I(N__18497));
    Odrv4 I__4326 (
            .O(N__18497),
            .I(\this_vram.mem_N_88 ));
    InMux I__4325 (
            .O(N__18494),
            .I(N__18491));
    LocalMux I__4324 (
            .O(N__18491),
            .I(N__18488));
    Odrv4 I__4323 (
            .O(N__18488),
            .I(\this_vram.mem_mem_0_1_RNISOI11Z0Z_0 ));
    InMux I__4322 (
            .O(N__18485),
            .I(N__18481));
    InMux I__4321 (
            .O(N__18484),
            .I(N__18478));
    LocalMux I__4320 (
            .O(N__18481),
            .I(N__18473));
    LocalMux I__4319 (
            .O(N__18478),
            .I(N__18473));
    Span4Mux_v I__4318 (
            .O(N__18473),
            .I(N__18470));
    Span4Mux_h I__4317 (
            .O(N__18470),
            .I(N__18467));
    Odrv4 I__4316 (
            .O(N__18467),
            .I(\this_vram.mem_N_105 ));
    CEMux I__4315 (
            .O(N__18464),
            .I(N__18461));
    LocalMux I__4314 (
            .O(N__18461),
            .I(N__18457));
    CEMux I__4313 (
            .O(N__18460),
            .I(N__18454));
    Span4Mux_h I__4312 (
            .O(N__18457),
            .I(N__18451));
    LocalMux I__4311 (
            .O(N__18454),
            .I(N__18448));
    Span4Mux_v I__4310 (
            .O(N__18451),
            .I(N__18445));
    Span4Mux_h I__4309 (
            .O(N__18448),
            .I(N__18442));
    Odrv4 I__4308 (
            .O(N__18445),
            .I(\this_vram.mem_WE_10 ));
    Odrv4 I__4307 (
            .O(N__18442),
            .I(\this_vram.mem_WE_10 ));
    CEMux I__4306 (
            .O(N__18437),
            .I(N__18433));
    CEMux I__4305 (
            .O(N__18436),
            .I(N__18430));
    LocalMux I__4304 (
            .O(N__18433),
            .I(N__18427));
    LocalMux I__4303 (
            .O(N__18430),
            .I(N__18424));
    Span4Mux_h I__4302 (
            .O(N__18427),
            .I(N__18421));
    Span12Mux_s2_v I__4301 (
            .O(N__18424),
            .I(N__18418));
    Span4Mux_v I__4300 (
            .O(N__18421),
            .I(N__18415));
    Span12Mux_v I__4299 (
            .O(N__18418),
            .I(N__18412));
    Span4Mux_v I__4298 (
            .O(N__18415),
            .I(N__18409));
    Odrv12 I__4297 (
            .O(N__18412),
            .I(\this_vram.mem_WE_14 ));
    Odrv4 I__4296 (
            .O(N__18409),
            .I(\this_vram.mem_WE_14 ));
    InMux I__4295 (
            .O(N__18404),
            .I(N__18401));
    LocalMux I__4294 (
            .O(N__18401),
            .I(N__18398));
    Span4Mux_v I__4293 (
            .O(N__18398),
            .I(N__18393));
    InMux I__4292 (
            .O(N__18397),
            .I(N__18390));
    InMux I__4291 (
            .O(N__18396),
            .I(N__18387));
    Sp12to4 I__4290 (
            .O(N__18393),
            .I(N__18382));
    LocalMux I__4289 (
            .O(N__18390),
            .I(N__18382));
    LocalMux I__4288 (
            .O(N__18387),
            .I(N__18379));
    Span12Mux_h I__4287 (
            .O(N__18382),
            .I(N__18374));
    Span12Mux_v I__4286 (
            .O(N__18379),
            .I(N__18374));
    Odrv12 I__4285 (
            .O(N__18374),
            .I(this_vram_mem_N_112));
    InMux I__4284 (
            .O(N__18371),
            .I(N__18367));
    InMux I__4283 (
            .O(N__18370),
            .I(N__18364));
    LocalMux I__4282 (
            .O(N__18367),
            .I(N__18360));
    LocalMux I__4281 (
            .O(N__18364),
            .I(N__18355));
    InMux I__4280 (
            .O(N__18363),
            .I(N__18352));
    Span4Mux_v I__4279 (
            .O(N__18360),
            .I(N__18349));
    InMux I__4278 (
            .O(N__18359),
            .I(N__18346));
    InMux I__4277 (
            .O(N__18358),
            .I(N__18343));
    Span4Mux_v I__4276 (
            .O(N__18355),
            .I(N__18332));
    LocalMux I__4275 (
            .O(N__18352),
            .I(N__18329));
    Sp12to4 I__4274 (
            .O(N__18349),
            .I(N__18326));
    LocalMux I__4273 (
            .O(N__18346),
            .I(N__18323));
    LocalMux I__4272 (
            .O(N__18343),
            .I(N__18319));
    InMux I__4271 (
            .O(N__18342),
            .I(N__18316));
    InMux I__4270 (
            .O(N__18341),
            .I(N__18309));
    InMux I__4269 (
            .O(N__18340),
            .I(N__18309));
    InMux I__4268 (
            .O(N__18339),
            .I(N__18309));
    InMux I__4267 (
            .O(N__18338),
            .I(N__18304));
    InMux I__4266 (
            .O(N__18337),
            .I(N__18304));
    InMux I__4265 (
            .O(N__18336),
            .I(N__18298));
    InMux I__4264 (
            .O(N__18335),
            .I(N__18298));
    Sp12to4 I__4263 (
            .O(N__18332),
            .I(N__18291));
    Span12Mux_v I__4262 (
            .O(N__18329),
            .I(N__18291));
    Span12Mux_h I__4261 (
            .O(N__18326),
            .I(N__18288));
    Span4Mux_h I__4260 (
            .O(N__18323),
            .I(N__18285));
    InMux I__4259 (
            .O(N__18322),
            .I(N__18282));
    Span4Mux_h I__4258 (
            .O(N__18319),
            .I(N__18275));
    LocalMux I__4257 (
            .O(N__18316),
            .I(N__18275));
    LocalMux I__4256 (
            .O(N__18309),
            .I(N__18275));
    LocalMux I__4255 (
            .O(N__18304),
            .I(N__18272));
    InMux I__4254 (
            .O(N__18303),
            .I(N__18269));
    LocalMux I__4253 (
            .O(N__18298),
            .I(N__18266));
    InMux I__4252 (
            .O(N__18297),
            .I(N__18263));
    InMux I__4251 (
            .O(N__18296),
            .I(N__18260));
    Odrv12 I__4250 (
            .O(N__18291),
            .I(\this_vga_signals.rgb_1_4 ));
    Odrv12 I__4249 (
            .O(N__18288),
            .I(\this_vga_signals.rgb_1_4 ));
    Odrv4 I__4248 (
            .O(N__18285),
            .I(\this_vga_signals.rgb_1_4 ));
    LocalMux I__4247 (
            .O(N__18282),
            .I(\this_vga_signals.rgb_1_4 ));
    Odrv4 I__4246 (
            .O(N__18275),
            .I(\this_vga_signals.rgb_1_4 ));
    Odrv4 I__4245 (
            .O(N__18272),
            .I(\this_vga_signals.rgb_1_4 ));
    LocalMux I__4244 (
            .O(N__18269),
            .I(\this_vga_signals.rgb_1_4 ));
    Odrv4 I__4243 (
            .O(N__18266),
            .I(\this_vga_signals.rgb_1_4 ));
    LocalMux I__4242 (
            .O(N__18263),
            .I(\this_vga_signals.rgb_1_4 ));
    LocalMux I__4241 (
            .O(N__18260),
            .I(\this_vga_signals.rgb_1_4 ));
    ClkMux I__4240 (
            .O(N__18239),
            .I(N__18056));
    ClkMux I__4239 (
            .O(N__18238),
            .I(N__18056));
    ClkMux I__4238 (
            .O(N__18237),
            .I(N__18056));
    ClkMux I__4237 (
            .O(N__18236),
            .I(N__18056));
    ClkMux I__4236 (
            .O(N__18235),
            .I(N__18056));
    ClkMux I__4235 (
            .O(N__18234),
            .I(N__18056));
    ClkMux I__4234 (
            .O(N__18233),
            .I(N__18056));
    ClkMux I__4233 (
            .O(N__18232),
            .I(N__18056));
    ClkMux I__4232 (
            .O(N__18231),
            .I(N__18056));
    ClkMux I__4231 (
            .O(N__18230),
            .I(N__18056));
    ClkMux I__4230 (
            .O(N__18229),
            .I(N__18056));
    ClkMux I__4229 (
            .O(N__18228),
            .I(N__18056));
    ClkMux I__4228 (
            .O(N__18227),
            .I(N__18056));
    ClkMux I__4227 (
            .O(N__18226),
            .I(N__18056));
    ClkMux I__4226 (
            .O(N__18225),
            .I(N__18056));
    ClkMux I__4225 (
            .O(N__18224),
            .I(N__18056));
    ClkMux I__4224 (
            .O(N__18223),
            .I(N__18056));
    ClkMux I__4223 (
            .O(N__18222),
            .I(N__18056));
    ClkMux I__4222 (
            .O(N__18221),
            .I(N__18056));
    ClkMux I__4221 (
            .O(N__18220),
            .I(N__18056));
    ClkMux I__4220 (
            .O(N__18219),
            .I(N__18056));
    ClkMux I__4219 (
            .O(N__18218),
            .I(N__18056));
    ClkMux I__4218 (
            .O(N__18217),
            .I(N__18056));
    ClkMux I__4217 (
            .O(N__18216),
            .I(N__18056));
    ClkMux I__4216 (
            .O(N__18215),
            .I(N__18056));
    ClkMux I__4215 (
            .O(N__18214),
            .I(N__18056));
    ClkMux I__4214 (
            .O(N__18213),
            .I(N__18056));
    ClkMux I__4213 (
            .O(N__18212),
            .I(N__18056));
    ClkMux I__4212 (
            .O(N__18211),
            .I(N__18056));
    ClkMux I__4211 (
            .O(N__18210),
            .I(N__18056));
    ClkMux I__4210 (
            .O(N__18209),
            .I(N__18056));
    ClkMux I__4209 (
            .O(N__18208),
            .I(N__18056));
    ClkMux I__4208 (
            .O(N__18207),
            .I(N__18056));
    ClkMux I__4207 (
            .O(N__18206),
            .I(N__18056));
    ClkMux I__4206 (
            .O(N__18205),
            .I(N__18056));
    ClkMux I__4205 (
            .O(N__18204),
            .I(N__18056));
    ClkMux I__4204 (
            .O(N__18203),
            .I(N__18056));
    ClkMux I__4203 (
            .O(N__18202),
            .I(N__18056));
    ClkMux I__4202 (
            .O(N__18201),
            .I(N__18056));
    ClkMux I__4201 (
            .O(N__18200),
            .I(N__18056));
    ClkMux I__4200 (
            .O(N__18199),
            .I(N__18056));
    ClkMux I__4199 (
            .O(N__18198),
            .I(N__18056));
    ClkMux I__4198 (
            .O(N__18197),
            .I(N__18056));
    ClkMux I__4197 (
            .O(N__18196),
            .I(N__18056));
    ClkMux I__4196 (
            .O(N__18195),
            .I(N__18056));
    ClkMux I__4195 (
            .O(N__18194),
            .I(N__18056));
    ClkMux I__4194 (
            .O(N__18193),
            .I(N__18056));
    ClkMux I__4193 (
            .O(N__18192),
            .I(N__18056));
    ClkMux I__4192 (
            .O(N__18191),
            .I(N__18056));
    ClkMux I__4191 (
            .O(N__18190),
            .I(N__18056));
    ClkMux I__4190 (
            .O(N__18189),
            .I(N__18056));
    ClkMux I__4189 (
            .O(N__18188),
            .I(N__18056));
    ClkMux I__4188 (
            .O(N__18187),
            .I(N__18056));
    ClkMux I__4187 (
            .O(N__18186),
            .I(N__18056));
    ClkMux I__4186 (
            .O(N__18185),
            .I(N__18056));
    ClkMux I__4185 (
            .O(N__18184),
            .I(N__18056));
    ClkMux I__4184 (
            .O(N__18183),
            .I(N__18056));
    ClkMux I__4183 (
            .O(N__18182),
            .I(N__18056));
    ClkMux I__4182 (
            .O(N__18181),
            .I(N__18056));
    ClkMux I__4181 (
            .O(N__18180),
            .I(N__18056));
    ClkMux I__4180 (
            .O(N__18179),
            .I(N__18056));
    GlobalMux I__4179 (
            .O(N__18056),
            .I(N__18053));
    gio2CtrlBuf I__4178 (
            .O(N__18053),
            .I(clk_0_c_g));
    CascadeMux I__4177 (
            .O(N__18050),
            .I(N__18046));
    InMux I__4176 (
            .O(N__18049),
            .I(N__18040));
    InMux I__4175 (
            .O(N__18046),
            .I(N__18040));
    InMux I__4174 (
            .O(N__18045),
            .I(N__18037));
    LocalMux I__4173 (
            .O(N__18040),
            .I(N__18034));
    LocalMux I__4172 (
            .O(N__18037),
            .I(N__18031));
    Sp12to4 I__4171 (
            .O(N__18034),
            .I(N__18028));
    Span4Mux_v I__4170 (
            .O(N__18031),
            .I(N__18025));
    Span12Mux_v I__4169 (
            .O(N__18028),
            .I(N__18022));
    Sp12to4 I__4168 (
            .O(N__18025),
            .I(N__18019));
    Span12Mux_h I__4167 (
            .O(N__18022),
            .I(N__18016));
    Span12Mux_h I__4166 (
            .O(N__18019),
            .I(N__18013));
    Odrv12 I__4165 (
            .O(N__18016),
            .I(port_data_c_3));
    Odrv12 I__4164 (
            .O(N__18013),
            .I(port_data_c_3));
    InMux I__4163 (
            .O(N__18008),
            .I(N__18005));
    LocalMux I__4162 (
            .O(N__18005),
            .I(N__18000));
    InMux I__4161 (
            .O(N__18004),
            .I(N__17997));
    InMux I__4160 (
            .O(N__18003),
            .I(N__17993));
    Span4Mux_h I__4159 (
            .O(N__18000),
            .I(N__17989));
    LocalMux I__4158 (
            .O(N__17997),
            .I(N__17986));
    InMux I__4157 (
            .O(N__17996),
            .I(N__17983));
    LocalMux I__4156 (
            .O(N__17993),
            .I(N__17979));
    InMux I__4155 (
            .O(N__17992),
            .I(N__17976));
    Span4Mux_v I__4154 (
            .O(N__17989),
            .I(N__17971));
    Span4Mux_h I__4153 (
            .O(N__17986),
            .I(N__17971));
    LocalMux I__4152 (
            .O(N__17983),
            .I(N__17968));
    InMux I__4151 (
            .O(N__17982),
            .I(N__17965));
    Span4Mux_h I__4150 (
            .O(N__17979),
            .I(N__17960));
    LocalMux I__4149 (
            .O(N__17976),
            .I(N__17957));
    Span4Mux_v I__4148 (
            .O(N__17971),
            .I(N__17952));
    Span4Mux_h I__4147 (
            .O(N__17968),
            .I(N__17952));
    LocalMux I__4146 (
            .O(N__17965),
            .I(N__17949));
    InMux I__4145 (
            .O(N__17964),
            .I(N__17946));
    InMux I__4144 (
            .O(N__17963),
            .I(N__17943));
    Span4Mux_v I__4143 (
            .O(N__17960),
            .I(N__17938));
    Span4Mux_h I__4142 (
            .O(N__17957),
            .I(N__17938));
    Span4Mux_v I__4141 (
            .O(N__17952),
            .I(N__17933));
    Span4Mux_h I__4140 (
            .O(N__17949),
            .I(N__17933));
    LocalMux I__4139 (
            .O(N__17946),
            .I(N__17930));
    LocalMux I__4138 (
            .O(N__17943),
            .I(N__17927));
    Span4Mux_v I__4137 (
            .O(N__17938),
            .I(N__17918));
    Span4Mux_v I__4136 (
            .O(N__17933),
            .I(N__17918));
    Span4Mux_h I__4135 (
            .O(N__17930),
            .I(N__17918));
    Span4Mux_h I__4134 (
            .O(N__17927),
            .I(N__17918));
    Odrv4 I__4133 (
            .O(N__17918),
            .I(M_this_vram_write_data_3));
    InMux I__4132 (
            .O(N__17915),
            .I(N__17912));
    LocalMux I__4131 (
            .O(N__17912),
            .I(N__17909));
    Span4Mux_v I__4130 (
            .O(N__17909),
            .I(N__17906));
    Odrv4 I__4129 (
            .O(N__17906),
            .I(\this_vram.mem_out_bus4_1 ));
    InMux I__4128 (
            .O(N__17903),
            .I(N__17900));
    LocalMux I__4127 (
            .O(N__17900),
            .I(N__17897));
    Span4Mux_v I__4126 (
            .O(N__17897),
            .I(N__17894));
    Span4Mux_v I__4125 (
            .O(N__17894),
            .I(N__17891));
    Odrv4 I__4124 (
            .O(N__17891),
            .I(\this_vram.mem_out_bus0_1 ));
    CascadeMux I__4123 (
            .O(N__17888),
            .I(rgbZ0Z_1_cascade_));
    InMux I__4122 (
            .O(N__17885),
            .I(N__17882));
    LocalMux I__4121 (
            .O(N__17882),
            .I(M_vcounter_q_esr_RNI2RH6LA_9));
    InMux I__4120 (
            .O(N__17879),
            .I(N__17875));
    CascadeMux I__4119 (
            .O(N__17878),
            .I(N__17870));
    LocalMux I__4118 (
            .O(N__17875),
            .I(N__17866));
    InMux I__4117 (
            .O(N__17874),
            .I(N__17862));
    InMux I__4116 (
            .O(N__17873),
            .I(N__17859));
    InMux I__4115 (
            .O(N__17870),
            .I(N__17854));
    InMux I__4114 (
            .O(N__17869),
            .I(N__17854));
    Span4Mux_v I__4113 (
            .O(N__17866),
            .I(N__17850));
    CascadeMux I__4112 (
            .O(N__17865),
            .I(N__17847));
    LocalMux I__4111 (
            .O(N__17862),
            .I(N__17843));
    LocalMux I__4110 (
            .O(N__17859),
            .I(N__17840));
    LocalMux I__4109 (
            .O(N__17854),
            .I(N__17837));
    CascadeMux I__4108 (
            .O(N__17853),
            .I(N__17834));
    Span4Mux_h I__4107 (
            .O(N__17850),
            .I(N__17828));
    InMux I__4106 (
            .O(N__17847),
            .I(N__17823));
    InMux I__4105 (
            .O(N__17846),
            .I(N__17823));
    Span4Mux_v I__4104 (
            .O(N__17843),
            .I(N__17816));
    Span4Mux_v I__4103 (
            .O(N__17840),
            .I(N__17816));
    Span4Mux_h I__4102 (
            .O(N__17837),
            .I(N__17816));
    InMux I__4101 (
            .O(N__17834),
            .I(N__17809));
    InMux I__4100 (
            .O(N__17833),
            .I(N__17809));
    InMux I__4099 (
            .O(N__17832),
            .I(N__17809));
    InMux I__4098 (
            .O(N__17831),
            .I(N__17806));
    Odrv4 I__4097 (
            .O(N__17828),
            .I(rgbZ0Z_1));
    LocalMux I__4096 (
            .O(N__17823),
            .I(rgbZ0Z_1));
    Odrv4 I__4095 (
            .O(N__17816),
            .I(rgbZ0Z_1));
    LocalMux I__4094 (
            .O(N__17809),
            .I(rgbZ0Z_1));
    LocalMux I__4093 (
            .O(N__17806),
            .I(rgbZ0Z_1));
    CascadeMux I__4092 (
            .O(N__17795),
            .I(N__17792));
    InMux I__4091 (
            .O(N__17792),
            .I(N__17789));
    LocalMux I__4090 (
            .O(N__17789),
            .I(N__17786));
    Odrv12 I__4089 (
            .O(N__17786),
            .I(M_vcounter_q_esr_RNIVLNKSA_9));
    InMux I__4088 (
            .O(N__17783),
            .I(N__17780));
    LocalMux I__4087 (
            .O(N__17780),
            .I(N__17776));
    CascadeMux I__4086 (
            .O(N__17779),
            .I(N__17771));
    Span4Mux_h I__4085 (
            .O(N__17776),
            .I(N__17766));
    InMux I__4084 (
            .O(N__17775),
            .I(N__17763));
    InMux I__4083 (
            .O(N__17774),
            .I(N__17754));
    InMux I__4082 (
            .O(N__17771),
            .I(N__17754));
    InMux I__4081 (
            .O(N__17770),
            .I(N__17754));
    InMux I__4080 (
            .O(N__17769),
            .I(N__17754));
    Odrv4 I__4079 (
            .O(N__17766),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__4078 (
            .O(N__17763),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__4077 (
            .O(N__17754),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    CascadeMux I__4076 (
            .O(N__17747),
            .I(N__17744));
    CascadeBuf I__4075 (
            .O(N__17744),
            .I(N__17741));
    CascadeMux I__4074 (
            .O(N__17741),
            .I(N__17738));
    CascadeBuf I__4073 (
            .O(N__17738),
            .I(N__17735));
    CascadeMux I__4072 (
            .O(N__17735),
            .I(N__17732));
    CascadeBuf I__4071 (
            .O(N__17732),
            .I(N__17729));
    CascadeMux I__4070 (
            .O(N__17729),
            .I(N__17726));
    CascadeBuf I__4069 (
            .O(N__17726),
            .I(N__17723));
    CascadeMux I__4068 (
            .O(N__17723),
            .I(N__17720));
    CascadeBuf I__4067 (
            .O(N__17720),
            .I(N__17717));
    CascadeMux I__4066 (
            .O(N__17717),
            .I(N__17714));
    CascadeBuf I__4065 (
            .O(N__17714),
            .I(N__17711));
    CascadeMux I__4064 (
            .O(N__17711),
            .I(N__17708));
    CascadeBuf I__4063 (
            .O(N__17708),
            .I(N__17705));
    CascadeMux I__4062 (
            .O(N__17705),
            .I(N__17702));
    CascadeBuf I__4061 (
            .O(N__17702),
            .I(N__17699));
    CascadeMux I__4060 (
            .O(N__17699),
            .I(N__17696));
    CascadeBuf I__4059 (
            .O(N__17696),
            .I(N__17693));
    CascadeMux I__4058 (
            .O(N__17693),
            .I(N__17690));
    CascadeBuf I__4057 (
            .O(N__17690),
            .I(N__17687));
    CascadeMux I__4056 (
            .O(N__17687),
            .I(N__17684));
    CascadeBuf I__4055 (
            .O(N__17684),
            .I(N__17681));
    CascadeMux I__4054 (
            .O(N__17681),
            .I(N__17678));
    CascadeBuf I__4053 (
            .O(N__17678),
            .I(N__17675));
    CascadeMux I__4052 (
            .O(N__17675),
            .I(N__17672));
    CascadeBuf I__4051 (
            .O(N__17672),
            .I(N__17669));
    CascadeMux I__4050 (
            .O(N__17669),
            .I(N__17666));
    CascadeBuf I__4049 (
            .O(N__17666),
            .I(N__17663));
    CascadeMux I__4048 (
            .O(N__17663),
            .I(N__17660));
    CascadeBuf I__4047 (
            .O(N__17660),
            .I(N__17657));
    CascadeMux I__4046 (
            .O(N__17657),
            .I(N__17654));
    InMux I__4045 (
            .O(N__17654),
            .I(N__17651));
    LocalMux I__4044 (
            .O(N__17651),
            .I(N__17648));
    Span4Mux_h I__4043 (
            .O(N__17648),
            .I(N__17644));
    InMux I__4042 (
            .O(N__17647),
            .I(N__17641));
    Span4Mux_v I__4041 (
            .O(N__17644),
            .I(N__17638));
    LocalMux I__4040 (
            .O(N__17641),
            .I(N__17635));
    Span4Mux_v I__4039 (
            .O(N__17638),
            .I(N__17632));
    Odrv4 I__4038 (
            .O(N__17635),
            .I(M_this_vga_signals_address_3));
    Odrv4 I__4037 (
            .O(N__17632),
            .I(M_this_vga_signals_address_3));
    InMux I__4036 (
            .O(N__17627),
            .I(N__17624));
    LocalMux I__4035 (
            .O(N__17624),
            .I(N__17619));
    InMux I__4034 (
            .O(N__17623),
            .I(N__17616));
    CascadeMux I__4033 (
            .O(N__17622),
            .I(N__17613));
    Span4Mux_v I__4032 (
            .O(N__17619),
            .I(N__17610));
    LocalMux I__4031 (
            .O(N__17616),
            .I(N__17607));
    InMux I__4030 (
            .O(N__17613),
            .I(N__17604));
    Sp12to4 I__4029 (
            .O(N__17610),
            .I(N__17601));
    Span4Mux_h I__4028 (
            .O(N__17607),
            .I(N__17598));
    LocalMux I__4027 (
            .O(N__17604),
            .I(N__17595));
    Span12Mux_h I__4026 (
            .O(N__17601),
            .I(N__17590));
    Sp12to4 I__4025 (
            .O(N__17598),
            .I(N__17590));
    Span12Mux_v I__4024 (
            .O(N__17595),
            .I(N__17587));
    Odrv12 I__4023 (
            .O(N__17590),
            .I(port_data_c_0));
    Odrv12 I__4022 (
            .O(N__17587),
            .I(port_data_c_0));
    InMux I__4021 (
            .O(N__17582),
            .I(N__17578));
    InMux I__4020 (
            .O(N__17581),
            .I(N__17574));
    LocalMux I__4019 (
            .O(N__17578),
            .I(N__17569));
    InMux I__4018 (
            .O(N__17577),
            .I(N__17566));
    LocalMux I__4017 (
            .O(N__17574),
            .I(N__17562));
    InMux I__4016 (
            .O(N__17573),
            .I(N__17559));
    InMux I__4015 (
            .O(N__17572),
            .I(N__17556));
    Span4Mux_s3_v I__4014 (
            .O(N__17569),
            .I(N__17550));
    LocalMux I__4013 (
            .O(N__17566),
            .I(N__17550));
    InMux I__4012 (
            .O(N__17565),
            .I(N__17547));
    Span4Mux_h I__4011 (
            .O(N__17562),
            .I(N__17544));
    LocalMux I__4010 (
            .O(N__17559),
            .I(N__17541));
    LocalMux I__4009 (
            .O(N__17556),
            .I(N__17538));
    InMux I__4008 (
            .O(N__17555),
            .I(N__17535));
    Span4Mux_v I__4007 (
            .O(N__17550),
            .I(N__17530));
    LocalMux I__4006 (
            .O(N__17547),
            .I(N__17530));
    Span4Mux_v I__4005 (
            .O(N__17544),
            .I(N__17525));
    Span4Mux_h I__4004 (
            .O(N__17541),
            .I(N__17525));
    Span4Mux_v I__4003 (
            .O(N__17538),
            .I(N__17520));
    LocalMux I__4002 (
            .O(N__17535),
            .I(N__17520));
    Sp12to4 I__4001 (
            .O(N__17530),
            .I(N__17516));
    Span4Mux_v I__4000 (
            .O(N__17525),
            .I(N__17511));
    Span4Mux_v I__3999 (
            .O(N__17520),
            .I(N__17511));
    InMux I__3998 (
            .O(N__17519),
            .I(N__17508));
    Span12Mux_v I__3997 (
            .O(N__17516),
            .I(N__17501));
    Sp12to4 I__3996 (
            .O(N__17511),
            .I(N__17501));
    LocalMux I__3995 (
            .O(N__17508),
            .I(N__17501));
    Odrv12 I__3994 (
            .O(N__17501),
            .I(M_this_vram_write_data_0));
    InMux I__3993 (
            .O(N__17498),
            .I(N__17495));
    LocalMux I__3992 (
            .O(N__17495),
            .I(N__17492));
    Span4Mux_h I__3991 (
            .O(N__17492),
            .I(N__17489));
    Span4Mux_h I__3990 (
            .O(N__17489),
            .I(N__17486));
    Odrv4 I__3989 (
            .O(N__17486),
            .I(\this_vga_signals.SUM_3_1 ));
    CascadeMux I__3988 (
            .O(N__17483),
            .I(N__17480));
    CascadeBuf I__3987 (
            .O(N__17480),
            .I(N__17477));
    CascadeMux I__3986 (
            .O(N__17477),
            .I(N__17474));
    CascadeBuf I__3985 (
            .O(N__17474),
            .I(N__17471));
    CascadeMux I__3984 (
            .O(N__17471),
            .I(N__17468));
    CascadeBuf I__3983 (
            .O(N__17468),
            .I(N__17465));
    CascadeMux I__3982 (
            .O(N__17465),
            .I(N__17462));
    CascadeBuf I__3981 (
            .O(N__17462),
            .I(N__17459));
    CascadeMux I__3980 (
            .O(N__17459),
            .I(N__17456));
    CascadeBuf I__3979 (
            .O(N__17456),
            .I(N__17453));
    CascadeMux I__3978 (
            .O(N__17453),
            .I(N__17450));
    CascadeBuf I__3977 (
            .O(N__17450),
            .I(N__17447));
    CascadeMux I__3976 (
            .O(N__17447),
            .I(N__17444));
    CascadeBuf I__3975 (
            .O(N__17444),
            .I(N__17441));
    CascadeMux I__3974 (
            .O(N__17441),
            .I(N__17438));
    CascadeBuf I__3973 (
            .O(N__17438),
            .I(N__17435));
    CascadeMux I__3972 (
            .O(N__17435),
            .I(N__17432));
    CascadeBuf I__3971 (
            .O(N__17432),
            .I(N__17429));
    CascadeMux I__3970 (
            .O(N__17429),
            .I(N__17426));
    CascadeBuf I__3969 (
            .O(N__17426),
            .I(N__17423));
    CascadeMux I__3968 (
            .O(N__17423),
            .I(N__17420));
    CascadeBuf I__3967 (
            .O(N__17420),
            .I(N__17417));
    CascadeMux I__3966 (
            .O(N__17417),
            .I(N__17414));
    CascadeBuf I__3965 (
            .O(N__17414),
            .I(N__17411));
    CascadeMux I__3964 (
            .O(N__17411),
            .I(N__17408));
    CascadeBuf I__3963 (
            .O(N__17408),
            .I(N__17405));
    CascadeMux I__3962 (
            .O(N__17405),
            .I(N__17402));
    CascadeBuf I__3961 (
            .O(N__17402),
            .I(N__17399));
    CascadeMux I__3960 (
            .O(N__17399),
            .I(N__17396));
    CascadeBuf I__3959 (
            .O(N__17396),
            .I(N__17393));
    CascadeMux I__3958 (
            .O(N__17393),
            .I(N__17390));
    InMux I__3957 (
            .O(N__17390),
            .I(N__17387));
    LocalMux I__3956 (
            .O(N__17387),
            .I(N__17384));
    Span4Mux_v I__3955 (
            .O(N__17384),
            .I(N__17381));
    Span4Mux_h I__3954 (
            .O(N__17381),
            .I(N__17378));
    Odrv4 I__3953 (
            .O(N__17378),
            .I(M_this_vga_signals_address_6));
    CEMux I__3952 (
            .O(N__17375),
            .I(N__17372));
    LocalMux I__3951 (
            .O(N__17372),
            .I(N__17368));
    CEMux I__3950 (
            .O(N__17371),
            .I(N__17365));
    Span4Mux_v I__3949 (
            .O(N__17368),
            .I(N__17360));
    LocalMux I__3948 (
            .O(N__17365),
            .I(N__17360));
    Span4Mux_v I__3947 (
            .O(N__17360),
            .I(N__17357));
    Span4Mux_v I__3946 (
            .O(N__17357),
            .I(N__17354));
    Odrv4 I__3945 (
            .O(N__17354),
            .I(\this_vram.mem_WE_12 ));
    InMux I__3944 (
            .O(N__17351),
            .I(N__17346));
    InMux I__3943 (
            .O(N__17350),
            .I(N__17343));
    InMux I__3942 (
            .O(N__17349),
            .I(N__17340));
    LocalMux I__3941 (
            .O(N__17346),
            .I(N__17334));
    LocalMux I__3940 (
            .O(N__17343),
            .I(N__17334));
    LocalMux I__3939 (
            .O(N__17340),
            .I(N__17331));
    InMux I__3938 (
            .O(N__17339),
            .I(N__17328));
    Span4Mux_v I__3937 (
            .O(N__17334),
            .I(N__17323));
    Span4Mux_h I__3936 (
            .O(N__17331),
            .I(N__17323));
    LocalMux I__3935 (
            .O(N__17328),
            .I(N__17315));
    Span4Mux_h I__3934 (
            .O(N__17323),
            .I(N__17312));
    InMux I__3933 (
            .O(N__17322),
            .I(N__17305));
    InMux I__3932 (
            .O(N__17321),
            .I(N__17305));
    InMux I__3931 (
            .O(N__17320),
            .I(N__17302));
    CascadeMux I__3930 (
            .O(N__17319),
            .I(N__17295));
    CascadeMux I__3929 (
            .O(N__17318),
            .I(N__17292));
    Span12Mux_h I__3928 (
            .O(N__17315),
            .I(N__17289));
    Span4Mux_h I__3927 (
            .O(N__17312),
            .I(N__17286));
    InMux I__3926 (
            .O(N__17311),
            .I(N__17281));
    InMux I__3925 (
            .O(N__17310),
            .I(N__17281));
    LocalMux I__3924 (
            .O(N__17305),
            .I(N__17278));
    LocalMux I__3923 (
            .O(N__17302),
            .I(N__17275));
    InMux I__3922 (
            .O(N__17301),
            .I(N__17266));
    InMux I__3921 (
            .O(N__17300),
            .I(N__17266));
    InMux I__3920 (
            .O(N__17299),
            .I(N__17266));
    InMux I__3919 (
            .O(N__17298),
            .I(N__17266));
    InMux I__3918 (
            .O(N__17295),
            .I(N__17263));
    InMux I__3917 (
            .O(N__17292),
            .I(N__17260));
    Odrv12 I__3916 (
            .O(N__17289),
            .I(\this_vga_signals.rgb_1_2 ));
    Odrv4 I__3915 (
            .O(N__17286),
            .I(\this_vga_signals.rgb_1_2 ));
    LocalMux I__3914 (
            .O(N__17281),
            .I(\this_vga_signals.rgb_1_2 ));
    Odrv4 I__3913 (
            .O(N__17278),
            .I(\this_vga_signals.rgb_1_2 ));
    Odrv4 I__3912 (
            .O(N__17275),
            .I(\this_vga_signals.rgb_1_2 ));
    LocalMux I__3911 (
            .O(N__17266),
            .I(\this_vga_signals.rgb_1_2 ));
    LocalMux I__3910 (
            .O(N__17263),
            .I(\this_vga_signals.rgb_1_2 ));
    LocalMux I__3909 (
            .O(N__17260),
            .I(\this_vga_signals.rgb_1_2 ));
    CEMux I__3908 (
            .O(N__17243),
            .I(N__17239));
    CEMux I__3907 (
            .O(N__17242),
            .I(N__17236));
    LocalMux I__3906 (
            .O(N__17239),
            .I(N__17233));
    LocalMux I__3905 (
            .O(N__17236),
            .I(N__17230));
    Span4Mux_v I__3904 (
            .O(N__17233),
            .I(N__17227));
    Span4Mux_h I__3903 (
            .O(N__17230),
            .I(N__17224));
    Odrv4 I__3902 (
            .O(N__17227),
            .I(\this_vram.mem_WE_8 ));
    Odrv4 I__3901 (
            .O(N__17224),
            .I(\this_vram.mem_WE_8 ));
    InMux I__3900 (
            .O(N__17219),
            .I(N__17216));
    LocalMux I__3899 (
            .O(N__17216),
            .I(N__17213));
    Span4Mux_v I__3898 (
            .O(N__17213),
            .I(N__17210));
    Span4Mux_v I__3897 (
            .O(N__17210),
            .I(N__17207));
    Span4Mux_v I__3896 (
            .O(N__17207),
            .I(N__17204));
    Odrv4 I__3895 (
            .O(N__17204),
            .I(\this_vram.mem_out_bus0_3 ));
    InMux I__3894 (
            .O(N__17201),
            .I(N__17194));
    InMux I__3893 (
            .O(N__17200),
            .I(N__17191));
    InMux I__3892 (
            .O(N__17199),
            .I(N__17188));
    InMux I__3891 (
            .O(N__17198),
            .I(N__17182));
    InMux I__3890 (
            .O(N__17197),
            .I(N__17182));
    LocalMux I__3889 (
            .O(N__17194),
            .I(N__17171));
    LocalMux I__3888 (
            .O(N__17191),
            .I(N__17171));
    LocalMux I__3887 (
            .O(N__17188),
            .I(N__17171));
    InMux I__3886 (
            .O(N__17187),
            .I(N__17165));
    LocalMux I__3885 (
            .O(N__17182),
            .I(N__17155));
    InMux I__3884 (
            .O(N__17181),
            .I(N__17152));
    InMux I__3883 (
            .O(N__17180),
            .I(N__17145));
    InMux I__3882 (
            .O(N__17179),
            .I(N__17145));
    InMux I__3881 (
            .O(N__17178),
            .I(N__17145));
    Span4Mux_v I__3880 (
            .O(N__17171),
            .I(N__17142));
    InMux I__3879 (
            .O(N__17170),
            .I(N__17139));
    InMux I__3878 (
            .O(N__17169),
            .I(N__17136));
    InMux I__3877 (
            .O(N__17168),
            .I(N__17133));
    LocalMux I__3876 (
            .O(N__17165),
            .I(N__17129));
    InMux I__3875 (
            .O(N__17164),
            .I(N__17126));
    InMux I__3874 (
            .O(N__17163),
            .I(N__17119));
    InMux I__3873 (
            .O(N__17162),
            .I(N__17119));
    InMux I__3872 (
            .O(N__17161),
            .I(N__17119));
    CascadeMux I__3871 (
            .O(N__17160),
            .I(N__17112));
    CascadeMux I__3870 (
            .O(N__17159),
            .I(N__17107));
    CascadeMux I__3869 (
            .O(N__17158),
            .I(N__17104));
    Span4Mux_h I__3868 (
            .O(N__17155),
            .I(N__17094));
    LocalMux I__3867 (
            .O(N__17152),
            .I(N__17094));
    LocalMux I__3866 (
            .O(N__17145),
            .I(N__17094));
    Sp12to4 I__3865 (
            .O(N__17142),
            .I(N__17087));
    LocalMux I__3864 (
            .O(N__17139),
            .I(N__17087));
    LocalMux I__3863 (
            .O(N__17136),
            .I(N__17087));
    LocalMux I__3862 (
            .O(N__17133),
            .I(N__17084));
    InMux I__3861 (
            .O(N__17132),
            .I(N__17081));
    Span4Mux_v I__3860 (
            .O(N__17129),
            .I(N__17074));
    LocalMux I__3859 (
            .O(N__17126),
            .I(N__17074));
    LocalMux I__3858 (
            .O(N__17119),
            .I(N__17074));
    InMux I__3857 (
            .O(N__17118),
            .I(N__17071));
    InMux I__3856 (
            .O(N__17117),
            .I(N__17064));
    InMux I__3855 (
            .O(N__17116),
            .I(N__17064));
    InMux I__3854 (
            .O(N__17115),
            .I(N__17064));
    InMux I__3853 (
            .O(N__17112),
            .I(N__17059));
    InMux I__3852 (
            .O(N__17111),
            .I(N__17059));
    InMux I__3851 (
            .O(N__17110),
            .I(N__17050));
    InMux I__3850 (
            .O(N__17107),
            .I(N__17050));
    InMux I__3849 (
            .O(N__17104),
            .I(N__17050));
    InMux I__3848 (
            .O(N__17103),
            .I(N__17050));
    InMux I__3847 (
            .O(N__17102),
            .I(N__17045));
    InMux I__3846 (
            .O(N__17101),
            .I(N__17045));
    Span4Mux_h I__3845 (
            .O(N__17094),
            .I(N__17042));
    Odrv12 I__3844 (
            .O(N__17087),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    Odrv4 I__3843 (
            .O(N__17084),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    LocalMux I__3842 (
            .O(N__17081),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    Odrv4 I__3841 (
            .O(N__17074),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    LocalMux I__3840 (
            .O(N__17071),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    LocalMux I__3839 (
            .O(N__17064),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    LocalMux I__3838 (
            .O(N__17059),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    LocalMux I__3837 (
            .O(N__17050),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    LocalMux I__3836 (
            .O(N__17045),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    Odrv4 I__3835 (
            .O(N__17042),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3));
    CascadeMux I__3834 (
            .O(N__17021),
            .I(N__17018));
    InMux I__3833 (
            .O(N__17018),
            .I(N__17015));
    LocalMux I__3832 (
            .O(N__17015),
            .I(rgb_1_cry_0_0_c_RNOZ0Z_0));
    InMux I__3831 (
            .O(N__17012),
            .I(N__17009));
    LocalMux I__3830 (
            .O(N__17009),
            .I(M_vcounter_q_esr_RNI1H9RHL_9));
    CascadeMux I__3829 (
            .O(N__17006),
            .I(N__17003));
    InMux I__3828 (
            .O(N__17003),
            .I(N__16994));
    InMux I__3827 (
            .O(N__17002),
            .I(N__16994));
    InMux I__3826 (
            .O(N__17001),
            .I(N__16987));
    InMux I__3825 (
            .O(N__17000),
            .I(N__16987));
    InMux I__3824 (
            .O(N__16999),
            .I(N__16987));
    LocalMux I__3823 (
            .O(N__16994),
            .I(N__16979));
    LocalMux I__3822 (
            .O(N__16987),
            .I(N__16979));
    InMux I__3821 (
            .O(N__16986),
            .I(N__16972));
    InMux I__3820 (
            .O(N__16985),
            .I(N__16972));
    InMux I__3819 (
            .O(N__16984),
            .I(N__16972));
    Span4Mux_v I__3818 (
            .O(N__16979),
            .I(N__16963));
    LocalMux I__3817 (
            .O(N__16972),
            .I(N__16960));
    InMux I__3816 (
            .O(N__16971),
            .I(N__16951));
    InMux I__3815 (
            .O(N__16970),
            .I(N__16951));
    InMux I__3814 (
            .O(N__16969),
            .I(N__16951));
    InMux I__3813 (
            .O(N__16968),
            .I(N__16951));
    InMux I__3812 (
            .O(N__16967),
            .I(N__16948));
    InMux I__3811 (
            .O(N__16966),
            .I(N__16945));
    Odrv4 I__3810 (
            .O(N__16963),
            .I(rgb_1_3));
    Odrv4 I__3809 (
            .O(N__16960),
            .I(rgb_1_3));
    LocalMux I__3808 (
            .O(N__16951),
            .I(rgb_1_3));
    LocalMux I__3807 (
            .O(N__16948),
            .I(rgb_1_3));
    LocalMux I__3806 (
            .O(N__16945),
            .I(rgb_1_3));
    CascadeMux I__3805 (
            .O(N__16934),
            .I(N__16928));
    CascadeMux I__3804 (
            .O(N__16933),
            .I(N__16925));
    CascadeMux I__3803 (
            .O(N__16932),
            .I(N__16921));
    InMux I__3802 (
            .O(N__16931),
            .I(N__16916));
    InMux I__3801 (
            .O(N__16928),
            .I(N__16916));
    InMux I__3800 (
            .O(N__16925),
            .I(N__16909));
    InMux I__3799 (
            .O(N__16924),
            .I(N__16909));
    InMux I__3798 (
            .O(N__16921),
            .I(N__16909));
    LocalMux I__3797 (
            .O(N__16916),
            .I(N__16898));
    LocalMux I__3796 (
            .O(N__16909),
            .I(N__16898));
    InMux I__3795 (
            .O(N__16908),
            .I(N__16891));
    InMux I__3794 (
            .O(N__16907),
            .I(N__16891));
    InMux I__3793 (
            .O(N__16906),
            .I(N__16891));
    CascadeMux I__3792 (
            .O(N__16905),
            .I(N__16888));
    CascadeMux I__3791 (
            .O(N__16904),
            .I(N__16884));
    CascadeMux I__3790 (
            .O(N__16903),
            .I(N__16881));
    Span4Mux_v I__3789 (
            .O(N__16898),
            .I(N__16876));
    LocalMux I__3788 (
            .O(N__16891),
            .I(N__16873));
    InMux I__3787 (
            .O(N__16888),
            .I(N__16864));
    InMux I__3786 (
            .O(N__16887),
            .I(N__16864));
    InMux I__3785 (
            .O(N__16884),
            .I(N__16864));
    InMux I__3784 (
            .O(N__16881),
            .I(N__16864));
    InMux I__3783 (
            .O(N__16880),
            .I(N__16861));
    InMux I__3782 (
            .O(N__16879),
            .I(N__16858));
    Odrv4 I__3781 (
            .O(N__16876),
            .I(rgb_1_4));
    Odrv4 I__3780 (
            .O(N__16873),
            .I(rgb_1_4));
    LocalMux I__3779 (
            .O(N__16864),
            .I(rgb_1_4));
    LocalMux I__3778 (
            .O(N__16861),
            .I(rgb_1_4));
    LocalMux I__3777 (
            .O(N__16858),
            .I(rgb_1_4));
    InMux I__3776 (
            .O(N__16847),
            .I(N__16837));
    InMux I__3775 (
            .O(N__16846),
            .I(N__16837));
    InMux I__3774 (
            .O(N__16845),
            .I(N__16830));
    InMux I__3773 (
            .O(N__16844),
            .I(N__16830));
    InMux I__3772 (
            .O(N__16843),
            .I(N__16830));
    CascadeMux I__3771 (
            .O(N__16842),
            .I(N__16827));
    LocalMux I__3770 (
            .O(N__16837),
            .I(N__16818));
    LocalMux I__3769 (
            .O(N__16830),
            .I(N__16818));
    InMux I__3768 (
            .O(N__16827),
            .I(N__16811));
    InMux I__3767 (
            .O(N__16826),
            .I(N__16811));
    InMux I__3766 (
            .O(N__16825),
            .I(N__16811));
    CascadeMux I__3765 (
            .O(N__16824),
            .I(N__16804));
    CascadeMux I__3764 (
            .O(N__16823),
            .I(N__16801));
    Span4Mux_v I__3763 (
            .O(N__16818),
            .I(N__16798));
    LocalMux I__3762 (
            .O(N__16811),
            .I(N__16795));
    InMux I__3761 (
            .O(N__16810),
            .I(N__16786));
    InMux I__3760 (
            .O(N__16809),
            .I(N__16786));
    InMux I__3759 (
            .O(N__16808),
            .I(N__16786));
    InMux I__3758 (
            .O(N__16807),
            .I(N__16786));
    InMux I__3757 (
            .O(N__16804),
            .I(N__16783));
    InMux I__3756 (
            .O(N__16801),
            .I(N__16780));
    Odrv4 I__3755 (
            .O(N__16798),
            .I(rgb_1_5));
    Odrv4 I__3754 (
            .O(N__16795),
            .I(rgb_1_5));
    LocalMux I__3753 (
            .O(N__16786),
            .I(rgb_1_5));
    LocalMux I__3752 (
            .O(N__16783),
            .I(rgb_1_5));
    LocalMux I__3751 (
            .O(N__16780),
            .I(rgb_1_5));
    CascadeMux I__3750 (
            .O(N__16769),
            .I(N__16763));
    InMux I__3749 (
            .O(N__16768),
            .I(N__16755));
    InMux I__3748 (
            .O(N__16767),
            .I(N__16755));
    InMux I__3747 (
            .O(N__16766),
            .I(N__16748));
    InMux I__3746 (
            .O(N__16763),
            .I(N__16748));
    InMux I__3745 (
            .O(N__16762),
            .I(N__16748));
    CascadeMux I__3744 (
            .O(N__16761),
            .I(N__16744));
    CascadeMux I__3743 (
            .O(N__16760),
            .I(N__16741));
    LocalMux I__3742 (
            .O(N__16755),
            .I(N__16735));
    LocalMux I__3741 (
            .O(N__16748),
            .I(N__16735));
    InMux I__3740 (
            .O(N__16747),
            .I(N__16728));
    InMux I__3739 (
            .O(N__16744),
            .I(N__16728));
    InMux I__3738 (
            .O(N__16741),
            .I(N__16728));
    CascadeMux I__3737 (
            .O(N__16740),
            .I(N__16724));
    Span4Mux_v I__3736 (
            .O(N__16735),
            .I(N__16717));
    LocalMux I__3735 (
            .O(N__16728),
            .I(N__16714));
    InMux I__3734 (
            .O(N__16727),
            .I(N__16705));
    InMux I__3733 (
            .O(N__16724),
            .I(N__16705));
    InMux I__3732 (
            .O(N__16723),
            .I(N__16705));
    InMux I__3731 (
            .O(N__16722),
            .I(N__16705));
    InMux I__3730 (
            .O(N__16721),
            .I(N__16702));
    InMux I__3729 (
            .O(N__16720),
            .I(N__16699));
    Odrv4 I__3728 (
            .O(N__16717),
            .I(rgb_1_6_THRU_CO));
    Odrv4 I__3727 (
            .O(N__16714),
            .I(rgb_1_6_THRU_CO));
    LocalMux I__3726 (
            .O(N__16705),
            .I(rgb_1_6_THRU_CO));
    LocalMux I__3725 (
            .O(N__16702),
            .I(rgb_1_6_THRU_CO));
    LocalMux I__3724 (
            .O(N__16699),
            .I(rgb_1_6_THRU_CO));
    InMux I__3723 (
            .O(N__16688),
            .I(N__16682));
    InMux I__3722 (
            .O(N__16687),
            .I(N__16682));
    LocalMux I__3721 (
            .O(N__16682),
            .I(m36));
    InMux I__3720 (
            .O(N__16679),
            .I(N__16675));
    InMux I__3719 (
            .O(N__16678),
            .I(N__16672));
    LocalMux I__3718 (
            .O(N__16675),
            .I(N__16669));
    LocalMux I__3717 (
            .O(N__16672),
            .I(N__16666));
    Span12Mux_h I__3716 (
            .O(N__16669),
            .I(N__16663));
    Span12Mux_v I__3715 (
            .O(N__16666),
            .I(N__16660));
    Odrv12 I__3714 (
            .O(N__16663),
            .I(port_address_c_0));
    Odrv12 I__3713 (
            .O(N__16660),
            .I(port_address_c_0));
    InMux I__3712 (
            .O(N__16655),
            .I(N__16652));
    LocalMux I__3711 (
            .O(N__16652),
            .I(N__16649));
    Span12Mux_h I__3710 (
            .O(N__16649),
            .I(N__16646));
    Odrv12 I__3709 (
            .O(N__16646),
            .I(port_address_c_1));
    InMux I__3708 (
            .O(N__16643),
            .I(N__16640));
    LocalMux I__3707 (
            .O(N__16640),
            .I(M_state_q_ns_0_a3_0_1_1));
    InMux I__3706 (
            .O(N__16637),
            .I(N__16632));
    InMux I__3705 (
            .O(N__16636),
            .I(N__16629));
    CascadeMux I__3704 (
            .O(N__16635),
            .I(N__16626));
    LocalMux I__3703 (
            .O(N__16632),
            .I(N__16623));
    LocalMux I__3702 (
            .O(N__16629),
            .I(N__16620));
    InMux I__3701 (
            .O(N__16626),
            .I(N__16617));
    Span4Mux_h I__3700 (
            .O(N__16623),
            .I(N__16614));
    Span4Mux_h I__3699 (
            .O(N__16620),
            .I(N__16611));
    LocalMux I__3698 (
            .O(N__16617),
            .I(N__16608));
    Span4Mux_v I__3697 (
            .O(N__16614),
            .I(N__16605));
    Span4Mux_v I__3696 (
            .O(N__16611),
            .I(N__16602));
    Span4Mux_h I__3695 (
            .O(N__16608),
            .I(N__16599));
    Span4Mux_v I__3694 (
            .O(N__16605),
            .I(N__16596));
    Span4Mux_v I__3693 (
            .O(N__16602),
            .I(N__16593));
    Span4Mux_v I__3692 (
            .O(N__16599),
            .I(N__16590));
    Span4Mux_h I__3691 (
            .O(N__16596),
            .I(N__16587));
    Span4Mux_v I__3690 (
            .O(N__16593),
            .I(N__16584));
    Span4Mux_v I__3689 (
            .O(N__16590),
            .I(N__16581));
    Odrv4 I__3688 (
            .O(N__16587),
            .I(port_data_c_1));
    Odrv4 I__3687 (
            .O(N__16584),
            .I(port_data_c_1));
    Odrv4 I__3686 (
            .O(N__16581),
            .I(port_data_c_1));
    InMux I__3685 (
            .O(N__16574),
            .I(N__16571));
    LocalMux I__3684 (
            .O(N__16571),
            .I(N__16567));
    InMux I__3683 (
            .O(N__16570),
            .I(N__16564));
    Span4Mux_h I__3682 (
            .O(N__16567),
            .I(N__16561));
    LocalMux I__3681 (
            .O(N__16564),
            .I(N__16558));
    Span4Mux_v I__3680 (
            .O(N__16561),
            .I(N__16551));
    Span4Mux_h I__3679 (
            .O(N__16558),
            .I(N__16551));
    InMux I__3678 (
            .O(N__16557),
            .I(N__16548));
    InMux I__3677 (
            .O(N__16556),
            .I(N__16543));
    Span4Mux_v I__3676 (
            .O(N__16551),
            .I(N__16539));
    LocalMux I__3675 (
            .O(N__16548),
            .I(N__16536));
    InMux I__3674 (
            .O(N__16547),
            .I(N__16533));
    InMux I__3673 (
            .O(N__16546),
            .I(N__16530));
    LocalMux I__3672 (
            .O(N__16543),
            .I(N__16527));
    InMux I__3671 (
            .O(N__16542),
            .I(N__16524));
    Span4Mux_v I__3670 (
            .O(N__16539),
            .I(N__16519));
    Span4Mux_h I__3669 (
            .O(N__16536),
            .I(N__16519));
    LocalMux I__3668 (
            .O(N__16533),
            .I(N__16516));
    LocalMux I__3667 (
            .O(N__16530),
            .I(N__16513));
    Span4Mux_v I__3666 (
            .O(N__16527),
            .I(N__16508));
    LocalMux I__3665 (
            .O(N__16524),
            .I(N__16508));
    Span4Mux_v I__3664 (
            .O(N__16519),
            .I(N__16502));
    Span4Mux_h I__3663 (
            .O(N__16516),
            .I(N__16502));
    Span12Mux_h I__3662 (
            .O(N__16513),
            .I(N__16499));
    Span4Mux_v I__3661 (
            .O(N__16508),
            .I(N__16496));
    InMux I__3660 (
            .O(N__16507),
            .I(N__16493));
    Span4Mux_h I__3659 (
            .O(N__16502),
            .I(N__16490));
    Span12Mux_v I__3658 (
            .O(N__16499),
            .I(N__16483));
    Sp12to4 I__3657 (
            .O(N__16496),
            .I(N__16483));
    LocalMux I__3656 (
            .O(N__16493),
            .I(N__16483));
    Odrv4 I__3655 (
            .O(N__16490),
            .I(M_this_vram_write_data_1));
    Odrv12 I__3654 (
            .O(N__16483),
            .I(M_this_vram_write_data_1));
    CascadeMux I__3653 (
            .O(N__16478),
            .I(N__16474));
    InMux I__3652 (
            .O(N__16477),
            .I(N__16466));
    InMux I__3651 (
            .O(N__16474),
            .I(N__16466));
    InMux I__3650 (
            .O(N__16473),
            .I(N__16463));
    InMux I__3649 (
            .O(N__16472),
            .I(N__16457));
    InMux I__3648 (
            .O(N__16471),
            .I(N__16454));
    LocalMux I__3647 (
            .O(N__16466),
            .I(N__16444));
    LocalMux I__3646 (
            .O(N__16463),
            .I(N__16444));
    InMux I__3645 (
            .O(N__16462),
            .I(N__16439));
    InMux I__3644 (
            .O(N__16461),
            .I(N__16439));
    InMux I__3643 (
            .O(N__16460),
            .I(N__16433));
    LocalMux I__3642 (
            .O(N__16457),
            .I(N__16430));
    LocalMux I__3641 (
            .O(N__16454),
            .I(N__16427));
    InMux I__3640 (
            .O(N__16453),
            .I(N__16422));
    InMux I__3639 (
            .O(N__16452),
            .I(N__16422));
    InMux I__3638 (
            .O(N__16451),
            .I(N__16419));
    InMux I__3637 (
            .O(N__16450),
            .I(N__16414));
    InMux I__3636 (
            .O(N__16449),
            .I(N__16414));
    Span4Mux_v I__3635 (
            .O(N__16444),
            .I(N__16411));
    LocalMux I__3634 (
            .O(N__16439),
            .I(N__16408));
    InMux I__3633 (
            .O(N__16438),
            .I(N__16401));
    InMux I__3632 (
            .O(N__16437),
            .I(N__16401));
    InMux I__3631 (
            .O(N__16436),
            .I(N__16401));
    LocalMux I__3630 (
            .O(N__16433),
            .I(N__16396));
    Span4Mux_h I__3629 (
            .O(N__16430),
            .I(N__16396));
    Span4Mux_v I__3628 (
            .O(N__16427),
            .I(N__16391));
    LocalMux I__3627 (
            .O(N__16422),
            .I(N__16391));
    LocalMux I__3626 (
            .O(N__16419),
            .I(N_349_0));
    LocalMux I__3625 (
            .O(N__16414),
            .I(N_349_0));
    Odrv4 I__3624 (
            .O(N__16411),
            .I(N_349_0));
    Odrv4 I__3623 (
            .O(N__16408),
            .I(N_349_0));
    LocalMux I__3622 (
            .O(N__16401),
            .I(N_349_0));
    Odrv4 I__3621 (
            .O(N__16396),
            .I(N_349_0));
    Odrv4 I__3620 (
            .O(N__16391),
            .I(N_349_0));
    CascadeMux I__3619 (
            .O(N__16376),
            .I(N__16372));
    CascadeMux I__3618 (
            .O(N__16375),
            .I(N__16369));
    InMux I__3617 (
            .O(N__16372),
            .I(N__16366));
    InMux I__3616 (
            .O(N__16369),
            .I(N__16363));
    LocalMux I__3615 (
            .O(N__16366),
            .I(N__16360));
    LocalMux I__3614 (
            .O(N__16363),
            .I(N__16357));
    Span4Mux_v I__3613 (
            .O(N__16360),
            .I(N__16354));
    Span4Mux_v I__3612 (
            .O(N__16357),
            .I(N__16351));
    Sp12to4 I__3611 (
            .O(N__16354),
            .I(N__16348));
    Sp12to4 I__3610 (
            .O(N__16351),
            .I(N__16345));
    Span12Mux_h I__3609 (
            .O(N__16348),
            .I(N__16342));
    Span12Mux_h I__3608 (
            .O(N__16345),
            .I(N__16339));
    Span12Mux_v I__3607 (
            .O(N__16342),
            .I(N__16336));
    Span12Mux_v I__3606 (
            .O(N__16339),
            .I(N__16333));
    Odrv12 I__3605 (
            .O(N__16336),
            .I(port_data_c_6));
    Odrv12 I__3604 (
            .O(N__16333),
            .I(port_data_c_6));
    InMux I__3603 (
            .O(N__16328),
            .I(N__16322));
    InMux I__3602 (
            .O(N__16327),
            .I(N__16306));
    InMux I__3601 (
            .O(N__16326),
            .I(N__16303));
    CascadeMux I__3600 (
            .O(N__16325),
            .I(N__16291));
    LocalMux I__3599 (
            .O(N__16322),
            .I(N__16288));
    InMux I__3598 (
            .O(N__16321),
            .I(N__16281));
    InMux I__3597 (
            .O(N__16320),
            .I(N__16270));
    InMux I__3596 (
            .O(N__16319),
            .I(N__16270));
    InMux I__3595 (
            .O(N__16318),
            .I(N__16270));
    InMux I__3594 (
            .O(N__16317),
            .I(N__16270));
    InMux I__3593 (
            .O(N__16316),
            .I(N__16270));
    InMux I__3592 (
            .O(N__16315),
            .I(N__16267));
    InMux I__3591 (
            .O(N__16314),
            .I(N__16258));
    InMux I__3590 (
            .O(N__16313),
            .I(N__16258));
    InMux I__3589 (
            .O(N__16312),
            .I(N__16258));
    InMux I__3588 (
            .O(N__16311),
            .I(N__16258));
    CascadeMux I__3587 (
            .O(N__16310),
            .I(N__16255));
    InMux I__3586 (
            .O(N__16309),
            .I(N__16252));
    LocalMux I__3585 (
            .O(N__16306),
            .I(N__16247));
    LocalMux I__3584 (
            .O(N__16303),
            .I(N__16247));
    InMux I__3583 (
            .O(N__16302),
            .I(N__16242));
    InMux I__3582 (
            .O(N__16301),
            .I(N__16242));
    InMux I__3581 (
            .O(N__16300),
            .I(N__16235));
    InMux I__3580 (
            .O(N__16299),
            .I(N__16235));
    InMux I__3579 (
            .O(N__16298),
            .I(N__16224));
    InMux I__3578 (
            .O(N__16297),
            .I(N__16224));
    InMux I__3577 (
            .O(N__16296),
            .I(N__16224));
    InMux I__3576 (
            .O(N__16295),
            .I(N__16224));
    InMux I__3575 (
            .O(N__16294),
            .I(N__16224));
    InMux I__3574 (
            .O(N__16291),
            .I(N__16221));
    Span4Mux_h I__3573 (
            .O(N__16288),
            .I(N__16218));
    InMux I__3572 (
            .O(N__16287),
            .I(N__16215));
    InMux I__3571 (
            .O(N__16286),
            .I(N__16208));
    InMux I__3570 (
            .O(N__16285),
            .I(N__16208));
    InMux I__3569 (
            .O(N__16284),
            .I(N__16208));
    LocalMux I__3568 (
            .O(N__16281),
            .I(N__16199));
    LocalMux I__3567 (
            .O(N__16270),
            .I(N__16199));
    LocalMux I__3566 (
            .O(N__16267),
            .I(N__16199));
    LocalMux I__3565 (
            .O(N__16258),
            .I(N__16199));
    InMux I__3564 (
            .O(N__16255),
            .I(N__16196));
    LocalMux I__3563 (
            .O(N__16252),
            .I(N__16193));
    Span4Mux_v I__3562 (
            .O(N__16247),
            .I(N__16188));
    LocalMux I__3561 (
            .O(N__16242),
            .I(N__16188));
    InMux I__3560 (
            .O(N__16241),
            .I(N__16183));
    InMux I__3559 (
            .O(N__16240),
            .I(N__16183));
    LocalMux I__3558 (
            .O(N__16235),
            .I(M_state_qZ0Z_0));
    LocalMux I__3557 (
            .O(N__16224),
            .I(M_state_qZ0Z_0));
    LocalMux I__3556 (
            .O(N__16221),
            .I(M_state_qZ0Z_0));
    Odrv4 I__3555 (
            .O(N__16218),
            .I(M_state_qZ0Z_0));
    LocalMux I__3554 (
            .O(N__16215),
            .I(M_state_qZ0Z_0));
    LocalMux I__3553 (
            .O(N__16208),
            .I(M_state_qZ0Z_0));
    Odrv4 I__3552 (
            .O(N__16199),
            .I(M_state_qZ0Z_0));
    LocalMux I__3551 (
            .O(N__16196),
            .I(M_state_qZ0Z_0));
    Odrv4 I__3550 (
            .O(N__16193),
            .I(M_state_qZ0Z_0));
    Odrv4 I__3549 (
            .O(N__16188),
            .I(M_state_qZ0Z_0));
    LocalMux I__3548 (
            .O(N__16183),
            .I(M_state_qZ0Z_0));
    CascadeMux I__3547 (
            .O(N__16160),
            .I(N__16157));
    InMux I__3546 (
            .O(N__16157),
            .I(N__16154));
    LocalMux I__3545 (
            .O(N__16154),
            .I(N__16151));
    Odrv4 I__3544 (
            .O(N__16151),
            .I(N_414));
    InMux I__3543 (
            .O(N__16148),
            .I(N__16143));
    CascadeMux I__3542 (
            .O(N__16147),
            .I(N__16137));
    CascadeMux I__3541 (
            .O(N__16146),
            .I(N__16133));
    LocalMux I__3540 (
            .O(N__16143),
            .I(N__16130));
    InMux I__3539 (
            .O(N__16142),
            .I(N__16125));
    InMux I__3538 (
            .O(N__16141),
            .I(N__16125));
    InMux I__3537 (
            .O(N__16140),
            .I(N__16122));
    InMux I__3536 (
            .O(N__16137),
            .I(N__16114));
    InMux I__3535 (
            .O(N__16136),
            .I(N__16114));
    InMux I__3534 (
            .O(N__16133),
            .I(N__16114));
    Span4Mux_h I__3533 (
            .O(N__16130),
            .I(N__16107));
    LocalMux I__3532 (
            .O(N__16125),
            .I(N__16107));
    LocalMux I__3531 (
            .O(N__16122),
            .I(N__16107));
    InMux I__3530 (
            .O(N__16121),
            .I(N__16104));
    LocalMux I__3529 (
            .O(N__16114),
            .I(N__16101));
    Odrv4 I__3528 (
            .O(N__16107),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1));
    LocalMux I__3527 (
            .O(N__16104),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1));
    Odrv4 I__3526 (
            .O(N__16101),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1));
    InMux I__3525 (
            .O(N__16094),
            .I(N__16090));
    InMux I__3524 (
            .O(N__16093),
            .I(N__16079));
    LocalMux I__3523 (
            .O(N__16090),
            .I(N__16076));
    InMux I__3522 (
            .O(N__16089),
            .I(N__16069));
    InMux I__3521 (
            .O(N__16088),
            .I(N__16069));
    InMux I__3520 (
            .O(N__16087),
            .I(N__16069));
    InMux I__3519 (
            .O(N__16086),
            .I(N__16062));
    InMux I__3518 (
            .O(N__16085),
            .I(N__16062));
    InMux I__3517 (
            .O(N__16084),
            .I(N__16062));
    InMux I__3516 (
            .O(N__16083),
            .I(N__16051));
    InMux I__3515 (
            .O(N__16082),
            .I(N__16051));
    LocalMux I__3514 (
            .O(N__16079),
            .I(N__16042));
    Span4Mux_h I__3513 (
            .O(N__16076),
            .I(N__16042));
    LocalMux I__3512 (
            .O(N__16069),
            .I(N__16042));
    LocalMux I__3511 (
            .O(N__16062),
            .I(N__16042));
    InMux I__3510 (
            .O(N__16061),
            .I(N__16033));
    InMux I__3509 (
            .O(N__16060),
            .I(N__16033));
    InMux I__3508 (
            .O(N__16059),
            .I(N__16033));
    InMux I__3507 (
            .O(N__16058),
            .I(N__16033));
    InMux I__3506 (
            .O(N__16057),
            .I(N__16028));
    InMux I__3505 (
            .O(N__16056),
            .I(N__16028));
    LocalMux I__3504 (
            .O(N__16051),
            .I(this_vga_signals_un16_address_if_i1_mux_0));
    Odrv4 I__3503 (
            .O(N__16042),
            .I(this_vga_signals_un16_address_if_i1_mux_0));
    LocalMux I__3502 (
            .O(N__16033),
            .I(this_vga_signals_un16_address_if_i1_mux_0));
    LocalMux I__3501 (
            .O(N__16028),
            .I(this_vga_signals_un16_address_if_i1_mux_0));
    CascadeMux I__3500 (
            .O(N__16019),
            .I(N__16016));
    CascadeBuf I__3499 (
            .O(N__16016),
            .I(N__16013));
    CascadeMux I__3498 (
            .O(N__16013),
            .I(N__16010));
    CascadeBuf I__3497 (
            .O(N__16010),
            .I(N__16007));
    CascadeMux I__3496 (
            .O(N__16007),
            .I(N__16004));
    CascadeBuf I__3495 (
            .O(N__16004),
            .I(N__16001));
    CascadeMux I__3494 (
            .O(N__16001),
            .I(N__15998));
    CascadeBuf I__3493 (
            .O(N__15998),
            .I(N__15995));
    CascadeMux I__3492 (
            .O(N__15995),
            .I(N__15992));
    CascadeBuf I__3491 (
            .O(N__15992),
            .I(N__15989));
    CascadeMux I__3490 (
            .O(N__15989),
            .I(N__15986));
    CascadeBuf I__3489 (
            .O(N__15986),
            .I(N__15983));
    CascadeMux I__3488 (
            .O(N__15983),
            .I(N__15980));
    CascadeBuf I__3487 (
            .O(N__15980),
            .I(N__15977));
    CascadeMux I__3486 (
            .O(N__15977),
            .I(N__15974));
    CascadeBuf I__3485 (
            .O(N__15974),
            .I(N__15971));
    CascadeMux I__3484 (
            .O(N__15971),
            .I(N__15968));
    CascadeBuf I__3483 (
            .O(N__15968),
            .I(N__15965));
    CascadeMux I__3482 (
            .O(N__15965),
            .I(N__15962));
    CascadeBuf I__3481 (
            .O(N__15962),
            .I(N__15959));
    CascadeMux I__3480 (
            .O(N__15959),
            .I(N__15956));
    CascadeBuf I__3479 (
            .O(N__15956),
            .I(N__15953));
    CascadeMux I__3478 (
            .O(N__15953),
            .I(N__15950));
    CascadeBuf I__3477 (
            .O(N__15950),
            .I(N__15947));
    CascadeMux I__3476 (
            .O(N__15947),
            .I(N__15944));
    CascadeBuf I__3475 (
            .O(N__15944),
            .I(N__15941));
    CascadeMux I__3474 (
            .O(N__15941),
            .I(N__15938));
    CascadeBuf I__3473 (
            .O(N__15938),
            .I(N__15935));
    CascadeMux I__3472 (
            .O(N__15935),
            .I(N__15932));
    CascadeBuf I__3471 (
            .O(N__15932),
            .I(N__15929));
    CascadeMux I__3470 (
            .O(N__15929),
            .I(N__15926));
    InMux I__3469 (
            .O(N__15926),
            .I(N__15923));
    LocalMux I__3468 (
            .O(N__15923),
            .I(N__15920));
    Span12Mux_h I__3467 (
            .O(N__15920),
            .I(N__15916));
    InMux I__3466 (
            .O(N__15919),
            .I(N__15913));
    Span12Mux_v I__3465 (
            .O(N__15916),
            .I(N__15910));
    LocalMux I__3464 (
            .O(N__15913),
            .I(M_this_vga_signals_address_10));
    Odrv12 I__3463 (
            .O(N__15910),
            .I(M_this_vga_signals_address_10));
    InMux I__3462 (
            .O(N__15905),
            .I(N__15899));
    InMux I__3461 (
            .O(N__15904),
            .I(N__15896));
    InMux I__3460 (
            .O(N__15903),
            .I(N__15893));
    InMux I__3459 (
            .O(N__15902),
            .I(N__15890));
    LocalMux I__3458 (
            .O(N__15899),
            .I(N__15887));
    LocalMux I__3457 (
            .O(N__15896),
            .I(N__15882));
    LocalMux I__3456 (
            .O(N__15893),
            .I(N__15882));
    LocalMux I__3455 (
            .O(N__15890),
            .I(N__15876));
    Span4Mux_v I__3454 (
            .O(N__15887),
            .I(N__15871));
    Span4Mux_v I__3453 (
            .O(N__15882),
            .I(N__15871));
    InMux I__3452 (
            .O(N__15881),
            .I(N__15866));
    InMux I__3451 (
            .O(N__15880),
            .I(N__15866));
    CascadeMux I__3450 (
            .O(N__15879),
            .I(N__15863));
    Span4Mux_v I__3449 (
            .O(N__15876),
            .I(N__15860));
    Sp12to4 I__3448 (
            .O(N__15871),
            .I(N__15855));
    LocalMux I__3447 (
            .O(N__15866),
            .I(N__15855));
    InMux I__3446 (
            .O(N__15863),
            .I(N__15852));
    Sp12to4 I__3445 (
            .O(N__15860),
            .I(N__15845));
    Span12Mux_h I__3444 (
            .O(N__15855),
            .I(N__15845));
    LocalMux I__3443 (
            .O(N__15852),
            .I(N__15845));
    Odrv12 I__3442 (
            .O(N__15845),
            .I(M_this_vram_read_data_2));
    InMux I__3441 (
            .O(N__15842),
            .I(N__15833));
    InMux I__3440 (
            .O(N__15841),
            .I(N__15830));
    InMux I__3439 (
            .O(N__15840),
            .I(N__15825));
    InMux I__3438 (
            .O(N__15839),
            .I(N__15825));
    InMux I__3437 (
            .O(N__15838),
            .I(N__15820));
    InMux I__3436 (
            .O(N__15837),
            .I(N__15820));
    InMux I__3435 (
            .O(N__15836),
            .I(N__15817));
    LocalMux I__3434 (
            .O(N__15833),
            .I(N__15807));
    LocalMux I__3433 (
            .O(N__15830),
            .I(N__15807));
    LocalMux I__3432 (
            .O(N__15825),
            .I(N__15807));
    LocalMux I__3431 (
            .O(N__15820),
            .I(N__15807));
    LocalMux I__3430 (
            .O(N__15817),
            .I(N__15804));
    InMux I__3429 (
            .O(N__15816),
            .I(N__15801));
    Span4Mux_v I__3428 (
            .O(N__15807),
            .I(N__15797));
    Span4Mux_v I__3427 (
            .O(N__15804),
            .I(N__15794));
    LocalMux I__3426 (
            .O(N__15801),
            .I(N__15791));
    InMux I__3425 (
            .O(N__15800),
            .I(N__15788));
    Sp12to4 I__3424 (
            .O(N__15797),
            .I(N__15783));
    Sp12to4 I__3423 (
            .O(N__15794),
            .I(N__15783));
    Span4Mux_v I__3422 (
            .O(N__15791),
            .I(N__15778));
    LocalMux I__3421 (
            .O(N__15788),
            .I(N__15778));
    Odrv12 I__3420 (
            .O(N__15783),
            .I(this_vram_mem_radreg_11));
    Odrv4 I__3419 (
            .O(N__15778),
            .I(this_vram_mem_radreg_11));
    InMux I__3418 (
            .O(N__15773),
            .I(N__15770));
    LocalMux I__3417 (
            .O(N__15770),
            .I(mem_radreg_RNIMTEJ4_11));
    InMux I__3416 (
            .O(N__15767),
            .I(N__15764));
    LocalMux I__3415 (
            .O(N__15764),
            .I(m14));
    InMux I__3414 (
            .O(N__15761),
            .I(N__15758));
    LocalMux I__3413 (
            .O(N__15758),
            .I(rgb_1_cry_0_0_c_RNOZ0));
    InMux I__3412 (
            .O(N__15755),
            .I(N__15752));
    LocalMux I__3411 (
            .O(N__15752),
            .I(M_vcounter_q_esr_RNIB9J4TN_9));
    CascadeMux I__3410 (
            .O(N__15749),
            .I(N__15746));
    InMux I__3409 (
            .O(N__15746),
            .I(N__15743));
    LocalMux I__3408 (
            .O(N__15743),
            .I(N__15740));
    Odrv4 I__3407 (
            .O(N__15740),
            .I(M_vcounter_q_esr_RNICJRF0D_9));
    InMux I__3406 (
            .O(N__15737),
            .I(rgb_1_cry_0));
    InMux I__3405 (
            .O(N__15734),
            .I(rgb_1_cry_1));
    InMux I__3404 (
            .O(N__15731),
            .I(rgb_1_cry_2));
    InMux I__3403 (
            .O(N__15728),
            .I(rgb_1_6));
    CascadeMux I__3402 (
            .O(N__15725),
            .I(N_403_cascade_));
    InMux I__3401 (
            .O(N__15722),
            .I(N__15719));
    LocalMux I__3400 (
            .O(N__15719),
            .I(N__15716));
    Span4Mux_h I__3399 (
            .O(N__15716),
            .I(N__15713));
    Odrv4 I__3398 (
            .O(N__15713),
            .I(M_current_address_q_RNO_1Z0Z_2));
    CascadeMux I__3397 (
            .O(N__15710),
            .I(N__15707));
    CascadeBuf I__3396 (
            .O(N__15707),
            .I(N__15704));
    CascadeMux I__3395 (
            .O(N__15704),
            .I(N__15701));
    CascadeBuf I__3394 (
            .O(N__15701),
            .I(N__15698));
    CascadeMux I__3393 (
            .O(N__15698),
            .I(N__15695));
    CascadeBuf I__3392 (
            .O(N__15695),
            .I(N__15692));
    CascadeMux I__3391 (
            .O(N__15692),
            .I(N__15689));
    CascadeBuf I__3390 (
            .O(N__15689),
            .I(N__15686));
    CascadeMux I__3389 (
            .O(N__15686),
            .I(N__15683));
    CascadeBuf I__3388 (
            .O(N__15683),
            .I(N__15680));
    CascadeMux I__3387 (
            .O(N__15680),
            .I(N__15677));
    CascadeBuf I__3386 (
            .O(N__15677),
            .I(N__15674));
    CascadeMux I__3385 (
            .O(N__15674),
            .I(N__15671));
    CascadeBuf I__3384 (
            .O(N__15671),
            .I(N__15668));
    CascadeMux I__3383 (
            .O(N__15668),
            .I(N__15665));
    CascadeBuf I__3382 (
            .O(N__15665),
            .I(N__15662));
    CascadeMux I__3381 (
            .O(N__15662),
            .I(N__15659));
    CascadeBuf I__3380 (
            .O(N__15659),
            .I(N__15656));
    CascadeMux I__3379 (
            .O(N__15656),
            .I(N__15653));
    CascadeBuf I__3378 (
            .O(N__15653),
            .I(N__15650));
    CascadeMux I__3377 (
            .O(N__15650),
            .I(N__15647));
    CascadeBuf I__3376 (
            .O(N__15647),
            .I(N__15644));
    CascadeMux I__3375 (
            .O(N__15644),
            .I(N__15641));
    CascadeBuf I__3374 (
            .O(N__15641),
            .I(N__15638));
    CascadeMux I__3373 (
            .O(N__15638),
            .I(N__15635));
    CascadeBuf I__3372 (
            .O(N__15635),
            .I(N__15632));
    CascadeMux I__3371 (
            .O(N__15632),
            .I(N__15629));
    CascadeBuf I__3370 (
            .O(N__15629),
            .I(N__15626));
    CascadeMux I__3369 (
            .O(N__15626),
            .I(N__15623));
    CascadeBuf I__3368 (
            .O(N__15623),
            .I(N__15620));
    CascadeMux I__3367 (
            .O(N__15620),
            .I(N__15616));
    InMux I__3366 (
            .O(N__15619),
            .I(N__15613));
    InMux I__3365 (
            .O(N__15616),
            .I(N__15610));
    LocalMux I__3364 (
            .O(N__15613),
            .I(N__15607));
    LocalMux I__3363 (
            .O(N__15610),
            .I(N__15603));
    Span4Mux_h I__3362 (
            .O(N__15607),
            .I(N__15600));
    InMux I__3361 (
            .O(N__15606),
            .I(N__15597));
    Span12Mux_h I__3360 (
            .O(N__15603),
            .I(N__15594));
    Odrv4 I__3359 (
            .O(N__15600),
            .I(M_current_address_qZ0Z_2));
    LocalMux I__3358 (
            .O(N__15597),
            .I(M_current_address_qZ0Z_2));
    Odrv12 I__3357 (
            .O(N__15594),
            .I(M_current_address_qZ0Z_2));
    InMux I__3356 (
            .O(N__15587),
            .I(N__15584));
    LocalMux I__3355 (
            .O(N__15584),
            .I(N__15581));
    Odrv4 I__3354 (
            .O(N__15581),
            .I(M_current_address_q_RNO_1Z0Z_13));
    CascadeMux I__3353 (
            .O(N__15578),
            .I(N__15570));
    CascadeMux I__3352 (
            .O(N__15577),
            .I(N__15566));
    InMux I__3351 (
            .O(N__15576),
            .I(N__15559));
    InMux I__3350 (
            .O(N__15575),
            .I(N__15548));
    InMux I__3349 (
            .O(N__15574),
            .I(N__15548));
    InMux I__3348 (
            .O(N__15573),
            .I(N__15548));
    InMux I__3347 (
            .O(N__15570),
            .I(N__15541));
    InMux I__3346 (
            .O(N__15569),
            .I(N__15541));
    InMux I__3345 (
            .O(N__15566),
            .I(N__15541));
    InMux I__3344 (
            .O(N__15565),
            .I(N__15538));
    InMux I__3343 (
            .O(N__15564),
            .I(N__15531));
    InMux I__3342 (
            .O(N__15563),
            .I(N__15531));
    InMux I__3341 (
            .O(N__15562),
            .I(N__15531));
    LocalMux I__3340 (
            .O(N__15559),
            .I(N__15526));
    InMux I__3339 (
            .O(N__15558),
            .I(N__15523));
    InMux I__3338 (
            .O(N__15557),
            .I(N__15517));
    InMux I__3337 (
            .O(N__15556),
            .I(N__15517));
    InMux I__3336 (
            .O(N__15555),
            .I(N__15514));
    LocalMux I__3335 (
            .O(N__15548),
            .I(N__15511));
    LocalMux I__3334 (
            .O(N__15541),
            .I(N__15504));
    LocalMux I__3333 (
            .O(N__15538),
            .I(N__15504));
    LocalMux I__3332 (
            .O(N__15531),
            .I(N__15504));
    InMux I__3331 (
            .O(N__15530),
            .I(N__15501));
    InMux I__3330 (
            .O(N__15529),
            .I(N__15498));
    Span4Mux_v I__3329 (
            .O(N__15526),
            .I(N__15493));
    LocalMux I__3328 (
            .O(N__15523),
            .I(N__15493));
    InMux I__3327 (
            .O(N__15522),
            .I(N__15490));
    LocalMux I__3326 (
            .O(N__15517),
            .I(M_state_qZ0Z_1));
    LocalMux I__3325 (
            .O(N__15514),
            .I(M_state_qZ0Z_1));
    Odrv4 I__3324 (
            .O(N__15511),
            .I(M_state_qZ0Z_1));
    Odrv4 I__3323 (
            .O(N__15504),
            .I(M_state_qZ0Z_1));
    LocalMux I__3322 (
            .O(N__15501),
            .I(M_state_qZ0Z_1));
    LocalMux I__3321 (
            .O(N__15498),
            .I(M_state_qZ0Z_1));
    Odrv4 I__3320 (
            .O(N__15493),
            .I(M_state_qZ0Z_1));
    LocalMux I__3319 (
            .O(N__15490),
            .I(M_state_qZ0Z_1));
    CascadeMux I__3318 (
            .O(N__15473),
            .I(N_407_cascade_));
    InMux I__3317 (
            .O(N__15470),
            .I(N__15467));
    LocalMux I__3316 (
            .O(N__15467),
            .I(N__15464));
    Span4Mux_h I__3315 (
            .O(N__15464),
            .I(N__15461));
    Odrv4 I__3314 (
            .O(N__15461),
            .I(M_current_address_q_RNO_1Z0Z_6));
    CascadeMux I__3313 (
            .O(N__15458),
            .I(N__15455));
    CascadeBuf I__3312 (
            .O(N__15455),
            .I(N__15452));
    CascadeMux I__3311 (
            .O(N__15452),
            .I(N__15449));
    CascadeBuf I__3310 (
            .O(N__15449),
            .I(N__15446));
    CascadeMux I__3309 (
            .O(N__15446),
            .I(N__15443));
    CascadeBuf I__3308 (
            .O(N__15443),
            .I(N__15440));
    CascadeMux I__3307 (
            .O(N__15440),
            .I(N__15437));
    CascadeBuf I__3306 (
            .O(N__15437),
            .I(N__15434));
    CascadeMux I__3305 (
            .O(N__15434),
            .I(N__15431));
    CascadeBuf I__3304 (
            .O(N__15431),
            .I(N__15428));
    CascadeMux I__3303 (
            .O(N__15428),
            .I(N__15425));
    CascadeBuf I__3302 (
            .O(N__15425),
            .I(N__15422));
    CascadeMux I__3301 (
            .O(N__15422),
            .I(N__15419));
    CascadeBuf I__3300 (
            .O(N__15419),
            .I(N__15416));
    CascadeMux I__3299 (
            .O(N__15416),
            .I(N__15413));
    CascadeBuf I__3298 (
            .O(N__15413),
            .I(N__15410));
    CascadeMux I__3297 (
            .O(N__15410),
            .I(N__15407));
    CascadeBuf I__3296 (
            .O(N__15407),
            .I(N__15404));
    CascadeMux I__3295 (
            .O(N__15404),
            .I(N__15401));
    CascadeBuf I__3294 (
            .O(N__15401),
            .I(N__15398));
    CascadeMux I__3293 (
            .O(N__15398),
            .I(N__15395));
    CascadeBuf I__3292 (
            .O(N__15395),
            .I(N__15392));
    CascadeMux I__3291 (
            .O(N__15392),
            .I(N__15389));
    CascadeBuf I__3290 (
            .O(N__15389),
            .I(N__15386));
    CascadeMux I__3289 (
            .O(N__15386),
            .I(N__15383));
    CascadeBuf I__3288 (
            .O(N__15383),
            .I(N__15380));
    CascadeMux I__3287 (
            .O(N__15380),
            .I(N__15377));
    CascadeBuf I__3286 (
            .O(N__15377),
            .I(N__15374));
    CascadeMux I__3285 (
            .O(N__15374),
            .I(N__15371));
    CascadeBuf I__3284 (
            .O(N__15371),
            .I(N__15368));
    CascadeMux I__3283 (
            .O(N__15368),
            .I(N__15365));
    InMux I__3282 (
            .O(N__15365),
            .I(N__15362));
    LocalMux I__3281 (
            .O(N__15362),
            .I(N__15359));
    Span4Mux_s2_v I__3280 (
            .O(N__15359),
            .I(N__15355));
    InMux I__3279 (
            .O(N__15358),
            .I(N__15352));
    Span4Mux_h I__3278 (
            .O(N__15355),
            .I(N__15349));
    LocalMux I__3277 (
            .O(N__15352),
            .I(N__15346));
    Span4Mux_v I__3276 (
            .O(N__15349),
            .I(N__15342));
    Span4Mux_h I__3275 (
            .O(N__15346),
            .I(N__15339));
    InMux I__3274 (
            .O(N__15345),
            .I(N__15336));
    Span4Mux_v I__3273 (
            .O(N__15342),
            .I(N__15333));
    Odrv4 I__3272 (
            .O(N__15339),
            .I(M_current_address_qZ0Z_6));
    LocalMux I__3271 (
            .O(N__15336),
            .I(M_current_address_qZ0Z_6));
    Odrv4 I__3270 (
            .O(N__15333),
            .I(M_current_address_qZ0Z_6));
    InMux I__3269 (
            .O(N__15326),
            .I(N__15316));
    InMux I__3268 (
            .O(N__15325),
            .I(N__15316));
    SRMux I__3267 (
            .O(N__15324),
            .I(N__15313));
    SRMux I__3266 (
            .O(N__15323),
            .I(N__15309));
    SRMux I__3265 (
            .O(N__15322),
            .I(N__15303));
    SRMux I__3264 (
            .O(N__15321),
            .I(N__15300));
    LocalMux I__3263 (
            .O(N__15316),
            .I(N__15295));
    LocalMux I__3262 (
            .O(N__15313),
            .I(N__15295));
    SRMux I__3261 (
            .O(N__15312),
            .I(N__15292));
    LocalMux I__3260 (
            .O(N__15309),
            .I(N__15289));
    InMux I__3259 (
            .O(N__15308),
            .I(N__15286));
    SRMux I__3258 (
            .O(N__15307),
            .I(N__15283));
    InMux I__3257 (
            .O(N__15306),
            .I(N__15280));
    LocalMux I__3256 (
            .O(N__15303),
            .I(N__15277));
    LocalMux I__3255 (
            .O(N__15300),
            .I(N__15274));
    Span4Mux_v I__3254 (
            .O(N__15295),
            .I(N__15271));
    LocalMux I__3253 (
            .O(N__15292),
            .I(N__15264));
    Span4Mux_v I__3252 (
            .O(N__15289),
            .I(N__15264));
    LocalMux I__3251 (
            .O(N__15286),
            .I(N__15264));
    LocalMux I__3250 (
            .O(N__15283),
            .I(N__15261));
    LocalMux I__3249 (
            .O(N__15280),
            .I(N__15258));
    Span4Mux_h I__3248 (
            .O(N__15277),
            .I(N__15249));
    Span4Mux_v I__3247 (
            .O(N__15274),
            .I(N__15249));
    Span4Mux_h I__3246 (
            .O(N__15271),
            .I(N__15249));
    Span4Mux_v I__3245 (
            .O(N__15264),
            .I(N__15244));
    Span4Mux_h I__3244 (
            .O(N__15261),
            .I(N__15244));
    Span4Mux_v I__3243 (
            .O(N__15258),
            .I(N__15241));
    InMux I__3242 (
            .O(N__15257),
            .I(N__15236));
    InMux I__3241 (
            .O(N__15256),
            .I(N__15236));
    Sp12to4 I__3240 (
            .O(N__15249),
            .I(N__15227));
    Sp12to4 I__3239 (
            .O(N__15244),
            .I(N__15227));
    Sp12to4 I__3238 (
            .O(N__15241),
            .I(N__15227));
    LocalMux I__3237 (
            .O(N__15236),
            .I(N__15227));
    Odrv12 I__3236 (
            .O(N__15227),
            .I(M_this_reset_cond_out_0));
    CascadeMux I__3235 (
            .O(N__15224),
            .I(N__15221));
    CascadeBuf I__3234 (
            .O(N__15221),
            .I(N__15218));
    CascadeMux I__3233 (
            .O(N__15218),
            .I(N__15215));
    CascadeBuf I__3232 (
            .O(N__15215),
            .I(N__15212));
    CascadeMux I__3231 (
            .O(N__15212),
            .I(N__15209));
    CascadeBuf I__3230 (
            .O(N__15209),
            .I(N__15206));
    CascadeMux I__3229 (
            .O(N__15206),
            .I(N__15203));
    CascadeBuf I__3228 (
            .O(N__15203),
            .I(N__15200));
    CascadeMux I__3227 (
            .O(N__15200),
            .I(N__15197));
    CascadeBuf I__3226 (
            .O(N__15197),
            .I(N__15194));
    CascadeMux I__3225 (
            .O(N__15194),
            .I(N__15191));
    CascadeBuf I__3224 (
            .O(N__15191),
            .I(N__15188));
    CascadeMux I__3223 (
            .O(N__15188),
            .I(N__15185));
    CascadeBuf I__3222 (
            .O(N__15185),
            .I(N__15182));
    CascadeMux I__3221 (
            .O(N__15182),
            .I(N__15179));
    CascadeBuf I__3220 (
            .O(N__15179),
            .I(N__15176));
    CascadeMux I__3219 (
            .O(N__15176),
            .I(N__15173));
    CascadeBuf I__3218 (
            .O(N__15173),
            .I(N__15170));
    CascadeMux I__3217 (
            .O(N__15170),
            .I(N__15167));
    CascadeBuf I__3216 (
            .O(N__15167),
            .I(N__15164));
    CascadeMux I__3215 (
            .O(N__15164),
            .I(N__15161));
    CascadeBuf I__3214 (
            .O(N__15161),
            .I(N__15158));
    CascadeMux I__3213 (
            .O(N__15158),
            .I(N__15155));
    CascadeBuf I__3212 (
            .O(N__15155),
            .I(N__15152));
    CascadeMux I__3211 (
            .O(N__15152),
            .I(N__15149));
    CascadeBuf I__3210 (
            .O(N__15149),
            .I(N__15146));
    CascadeMux I__3209 (
            .O(N__15146),
            .I(N__15143));
    CascadeBuf I__3208 (
            .O(N__15143),
            .I(N__15140));
    CascadeMux I__3207 (
            .O(N__15140),
            .I(N__15137));
    CascadeBuf I__3206 (
            .O(N__15137),
            .I(N__15134));
    CascadeMux I__3205 (
            .O(N__15134),
            .I(N__15131));
    InMux I__3204 (
            .O(N__15131),
            .I(N__15128));
    LocalMux I__3203 (
            .O(N__15128),
            .I(N__15123));
    InMux I__3202 (
            .O(N__15127),
            .I(N__15120));
    InMux I__3201 (
            .O(N__15126),
            .I(N__15117));
    Span12Mux_s9_v I__3200 (
            .O(N__15123),
            .I(N__15114));
    LocalMux I__3199 (
            .O(N__15120),
            .I(M_current_address_qZ0Z_9));
    LocalMux I__3198 (
            .O(N__15117),
            .I(M_current_address_qZ0Z_9));
    Odrv12 I__3197 (
            .O(N__15114),
            .I(M_current_address_qZ0Z_9));
    CascadeMux I__3196 (
            .O(N__15107),
            .I(N__15104));
    InMux I__3195 (
            .O(N__15104),
            .I(N__15101));
    LocalMux I__3194 (
            .O(N__15101),
            .I(N_410));
    InMux I__3193 (
            .O(N__15098),
            .I(N__15095));
    LocalMux I__3192 (
            .O(N__15095),
            .I(N__15092));
    Odrv12 I__3191 (
            .O(N__15092),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    CascadeMux I__3190 (
            .O(N__15089),
            .I(N__15086));
    CascadeBuf I__3189 (
            .O(N__15086),
            .I(N__15083));
    CascadeMux I__3188 (
            .O(N__15083),
            .I(N__15080));
    CascadeBuf I__3187 (
            .O(N__15080),
            .I(N__15077));
    CascadeMux I__3186 (
            .O(N__15077),
            .I(N__15074));
    CascadeBuf I__3185 (
            .O(N__15074),
            .I(N__15071));
    CascadeMux I__3184 (
            .O(N__15071),
            .I(N__15068));
    CascadeBuf I__3183 (
            .O(N__15068),
            .I(N__15065));
    CascadeMux I__3182 (
            .O(N__15065),
            .I(N__15062));
    CascadeBuf I__3181 (
            .O(N__15062),
            .I(N__15059));
    CascadeMux I__3180 (
            .O(N__15059),
            .I(N__15056));
    CascadeBuf I__3179 (
            .O(N__15056),
            .I(N__15053));
    CascadeMux I__3178 (
            .O(N__15053),
            .I(N__15050));
    CascadeBuf I__3177 (
            .O(N__15050),
            .I(N__15047));
    CascadeMux I__3176 (
            .O(N__15047),
            .I(N__15044));
    CascadeBuf I__3175 (
            .O(N__15044),
            .I(N__15041));
    CascadeMux I__3174 (
            .O(N__15041),
            .I(N__15038));
    CascadeBuf I__3173 (
            .O(N__15038),
            .I(N__15035));
    CascadeMux I__3172 (
            .O(N__15035),
            .I(N__15032));
    CascadeBuf I__3171 (
            .O(N__15032),
            .I(N__15029));
    CascadeMux I__3170 (
            .O(N__15029),
            .I(N__15026));
    CascadeBuf I__3169 (
            .O(N__15026),
            .I(N__15023));
    CascadeMux I__3168 (
            .O(N__15023),
            .I(N__15020));
    CascadeBuf I__3167 (
            .O(N__15020),
            .I(N__15017));
    CascadeMux I__3166 (
            .O(N__15017),
            .I(N__15014));
    CascadeBuf I__3165 (
            .O(N__15014),
            .I(N__15011));
    CascadeMux I__3164 (
            .O(N__15011),
            .I(N__15008));
    CascadeBuf I__3163 (
            .O(N__15008),
            .I(N__15005));
    CascadeMux I__3162 (
            .O(N__15005),
            .I(N__15002));
    CascadeBuf I__3161 (
            .O(N__15002),
            .I(N__14999));
    CascadeMux I__3160 (
            .O(N__14999),
            .I(N__14996));
    InMux I__3159 (
            .O(N__14996),
            .I(N__14993));
    LocalMux I__3158 (
            .O(N__14993),
            .I(N__14990));
    Span4Mux_h I__3157 (
            .O(N__14990),
            .I(N__14987));
    Sp12to4 I__3156 (
            .O(N__14987),
            .I(N__14984));
    Span12Mux_s9_v I__3155 (
            .O(N__14984),
            .I(N__14981));
    Odrv12 I__3154 (
            .O(N__14981),
            .I(M_this_vga_signals_address_5));
    CascadeMux I__3153 (
            .O(N__14978),
            .I(N__14975));
    InMux I__3152 (
            .O(N__14975),
            .I(N__14972));
    LocalMux I__3151 (
            .O(N__14972),
            .I(N__14969));
    Span4Mux_h I__3150 (
            .O(N__14969),
            .I(N__14966));
    Odrv4 I__3149 (
            .O(N__14966),
            .I(mem_radreg_RNIETEJ4_11));
    InMux I__3148 (
            .O(N__14963),
            .I(N__14959));
    InMux I__3147 (
            .O(N__14962),
            .I(N__14956));
    LocalMux I__3146 (
            .O(N__14959),
            .I(m19));
    LocalMux I__3145 (
            .O(N__14956),
            .I(m19));
    InMux I__3144 (
            .O(N__14951),
            .I(N__14944));
    InMux I__3143 (
            .O(N__14950),
            .I(N__14939));
    InMux I__3142 (
            .O(N__14949),
            .I(N__14939));
    InMux I__3141 (
            .O(N__14948),
            .I(N__14931));
    InMux I__3140 (
            .O(N__14947),
            .I(N__14931));
    LocalMux I__3139 (
            .O(N__14944),
            .I(N__14926));
    LocalMux I__3138 (
            .O(N__14939),
            .I(N__14926));
    InMux I__3137 (
            .O(N__14938),
            .I(N__14923));
    InMux I__3136 (
            .O(N__14937),
            .I(N__14920));
    InMux I__3135 (
            .O(N__14936),
            .I(N__14917));
    LocalMux I__3134 (
            .O(N__14931),
            .I(rgb_1_axb_0));
    Odrv4 I__3133 (
            .O(N__14926),
            .I(rgb_1_axb_0));
    LocalMux I__3132 (
            .O(N__14923),
            .I(rgb_1_axb_0));
    LocalMux I__3131 (
            .O(N__14920),
            .I(rgb_1_axb_0));
    LocalMux I__3130 (
            .O(N__14917),
            .I(rgb_1_axb_0));
    InMux I__3129 (
            .O(N__14906),
            .I(N__14901));
    InMux I__3128 (
            .O(N__14905),
            .I(N__14898));
    InMux I__3127 (
            .O(N__14904),
            .I(N__14895));
    LocalMux I__3126 (
            .O(N__14901),
            .I(N__14892));
    LocalMux I__3125 (
            .O(N__14898),
            .I(N__14884));
    LocalMux I__3124 (
            .O(N__14895),
            .I(N__14884));
    Span4Mux_v I__3123 (
            .O(N__14892),
            .I(N__14881));
    InMux I__3122 (
            .O(N__14891),
            .I(N__14878));
    InMux I__3121 (
            .O(N__14890),
            .I(N__14875));
    InMux I__3120 (
            .O(N__14889),
            .I(N__14872));
    Odrv4 I__3119 (
            .O(N__14884),
            .I(a0_b_0));
    Odrv4 I__3118 (
            .O(N__14881),
            .I(a0_b_0));
    LocalMux I__3117 (
            .O(N__14878),
            .I(a0_b_0));
    LocalMux I__3116 (
            .O(N__14875),
            .I(a0_b_0));
    LocalMux I__3115 (
            .O(N__14872),
            .I(a0_b_0));
    CascadeMux I__3114 (
            .O(N__14861),
            .I(m46_am_cascade_));
    InMux I__3113 (
            .O(N__14858),
            .I(N__14855));
    LocalMux I__3112 (
            .O(N__14855),
            .I(N__14852));
    Odrv4 I__3111 (
            .O(N__14852),
            .I(m46_bm));
    CascadeMux I__3110 (
            .O(N__14849),
            .I(N__14846));
    InMux I__3109 (
            .O(N__14846),
            .I(N__14843));
    LocalMux I__3108 (
            .O(N__14843),
            .I(N__14840));
    Span12Mux_h I__3107 (
            .O(N__14840),
            .I(N__14837));
    Odrv12 I__3106 (
            .O(N__14837),
            .I(rgb_2_5));
    InMux I__3105 (
            .O(N__14834),
            .I(N__14831));
    LocalMux I__3104 (
            .O(N__14831),
            .I(N_352));
    CascadeMux I__3103 (
            .O(N__14828),
            .I(N_408_cascade_));
    InMux I__3102 (
            .O(N__14825),
            .I(N__14822));
    LocalMux I__3101 (
            .O(N__14822),
            .I(N__14819));
    Odrv4 I__3100 (
            .O(N__14819),
            .I(M_current_address_q_RNO_1Z0Z_7));
    CascadeMux I__3099 (
            .O(N__14816),
            .I(N__14813));
    CascadeBuf I__3098 (
            .O(N__14813),
            .I(N__14810));
    CascadeMux I__3097 (
            .O(N__14810),
            .I(N__14807));
    CascadeBuf I__3096 (
            .O(N__14807),
            .I(N__14804));
    CascadeMux I__3095 (
            .O(N__14804),
            .I(N__14801));
    CascadeBuf I__3094 (
            .O(N__14801),
            .I(N__14798));
    CascadeMux I__3093 (
            .O(N__14798),
            .I(N__14795));
    CascadeBuf I__3092 (
            .O(N__14795),
            .I(N__14792));
    CascadeMux I__3091 (
            .O(N__14792),
            .I(N__14789));
    CascadeBuf I__3090 (
            .O(N__14789),
            .I(N__14786));
    CascadeMux I__3089 (
            .O(N__14786),
            .I(N__14783));
    CascadeBuf I__3088 (
            .O(N__14783),
            .I(N__14780));
    CascadeMux I__3087 (
            .O(N__14780),
            .I(N__14777));
    CascadeBuf I__3086 (
            .O(N__14777),
            .I(N__14774));
    CascadeMux I__3085 (
            .O(N__14774),
            .I(N__14771));
    CascadeBuf I__3084 (
            .O(N__14771),
            .I(N__14768));
    CascadeMux I__3083 (
            .O(N__14768),
            .I(N__14765));
    CascadeBuf I__3082 (
            .O(N__14765),
            .I(N__14762));
    CascadeMux I__3081 (
            .O(N__14762),
            .I(N__14759));
    CascadeBuf I__3080 (
            .O(N__14759),
            .I(N__14756));
    CascadeMux I__3079 (
            .O(N__14756),
            .I(N__14753));
    CascadeBuf I__3078 (
            .O(N__14753),
            .I(N__14750));
    CascadeMux I__3077 (
            .O(N__14750),
            .I(N__14747));
    CascadeBuf I__3076 (
            .O(N__14747),
            .I(N__14744));
    CascadeMux I__3075 (
            .O(N__14744),
            .I(N__14741));
    CascadeBuf I__3074 (
            .O(N__14741),
            .I(N__14738));
    CascadeMux I__3073 (
            .O(N__14738),
            .I(N__14735));
    CascadeBuf I__3072 (
            .O(N__14735),
            .I(N__14732));
    CascadeMux I__3071 (
            .O(N__14732),
            .I(N__14729));
    CascadeBuf I__3070 (
            .O(N__14729),
            .I(N__14726));
    CascadeMux I__3069 (
            .O(N__14726),
            .I(N__14723));
    InMux I__3068 (
            .O(N__14723),
            .I(N__14720));
    LocalMux I__3067 (
            .O(N__14720),
            .I(N__14717));
    Span4Mux_h I__3066 (
            .O(N__14717),
            .I(N__14713));
    InMux I__3065 (
            .O(N__14716),
            .I(N__14709));
    Sp12to4 I__3064 (
            .O(N__14713),
            .I(N__14706));
    InMux I__3063 (
            .O(N__14712),
            .I(N__14703));
    LocalMux I__3062 (
            .O(N__14709),
            .I(N__14698));
    Span12Mux_s11_v I__3061 (
            .O(N__14706),
            .I(N__14698));
    LocalMux I__3060 (
            .O(N__14703),
            .I(M_current_address_qZ0Z_7));
    Odrv12 I__3059 (
            .O(N__14698),
            .I(M_current_address_qZ0Z_7));
    CascadeMux I__3058 (
            .O(N__14693),
            .I(N__14690));
    InMux I__3057 (
            .O(N__14690),
            .I(N__14687));
    LocalMux I__3056 (
            .O(N__14687),
            .I(N_405));
    InMux I__3055 (
            .O(N__14684),
            .I(N__14681));
    LocalMux I__3054 (
            .O(N__14681),
            .I(N__14678));
    Odrv4 I__3053 (
            .O(N__14678),
            .I(M_current_address_q_RNO_1Z0Z_4));
    CascadeMux I__3052 (
            .O(N__14675),
            .I(N__14672));
    CascadeBuf I__3051 (
            .O(N__14672),
            .I(N__14669));
    CascadeMux I__3050 (
            .O(N__14669),
            .I(N__14666));
    CascadeBuf I__3049 (
            .O(N__14666),
            .I(N__14663));
    CascadeMux I__3048 (
            .O(N__14663),
            .I(N__14660));
    CascadeBuf I__3047 (
            .O(N__14660),
            .I(N__14657));
    CascadeMux I__3046 (
            .O(N__14657),
            .I(N__14654));
    CascadeBuf I__3045 (
            .O(N__14654),
            .I(N__14651));
    CascadeMux I__3044 (
            .O(N__14651),
            .I(N__14648));
    CascadeBuf I__3043 (
            .O(N__14648),
            .I(N__14645));
    CascadeMux I__3042 (
            .O(N__14645),
            .I(N__14642));
    CascadeBuf I__3041 (
            .O(N__14642),
            .I(N__14639));
    CascadeMux I__3040 (
            .O(N__14639),
            .I(N__14636));
    CascadeBuf I__3039 (
            .O(N__14636),
            .I(N__14633));
    CascadeMux I__3038 (
            .O(N__14633),
            .I(N__14630));
    CascadeBuf I__3037 (
            .O(N__14630),
            .I(N__14627));
    CascadeMux I__3036 (
            .O(N__14627),
            .I(N__14624));
    CascadeBuf I__3035 (
            .O(N__14624),
            .I(N__14621));
    CascadeMux I__3034 (
            .O(N__14621),
            .I(N__14618));
    CascadeBuf I__3033 (
            .O(N__14618),
            .I(N__14615));
    CascadeMux I__3032 (
            .O(N__14615),
            .I(N__14612));
    CascadeBuf I__3031 (
            .O(N__14612),
            .I(N__14609));
    CascadeMux I__3030 (
            .O(N__14609),
            .I(N__14606));
    CascadeBuf I__3029 (
            .O(N__14606),
            .I(N__14603));
    CascadeMux I__3028 (
            .O(N__14603),
            .I(N__14600));
    CascadeBuf I__3027 (
            .O(N__14600),
            .I(N__14597));
    CascadeMux I__3026 (
            .O(N__14597),
            .I(N__14594));
    CascadeBuf I__3025 (
            .O(N__14594),
            .I(N__14591));
    CascadeMux I__3024 (
            .O(N__14591),
            .I(N__14588));
    CascadeBuf I__3023 (
            .O(N__14588),
            .I(N__14585));
    CascadeMux I__3022 (
            .O(N__14585),
            .I(N__14582));
    InMux I__3021 (
            .O(N__14582),
            .I(N__14579));
    LocalMux I__3020 (
            .O(N__14579),
            .I(N__14576));
    Span4Mux_s1_v I__3019 (
            .O(N__14576),
            .I(N__14572));
    InMux I__3018 (
            .O(N__14575),
            .I(N__14569));
    Sp12to4 I__3017 (
            .O(N__14572),
            .I(N__14565));
    LocalMux I__3016 (
            .O(N__14569),
            .I(N__14562));
    InMux I__3015 (
            .O(N__14568),
            .I(N__14559));
    Span12Mux_h I__3014 (
            .O(N__14565),
            .I(N__14556));
    Odrv4 I__3013 (
            .O(N__14562),
            .I(M_current_address_qZ0Z_4));
    LocalMux I__3012 (
            .O(N__14559),
            .I(M_current_address_qZ0Z_4));
    Odrv12 I__3011 (
            .O(N__14556),
            .I(M_current_address_qZ0Z_4));
    CascadeMux I__3010 (
            .O(N__14549),
            .I(N__14546));
    InMux I__3009 (
            .O(N__14546),
            .I(N__14542));
    InMux I__3008 (
            .O(N__14545),
            .I(N__14539));
    LocalMux I__3007 (
            .O(N__14542),
            .I(N__14536));
    LocalMux I__3006 (
            .O(N__14539),
            .I(N__14533));
    Span4Mux_h I__3005 (
            .O(N__14536),
            .I(N__14530));
    Span4Mux_h I__3004 (
            .O(N__14533),
            .I(N__14527));
    Odrv4 I__3003 (
            .O(N__14530),
            .I(M_state_q_ns_0_a3_0_2_0));
    Odrv4 I__3002 (
            .O(N__14527),
            .I(M_state_q_ns_0_a3_0_2_0));
    CascadeMux I__3001 (
            .O(N__14522),
            .I(N__14519));
    InMux I__3000 (
            .O(N__14519),
            .I(N__14516));
    LocalMux I__2999 (
            .O(N__14516),
            .I(N_351));
    InMux I__2998 (
            .O(N__14513),
            .I(N__14509));
    InMux I__2997 (
            .O(N__14512),
            .I(N__14506));
    LocalMux I__2996 (
            .O(N__14509),
            .I(m24));
    LocalMux I__2995 (
            .O(N__14506),
            .I(m24));
    CascadeMux I__2994 (
            .O(N__14501),
            .I(m40_cascade_));
    InMux I__2993 (
            .O(N__14498),
            .I(N__14495));
    LocalMux I__2992 (
            .O(N__14495),
            .I(m41));
    InMux I__2991 (
            .O(N__14492),
            .I(N__14486));
    InMux I__2990 (
            .O(N__14491),
            .I(N__14486));
    LocalMux I__2989 (
            .O(N__14486),
            .I(m10));
    CascadeMux I__2988 (
            .O(N__14483),
            .I(rgb_1_axb_0_cascade_));
    InMux I__2987 (
            .O(N__14480),
            .I(N__14474));
    InMux I__2986 (
            .O(N__14479),
            .I(N__14474));
    LocalMux I__2985 (
            .O(N__14474),
            .I(N__14471));
    Span4Mux_v I__2984 (
            .O(N__14471),
            .I(N__14468));
    Odrv4 I__2983 (
            .O(N__14468),
            .I(m15));
    InMux I__2982 (
            .O(N__14465),
            .I(N__14462));
    LocalMux I__2981 (
            .O(N__14462),
            .I(N__14458));
    InMux I__2980 (
            .O(N__14461),
            .I(N__14455));
    Span4Mux_v I__2979 (
            .O(N__14458),
            .I(N__14450));
    LocalMux I__2978 (
            .O(N__14455),
            .I(N__14450));
    Odrv4 I__2977 (
            .O(N__14450),
            .I(rgb_1_0));
    InMux I__2976 (
            .O(N__14447),
            .I(N__14444));
    LocalMux I__2975 (
            .O(N__14444),
            .I(m37));
    SRMux I__2974 (
            .O(N__14441),
            .I(N__14437));
    SRMux I__2973 (
            .O(N__14440),
            .I(N__14431));
    LocalMux I__2972 (
            .O(N__14437),
            .I(N__14427));
    SRMux I__2971 (
            .O(N__14436),
            .I(N__14423));
    SRMux I__2970 (
            .O(N__14435),
            .I(N__14420));
    SRMux I__2969 (
            .O(N__14434),
            .I(N__14415));
    LocalMux I__2968 (
            .O(N__14431),
            .I(N__14409));
    SRMux I__2967 (
            .O(N__14430),
            .I(N__14406));
    Span4Mux_s3_v I__2966 (
            .O(N__14427),
            .I(N__14403));
    SRMux I__2965 (
            .O(N__14426),
            .I(N__14400));
    LocalMux I__2964 (
            .O(N__14423),
            .I(N__14393));
    LocalMux I__2963 (
            .O(N__14420),
            .I(N__14393));
    SRMux I__2962 (
            .O(N__14419),
            .I(N__14390));
    SRMux I__2961 (
            .O(N__14418),
            .I(N__14382));
    LocalMux I__2960 (
            .O(N__14415),
            .I(N__14379));
    SRMux I__2959 (
            .O(N__14414),
            .I(N__14376));
    SRMux I__2958 (
            .O(N__14413),
            .I(N__14373));
    SRMux I__2957 (
            .O(N__14412),
            .I(N__14370));
    Span4Mux_h I__2956 (
            .O(N__14409),
            .I(N__14363));
    LocalMux I__2955 (
            .O(N__14406),
            .I(N__14363));
    Span4Mux_v I__2954 (
            .O(N__14403),
            .I(N__14358));
    LocalMux I__2953 (
            .O(N__14400),
            .I(N__14358));
    SRMux I__2952 (
            .O(N__14399),
            .I(N__14355));
    SRMux I__2951 (
            .O(N__14398),
            .I(N__14352));
    Span4Mux_s3_v I__2950 (
            .O(N__14393),
            .I(N__14346));
    LocalMux I__2949 (
            .O(N__14390),
            .I(N__14346));
    SRMux I__2948 (
            .O(N__14389),
            .I(N__14343));
    SRMux I__2947 (
            .O(N__14388),
            .I(N__14340));
    IoInMux I__2946 (
            .O(N__14387),
            .I(N__14334));
    SRMux I__2945 (
            .O(N__14386),
            .I(N__14331));
    SRMux I__2944 (
            .O(N__14385),
            .I(N__14328));
    LocalMux I__2943 (
            .O(N__14382),
            .I(N__14320));
    Span4Mux_h I__2942 (
            .O(N__14379),
            .I(N__14320));
    LocalMux I__2941 (
            .O(N__14376),
            .I(N__14320));
    LocalMux I__2940 (
            .O(N__14373),
            .I(N__14315));
    LocalMux I__2939 (
            .O(N__14370),
            .I(N__14315));
    SRMux I__2938 (
            .O(N__14369),
            .I(N__14312));
    SRMux I__2937 (
            .O(N__14368),
            .I(N__14308));
    Span4Mux_v I__2936 (
            .O(N__14363),
            .I(N__14298));
    Span4Mux_h I__2935 (
            .O(N__14358),
            .I(N__14298));
    LocalMux I__2934 (
            .O(N__14355),
            .I(N__14298));
    LocalMux I__2933 (
            .O(N__14352),
            .I(N__14295));
    SRMux I__2932 (
            .O(N__14351),
            .I(N__14292));
    Span4Mux_v I__2931 (
            .O(N__14346),
            .I(N__14285));
    LocalMux I__2930 (
            .O(N__14343),
            .I(N__14285));
    LocalMux I__2929 (
            .O(N__14340),
            .I(N__14285));
    SRMux I__2928 (
            .O(N__14339),
            .I(N__14282));
    SRMux I__2927 (
            .O(N__14338),
            .I(N__14279));
    InMux I__2926 (
            .O(N__14337),
            .I(N__14275));
    LocalMux I__2925 (
            .O(N__14334),
            .I(N__14272));
    LocalMux I__2924 (
            .O(N__14331),
            .I(N__14266));
    LocalMux I__2923 (
            .O(N__14328),
            .I(N__14266));
    SRMux I__2922 (
            .O(N__14327),
            .I(N__14263));
    Span4Mux_v I__2921 (
            .O(N__14320),
            .I(N__14256));
    Span4Mux_v I__2920 (
            .O(N__14315),
            .I(N__14256));
    LocalMux I__2919 (
            .O(N__14312),
            .I(N__14256));
    SRMux I__2918 (
            .O(N__14311),
            .I(N__14253));
    LocalMux I__2917 (
            .O(N__14308),
            .I(N__14250));
    SRMux I__2916 (
            .O(N__14307),
            .I(N__14247));
    SRMux I__2915 (
            .O(N__14306),
            .I(N__14244));
    SRMux I__2914 (
            .O(N__14305),
            .I(N__14241));
    Span4Mux_v I__2913 (
            .O(N__14298),
            .I(N__14234));
    Span4Mux_h I__2912 (
            .O(N__14295),
            .I(N__14234));
    LocalMux I__2911 (
            .O(N__14292),
            .I(N__14234));
    Span4Mux_v I__2910 (
            .O(N__14285),
            .I(N__14227));
    LocalMux I__2909 (
            .O(N__14282),
            .I(N__14227));
    LocalMux I__2908 (
            .O(N__14279),
            .I(N__14227));
    SRMux I__2907 (
            .O(N__14278),
            .I(N__14224));
    LocalMux I__2906 (
            .O(N__14275),
            .I(N__14220));
    Span4Mux_s2_h I__2905 (
            .O(N__14272),
            .I(N__14217));
    SRMux I__2904 (
            .O(N__14271),
            .I(N__14214));
    Span4Mux_v I__2903 (
            .O(N__14266),
            .I(N__14209));
    LocalMux I__2902 (
            .O(N__14263),
            .I(N__14209));
    Span4Mux_v I__2901 (
            .O(N__14256),
            .I(N__14204));
    LocalMux I__2900 (
            .O(N__14253),
            .I(N__14204));
    Span4Mux_h I__2899 (
            .O(N__14250),
            .I(N__14199));
    LocalMux I__2898 (
            .O(N__14247),
            .I(N__14199));
    LocalMux I__2897 (
            .O(N__14244),
            .I(N__14194));
    LocalMux I__2896 (
            .O(N__14241),
            .I(N__14194));
    Span4Mux_v I__2895 (
            .O(N__14234),
            .I(N__14187));
    Span4Mux_v I__2894 (
            .O(N__14227),
            .I(N__14187));
    LocalMux I__2893 (
            .O(N__14224),
            .I(N__14187));
    SRMux I__2892 (
            .O(N__14223),
            .I(N__14184));
    Span4Mux_h I__2891 (
            .O(N__14220),
            .I(N__14179));
    Sp12to4 I__2890 (
            .O(N__14217),
            .I(N__14176));
    LocalMux I__2889 (
            .O(N__14214),
            .I(N__14173));
    Span4Mux_h I__2888 (
            .O(N__14209),
            .I(N__14169));
    Span4Mux_v I__2887 (
            .O(N__14204),
            .I(N__14164));
    Span4Mux_v I__2886 (
            .O(N__14199),
            .I(N__14164));
    Span4Mux_v I__2885 (
            .O(N__14194),
            .I(N__14157));
    Span4Mux_v I__2884 (
            .O(N__14187),
            .I(N__14157));
    LocalMux I__2883 (
            .O(N__14184),
            .I(N__14157));
    CascadeMux I__2882 (
            .O(N__14183),
            .I(N__14154));
    CascadeMux I__2881 (
            .O(N__14182),
            .I(N__14151));
    Span4Mux_v I__2880 (
            .O(N__14179),
            .I(N__14147));
    Span12Mux_v I__2879 (
            .O(N__14176),
            .I(N__14144));
    Span12Mux_h I__2878 (
            .O(N__14173),
            .I(N__14141));
    SRMux I__2877 (
            .O(N__14172),
            .I(N__14138));
    Span4Mux_v I__2876 (
            .O(N__14169),
            .I(N__14131));
    Span4Mux_h I__2875 (
            .O(N__14164),
            .I(N__14131));
    Span4Mux_h I__2874 (
            .O(N__14157),
            .I(N__14131));
    InMux I__2873 (
            .O(N__14154),
            .I(N__14128));
    InMux I__2872 (
            .O(N__14151),
            .I(N__14123));
    InMux I__2871 (
            .O(N__14150),
            .I(N__14123));
    Span4Mux_v I__2870 (
            .O(N__14147),
            .I(N__14120));
    Span12Mux_h I__2869 (
            .O(N__14144),
            .I(N__14113));
    Span12Mux_v I__2868 (
            .O(N__14141),
            .I(N__14113));
    LocalMux I__2867 (
            .O(N__14138),
            .I(N__14113));
    Span4Mux_h I__2866 (
            .O(N__14131),
            .I(N__14110));
    LocalMux I__2865 (
            .O(N__14128),
            .I(N__14105));
    LocalMux I__2864 (
            .O(N__14123),
            .I(N__14105));
    Odrv4 I__2863 (
            .O(N__14120),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__2862 (
            .O(N__14113),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2861 (
            .O(N__14110),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2860 (
            .O(N__14105),
            .I(CONSTANT_ONE_NET));
    InMux I__2859 (
            .O(N__14096),
            .I(rgb291));
    InMux I__2858 (
            .O(N__14093),
            .I(N__14085));
    InMux I__2857 (
            .O(N__14092),
            .I(N__14085));
    InMux I__2856 (
            .O(N__14091),
            .I(N__14081));
    InMux I__2855 (
            .O(N__14090),
            .I(N__14078));
    LocalMux I__2854 (
            .O(N__14085),
            .I(N__14074));
    InMux I__2853 (
            .O(N__14084),
            .I(N__14071));
    LocalMux I__2852 (
            .O(N__14081),
            .I(N__14068));
    LocalMux I__2851 (
            .O(N__14078),
            .I(N__14065));
    InMux I__2850 (
            .O(N__14077),
            .I(N__14062));
    Span4Mux_h I__2849 (
            .O(N__14074),
            .I(N__14057));
    LocalMux I__2848 (
            .O(N__14071),
            .I(N__14057));
    Span4Mux_v I__2847 (
            .O(N__14068),
            .I(N__14054));
    Span4Mux_v I__2846 (
            .O(N__14065),
            .I(N__14049));
    LocalMux I__2845 (
            .O(N__14062),
            .I(N__14049));
    Span4Mux_v I__2844 (
            .O(N__14057),
            .I(N__14046));
    Sp12to4 I__2843 (
            .O(N__14054),
            .I(N__14043));
    Span4Mux_v I__2842 (
            .O(N__14049),
            .I(N__14040));
    Sp12to4 I__2841 (
            .O(N__14046),
            .I(N__14037));
    Span12Mux_h I__2840 (
            .O(N__14043),
            .I(N__14034));
    Span4Mux_h I__2839 (
            .O(N__14040),
            .I(N__14031));
    Odrv12 I__2838 (
            .O(N__14037),
            .I(\this_vga_signals.rgb_1_sqmuxa ));
    Odrv12 I__2837 (
            .O(N__14034),
            .I(\this_vga_signals.rgb_1_sqmuxa ));
    Odrv4 I__2836 (
            .O(N__14031),
            .I(\this_vga_signals.rgb_1_sqmuxa ));
    InMux I__2835 (
            .O(N__14024),
            .I(N__14021));
    LocalMux I__2834 (
            .O(N__14021),
            .I(mem_radreg_RNIMTEJ4_0_11));
    InMux I__2833 (
            .O(N__14018),
            .I(N__14015));
    LocalMux I__2832 (
            .O(N__14015),
            .I(mem_radreg_RNIETEJ4_0_11));
    CascadeMux I__2831 (
            .O(N__14012),
            .I(m44_cascade_));
    CascadeMux I__2830 (
            .O(N__14009),
            .I(m22_am_cascade_));
    InMux I__2829 (
            .O(N__14006),
            .I(N__14003));
    LocalMux I__2828 (
            .O(N__14003),
            .I(N__14000));
    Odrv4 I__2827 (
            .O(N__14000),
            .I(m22_ns));
    InMux I__2826 (
            .O(N__13997),
            .I(N__13994));
    LocalMux I__2825 (
            .O(N__13994),
            .I(m22_bm));
    InMux I__2824 (
            .O(N__13991),
            .I(N__13988));
    LocalMux I__2823 (
            .O(N__13988),
            .I(M_current_address_q_RNO_1Z0Z_8));
    InMux I__2822 (
            .O(N__13985),
            .I(N__13982));
    LocalMux I__2821 (
            .O(N__13982),
            .I(N__13979));
    Span4Mux_h I__2820 (
            .O(N__13979),
            .I(N__13976));
    Odrv4 I__2819 (
            .O(N__13976),
            .I(N_409));
    CascadeMux I__2818 (
            .O(N__13973),
            .I(N__13970));
    CascadeBuf I__2817 (
            .O(N__13970),
            .I(N__13967));
    CascadeMux I__2816 (
            .O(N__13967),
            .I(N__13964));
    CascadeBuf I__2815 (
            .O(N__13964),
            .I(N__13961));
    CascadeMux I__2814 (
            .O(N__13961),
            .I(N__13958));
    CascadeBuf I__2813 (
            .O(N__13958),
            .I(N__13955));
    CascadeMux I__2812 (
            .O(N__13955),
            .I(N__13952));
    CascadeBuf I__2811 (
            .O(N__13952),
            .I(N__13949));
    CascadeMux I__2810 (
            .O(N__13949),
            .I(N__13946));
    CascadeBuf I__2809 (
            .O(N__13946),
            .I(N__13943));
    CascadeMux I__2808 (
            .O(N__13943),
            .I(N__13940));
    CascadeBuf I__2807 (
            .O(N__13940),
            .I(N__13937));
    CascadeMux I__2806 (
            .O(N__13937),
            .I(N__13934));
    CascadeBuf I__2805 (
            .O(N__13934),
            .I(N__13931));
    CascadeMux I__2804 (
            .O(N__13931),
            .I(N__13928));
    CascadeBuf I__2803 (
            .O(N__13928),
            .I(N__13925));
    CascadeMux I__2802 (
            .O(N__13925),
            .I(N__13922));
    CascadeBuf I__2801 (
            .O(N__13922),
            .I(N__13919));
    CascadeMux I__2800 (
            .O(N__13919),
            .I(N__13916));
    CascadeBuf I__2799 (
            .O(N__13916),
            .I(N__13913));
    CascadeMux I__2798 (
            .O(N__13913),
            .I(N__13910));
    CascadeBuf I__2797 (
            .O(N__13910),
            .I(N__13907));
    CascadeMux I__2796 (
            .O(N__13907),
            .I(N__13904));
    CascadeBuf I__2795 (
            .O(N__13904),
            .I(N__13901));
    CascadeMux I__2794 (
            .O(N__13901),
            .I(N__13898));
    CascadeBuf I__2793 (
            .O(N__13898),
            .I(N__13895));
    CascadeMux I__2792 (
            .O(N__13895),
            .I(N__13892));
    CascadeBuf I__2791 (
            .O(N__13892),
            .I(N__13889));
    CascadeMux I__2790 (
            .O(N__13889),
            .I(N__13886));
    CascadeBuf I__2789 (
            .O(N__13886),
            .I(N__13883));
    CascadeMux I__2788 (
            .O(N__13883),
            .I(N__13880));
    InMux I__2787 (
            .O(N__13880),
            .I(N__13877));
    LocalMux I__2786 (
            .O(N__13877),
            .I(N__13874));
    Span4Mux_s3_v I__2785 (
            .O(N__13874),
            .I(N__13871));
    Span4Mux_h I__2784 (
            .O(N__13871),
            .I(N__13867));
    InMux I__2783 (
            .O(N__13870),
            .I(N__13863));
    Span4Mux_h I__2782 (
            .O(N__13867),
            .I(N__13860));
    InMux I__2781 (
            .O(N__13866),
            .I(N__13857));
    LocalMux I__2780 (
            .O(N__13863),
            .I(N__13854));
    Span4Mux_v I__2779 (
            .O(N__13860),
            .I(N__13851));
    LocalMux I__2778 (
            .O(N__13857),
            .I(M_current_address_qZ0Z_8));
    Odrv4 I__2777 (
            .O(N__13854),
            .I(M_current_address_qZ0Z_8));
    Odrv4 I__2776 (
            .O(N__13851),
            .I(M_current_address_qZ0Z_8));
    InMux I__2775 (
            .O(N__13844),
            .I(N__13841));
    LocalMux I__2774 (
            .O(N__13841),
            .I(N__13838));
    Odrv12 I__2773 (
            .O(N__13838),
            .I(N_412));
    InMux I__2772 (
            .O(N__13835),
            .I(N__13832));
    LocalMux I__2771 (
            .O(N__13832),
            .I(M_current_address_q_RNO_1Z0Z_11));
    CascadeMux I__2770 (
            .O(N__13829),
            .I(N__13825));
    InMux I__2769 (
            .O(N__13828),
            .I(N__13822));
    InMux I__2768 (
            .O(N__13825),
            .I(N__13819));
    LocalMux I__2767 (
            .O(N__13822),
            .I(N__13814));
    LocalMux I__2766 (
            .O(N__13819),
            .I(N__13814));
    Span4Mux_v I__2765 (
            .O(N__13814),
            .I(N__13811));
    Span4Mux_v I__2764 (
            .O(N__13811),
            .I(N__13808));
    Sp12to4 I__2763 (
            .O(N__13808),
            .I(N__13805));
    Span12Mux_h I__2762 (
            .O(N__13805),
            .I(N__13802));
    Odrv12 I__2761 (
            .O(N__13802),
            .I(port_data_c_4));
    InMux I__2760 (
            .O(N__13799),
            .I(N__13796));
    LocalMux I__2759 (
            .O(N__13796),
            .I(M_current_address_q_RNO_1Z0Z_9));
    CascadeMux I__2758 (
            .O(N__13793),
            .I(N__13789));
    CascadeMux I__2757 (
            .O(N__13792),
            .I(N__13784));
    InMux I__2756 (
            .O(N__13789),
            .I(N__13779));
    InMux I__2755 (
            .O(N__13788),
            .I(N__13779));
    CascadeMux I__2754 (
            .O(N__13787),
            .I(N__13776));
    InMux I__2753 (
            .O(N__13784),
            .I(N__13771));
    LocalMux I__2752 (
            .O(N__13779),
            .I(N__13766));
    InMux I__2751 (
            .O(N__13776),
            .I(N__13761));
    InMux I__2750 (
            .O(N__13775),
            .I(N__13761));
    InMux I__2749 (
            .O(N__13774),
            .I(N__13758));
    LocalMux I__2748 (
            .O(N__13771),
            .I(N__13755));
    CascadeMux I__2747 (
            .O(N__13770),
            .I(N__13752));
    CascadeMux I__2746 (
            .O(N__13769),
            .I(N__13747));
    Span4Mux_v I__2745 (
            .O(N__13766),
            .I(N__13742));
    LocalMux I__2744 (
            .O(N__13761),
            .I(N__13742));
    LocalMux I__2743 (
            .O(N__13758),
            .I(N__13739));
    Span4Mux_v I__2742 (
            .O(N__13755),
            .I(N__13736));
    InMux I__2741 (
            .O(N__13752),
            .I(N__13731));
    InMux I__2740 (
            .O(N__13751),
            .I(N__13731));
    InMux I__2739 (
            .O(N__13750),
            .I(N__13726));
    InMux I__2738 (
            .O(N__13747),
            .I(N__13726));
    Span4Mux_v I__2737 (
            .O(N__13742),
            .I(N__13721));
    Span4Mux_v I__2736 (
            .O(N__13739),
            .I(N__13721));
    Span4Mux_h I__2735 (
            .O(N__13736),
            .I(N__13714));
    LocalMux I__2734 (
            .O(N__13731),
            .I(N__13714));
    LocalMux I__2733 (
            .O(N__13726),
            .I(N__13714));
    Span4Mux_h I__2732 (
            .O(N__13721),
            .I(N__13711));
    Span4Mux_v I__2731 (
            .O(N__13714),
            .I(N__13708));
    Span4Mux_h I__2730 (
            .O(N__13711),
            .I(N__13705));
    Span4Mux_h I__2729 (
            .O(N__13708),
            .I(N__13702));
    Odrv4 I__2728 (
            .O(N__13705),
            .I(M_this_vram_read_data_1));
    Odrv4 I__2727 (
            .O(N__13702),
            .I(M_this_vram_read_data_1));
    CascadeMux I__2726 (
            .O(N__13697),
            .I(N__13693));
    CascadeMux I__2725 (
            .O(N__13696),
            .I(N__13690));
    InMux I__2724 (
            .O(N__13693),
            .I(N__13687));
    InMux I__2723 (
            .O(N__13690),
            .I(N__13684));
    LocalMux I__2722 (
            .O(N__13687),
            .I(N__13681));
    LocalMux I__2721 (
            .O(N__13684),
            .I(N__13678));
    Span4Mux_v I__2720 (
            .O(N__13681),
            .I(N__13673));
    Span4Mux_v I__2719 (
            .O(N__13678),
            .I(N__13673));
    Sp12to4 I__2718 (
            .O(N__13673),
            .I(N__13670));
    Span12Mux_h I__2717 (
            .O(N__13670),
            .I(N__13667));
    Odrv12 I__2716 (
            .O(N__13667),
            .I(port_data_c_5));
    CascadeMux I__2715 (
            .O(N__13664),
            .I(N_413_cascade_));
    InMux I__2714 (
            .O(N__13661),
            .I(N__13658));
    LocalMux I__2713 (
            .O(N__13658),
            .I(M_current_address_q_RNO_1Z0Z_12));
    CascadeMux I__2712 (
            .O(N__13655),
            .I(N__13652));
    InMux I__2711 (
            .O(N__13652),
            .I(N__13649));
    LocalMux I__2710 (
            .O(N__13649),
            .I(N_411));
    InMux I__2709 (
            .O(N__13646),
            .I(N__13643));
    LocalMux I__2708 (
            .O(N__13643),
            .I(M_current_address_q_RNO_1Z0Z_10));
    CascadeMux I__2707 (
            .O(N__13640),
            .I(N__13637));
    CascadeBuf I__2706 (
            .O(N__13637),
            .I(N__13634));
    CascadeMux I__2705 (
            .O(N__13634),
            .I(N__13631));
    CascadeBuf I__2704 (
            .O(N__13631),
            .I(N__13628));
    CascadeMux I__2703 (
            .O(N__13628),
            .I(N__13625));
    CascadeBuf I__2702 (
            .O(N__13625),
            .I(N__13622));
    CascadeMux I__2701 (
            .O(N__13622),
            .I(N__13619));
    CascadeBuf I__2700 (
            .O(N__13619),
            .I(N__13616));
    CascadeMux I__2699 (
            .O(N__13616),
            .I(N__13613));
    CascadeBuf I__2698 (
            .O(N__13613),
            .I(N__13610));
    CascadeMux I__2697 (
            .O(N__13610),
            .I(N__13607));
    CascadeBuf I__2696 (
            .O(N__13607),
            .I(N__13604));
    CascadeMux I__2695 (
            .O(N__13604),
            .I(N__13601));
    CascadeBuf I__2694 (
            .O(N__13601),
            .I(N__13598));
    CascadeMux I__2693 (
            .O(N__13598),
            .I(N__13595));
    CascadeBuf I__2692 (
            .O(N__13595),
            .I(N__13592));
    CascadeMux I__2691 (
            .O(N__13592),
            .I(N__13589));
    CascadeBuf I__2690 (
            .O(N__13589),
            .I(N__13586));
    CascadeMux I__2689 (
            .O(N__13586),
            .I(N__13583));
    CascadeBuf I__2688 (
            .O(N__13583),
            .I(N__13580));
    CascadeMux I__2687 (
            .O(N__13580),
            .I(N__13577));
    CascadeBuf I__2686 (
            .O(N__13577),
            .I(N__13574));
    CascadeMux I__2685 (
            .O(N__13574),
            .I(N__13571));
    CascadeBuf I__2684 (
            .O(N__13571),
            .I(N__13568));
    CascadeMux I__2683 (
            .O(N__13568),
            .I(N__13565));
    CascadeBuf I__2682 (
            .O(N__13565),
            .I(N__13562));
    CascadeMux I__2681 (
            .O(N__13562),
            .I(N__13559));
    CascadeBuf I__2680 (
            .O(N__13559),
            .I(N__13556));
    CascadeMux I__2679 (
            .O(N__13556),
            .I(N__13553));
    CascadeBuf I__2678 (
            .O(N__13553),
            .I(N__13550));
    CascadeMux I__2677 (
            .O(N__13550),
            .I(N__13547));
    InMux I__2676 (
            .O(N__13547),
            .I(N__13544));
    LocalMux I__2675 (
            .O(N__13544),
            .I(N__13539));
    InMux I__2674 (
            .O(N__13543),
            .I(N__13536));
    InMux I__2673 (
            .O(N__13542),
            .I(N__13533));
    Span12Mux_h I__2672 (
            .O(N__13539),
            .I(N__13530));
    LocalMux I__2671 (
            .O(N__13536),
            .I(M_current_address_qZ0Z_10));
    LocalMux I__2670 (
            .O(N__13533),
            .I(M_current_address_qZ0Z_10));
    Odrv12 I__2669 (
            .O(N__13530),
            .I(M_current_address_qZ0Z_10));
    CascadeMux I__2668 (
            .O(N__13523),
            .I(N__13520));
    InMux I__2667 (
            .O(N__13520),
            .I(N__13517));
    LocalMux I__2666 (
            .O(N__13517),
            .I(N_404));
    InMux I__2665 (
            .O(N__13514),
            .I(N__13511));
    LocalMux I__2664 (
            .O(N__13511),
            .I(M_current_address_q_RNO_1Z0Z_3));
    CascadeMux I__2663 (
            .O(N__13508),
            .I(N__13505));
    CascadeBuf I__2662 (
            .O(N__13505),
            .I(N__13502));
    CascadeMux I__2661 (
            .O(N__13502),
            .I(N__13499));
    CascadeBuf I__2660 (
            .O(N__13499),
            .I(N__13496));
    CascadeMux I__2659 (
            .O(N__13496),
            .I(N__13493));
    CascadeBuf I__2658 (
            .O(N__13493),
            .I(N__13490));
    CascadeMux I__2657 (
            .O(N__13490),
            .I(N__13487));
    CascadeBuf I__2656 (
            .O(N__13487),
            .I(N__13484));
    CascadeMux I__2655 (
            .O(N__13484),
            .I(N__13481));
    CascadeBuf I__2654 (
            .O(N__13481),
            .I(N__13478));
    CascadeMux I__2653 (
            .O(N__13478),
            .I(N__13475));
    CascadeBuf I__2652 (
            .O(N__13475),
            .I(N__13472));
    CascadeMux I__2651 (
            .O(N__13472),
            .I(N__13469));
    CascadeBuf I__2650 (
            .O(N__13469),
            .I(N__13466));
    CascadeMux I__2649 (
            .O(N__13466),
            .I(N__13463));
    CascadeBuf I__2648 (
            .O(N__13463),
            .I(N__13460));
    CascadeMux I__2647 (
            .O(N__13460),
            .I(N__13457));
    CascadeBuf I__2646 (
            .O(N__13457),
            .I(N__13454));
    CascadeMux I__2645 (
            .O(N__13454),
            .I(N__13451));
    CascadeBuf I__2644 (
            .O(N__13451),
            .I(N__13448));
    CascadeMux I__2643 (
            .O(N__13448),
            .I(N__13445));
    CascadeBuf I__2642 (
            .O(N__13445),
            .I(N__13442));
    CascadeMux I__2641 (
            .O(N__13442),
            .I(N__13439));
    CascadeBuf I__2640 (
            .O(N__13439),
            .I(N__13436));
    CascadeMux I__2639 (
            .O(N__13436),
            .I(N__13433));
    CascadeBuf I__2638 (
            .O(N__13433),
            .I(N__13430));
    CascadeMux I__2637 (
            .O(N__13430),
            .I(N__13427));
    CascadeBuf I__2636 (
            .O(N__13427),
            .I(N__13424));
    CascadeMux I__2635 (
            .O(N__13424),
            .I(N__13421));
    CascadeBuf I__2634 (
            .O(N__13421),
            .I(N__13418));
    CascadeMux I__2633 (
            .O(N__13418),
            .I(N__13415));
    InMux I__2632 (
            .O(N__13415),
            .I(N__13412));
    LocalMux I__2631 (
            .O(N__13412),
            .I(N__13409));
    Span4Mux_h I__2630 (
            .O(N__13409),
            .I(N__13404));
    CascadeMux I__2629 (
            .O(N__13408),
            .I(N__13401));
    InMux I__2628 (
            .O(N__13407),
            .I(N__13398));
    Sp12to4 I__2627 (
            .O(N__13404),
            .I(N__13395));
    InMux I__2626 (
            .O(N__13401),
            .I(N__13392));
    LocalMux I__2625 (
            .O(N__13398),
            .I(N__13387));
    Span12Mux_s11_v I__2624 (
            .O(N__13395),
            .I(N__13387));
    LocalMux I__2623 (
            .O(N__13392),
            .I(M_current_address_qZ0Z_3));
    Odrv12 I__2622 (
            .O(N__13387),
            .I(M_current_address_qZ0Z_3));
    InMux I__2621 (
            .O(N__13382),
            .I(N__13379));
    LocalMux I__2620 (
            .O(N__13379),
            .I(M_current_address_q_RNO_1Z0Z_5));
    CascadeMux I__2619 (
            .O(N__13376),
            .I(N__13373));
    InMux I__2618 (
            .O(N__13373),
            .I(N__13370));
    LocalMux I__2617 (
            .O(N__13370),
            .I(N_406));
    CascadeMux I__2616 (
            .O(N__13367),
            .I(N__13364));
    CascadeBuf I__2615 (
            .O(N__13364),
            .I(N__13361));
    CascadeMux I__2614 (
            .O(N__13361),
            .I(N__13358));
    CascadeBuf I__2613 (
            .O(N__13358),
            .I(N__13355));
    CascadeMux I__2612 (
            .O(N__13355),
            .I(N__13352));
    CascadeBuf I__2611 (
            .O(N__13352),
            .I(N__13349));
    CascadeMux I__2610 (
            .O(N__13349),
            .I(N__13346));
    CascadeBuf I__2609 (
            .O(N__13346),
            .I(N__13343));
    CascadeMux I__2608 (
            .O(N__13343),
            .I(N__13340));
    CascadeBuf I__2607 (
            .O(N__13340),
            .I(N__13337));
    CascadeMux I__2606 (
            .O(N__13337),
            .I(N__13334));
    CascadeBuf I__2605 (
            .O(N__13334),
            .I(N__13331));
    CascadeMux I__2604 (
            .O(N__13331),
            .I(N__13328));
    CascadeBuf I__2603 (
            .O(N__13328),
            .I(N__13325));
    CascadeMux I__2602 (
            .O(N__13325),
            .I(N__13322));
    CascadeBuf I__2601 (
            .O(N__13322),
            .I(N__13319));
    CascadeMux I__2600 (
            .O(N__13319),
            .I(N__13316));
    CascadeBuf I__2599 (
            .O(N__13316),
            .I(N__13313));
    CascadeMux I__2598 (
            .O(N__13313),
            .I(N__13310));
    CascadeBuf I__2597 (
            .O(N__13310),
            .I(N__13307));
    CascadeMux I__2596 (
            .O(N__13307),
            .I(N__13304));
    CascadeBuf I__2595 (
            .O(N__13304),
            .I(N__13301));
    CascadeMux I__2594 (
            .O(N__13301),
            .I(N__13298));
    CascadeBuf I__2593 (
            .O(N__13298),
            .I(N__13295));
    CascadeMux I__2592 (
            .O(N__13295),
            .I(N__13292));
    CascadeBuf I__2591 (
            .O(N__13292),
            .I(N__13289));
    CascadeMux I__2590 (
            .O(N__13289),
            .I(N__13286));
    CascadeBuf I__2589 (
            .O(N__13286),
            .I(N__13283));
    CascadeMux I__2588 (
            .O(N__13283),
            .I(N__13280));
    CascadeBuf I__2587 (
            .O(N__13280),
            .I(N__13277));
    CascadeMux I__2586 (
            .O(N__13277),
            .I(N__13274));
    InMux I__2585 (
            .O(N__13274),
            .I(N__13271));
    LocalMux I__2584 (
            .O(N__13271),
            .I(N__13266));
    InMux I__2583 (
            .O(N__13270),
            .I(N__13263));
    InMux I__2582 (
            .O(N__13269),
            .I(N__13260));
    Span12Mux_s11_v I__2581 (
            .O(N__13266),
            .I(N__13257));
    LocalMux I__2580 (
            .O(N__13263),
            .I(M_current_address_qZ0Z_5));
    LocalMux I__2579 (
            .O(N__13260),
            .I(M_current_address_qZ0Z_5));
    Odrv12 I__2578 (
            .O(N__13257),
            .I(M_current_address_qZ0Z_5));
    CascadeMux I__2577 (
            .O(N__13250),
            .I(N_402_cascade_));
    InMux I__2576 (
            .O(N__13247),
            .I(N__13244));
    LocalMux I__2575 (
            .O(N__13244),
            .I(M_current_address_q_RNO_1Z0Z_1));
    CascadeMux I__2574 (
            .O(N__13241),
            .I(N__13238));
    CascadeBuf I__2573 (
            .O(N__13238),
            .I(N__13235));
    CascadeMux I__2572 (
            .O(N__13235),
            .I(N__13232));
    CascadeBuf I__2571 (
            .O(N__13232),
            .I(N__13229));
    CascadeMux I__2570 (
            .O(N__13229),
            .I(N__13226));
    CascadeBuf I__2569 (
            .O(N__13226),
            .I(N__13223));
    CascadeMux I__2568 (
            .O(N__13223),
            .I(N__13220));
    CascadeBuf I__2567 (
            .O(N__13220),
            .I(N__13217));
    CascadeMux I__2566 (
            .O(N__13217),
            .I(N__13214));
    CascadeBuf I__2565 (
            .O(N__13214),
            .I(N__13211));
    CascadeMux I__2564 (
            .O(N__13211),
            .I(N__13208));
    CascadeBuf I__2563 (
            .O(N__13208),
            .I(N__13205));
    CascadeMux I__2562 (
            .O(N__13205),
            .I(N__13202));
    CascadeBuf I__2561 (
            .O(N__13202),
            .I(N__13199));
    CascadeMux I__2560 (
            .O(N__13199),
            .I(N__13196));
    CascadeBuf I__2559 (
            .O(N__13196),
            .I(N__13193));
    CascadeMux I__2558 (
            .O(N__13193),
            .I(N__13190));
    CascadeBuf I__2557 (
            .O(N__13190),
            .I(N__13187));
    CascadeMux I__2556 (
            .O(N__13187),
            .I(N__13184));
    CascadeBuf I__2555 (
            .O(N__13184),
            .I(N__13181));
    CascadeMux I__2554 (
            .O(N__13181),
            .I(N__13178));
    CascadeBuf I__2553 (
            .O(N__13178),
            .I(N__13175));
    CascadeMux I__2552 (
            .O(N__13175),
            .I(N__13172));
    CascadeBuf I__2551 (
            .O(N__13172),
            .I(N__13169));
    CascadeMux I__2550 (
            .O(N__13169),
            .I(N__13166));
    CascadeBuf I__2549 (
            .O(N__13166),
            .I(N__13163));
    CascadeMux I__2548 (
            .O(N__13163),
            .I(N__13160));
    CascadeBuf I__2547 (
            .O(N__13160),
            .I(N__13157));
    CascadeMux I__2546 (
            .O(N__13157),
            .I(N__13154));
    CascadeBuf I__2545 (
            .O(N__13154),
            .I(N__13151));
    CascadeMux I__2544 (
            .O(N__13151),
            .I(N__13148));
    InMux I__2543 (
            .O(N__13148),
            .I(N__13145));
    LocalMux I__2542 (
            .O(N__13145),
            .I(N__13142));
    Span4Mux_v I__2541 (
            .O(N__13142),
            .I(N__13139));
    Span4Mux_h I__2540 (
            .O(N__13139),
            .I(N__13136));
    Span4Mux_h I__2539 (
            .O(N__13136),
            .I(N__13131));
    InMux I__2538 (
            .O(N__13135),
            .I(N__13128));
    InMux I__2537 (
            .O(N__13134),
            .I(N__13125));
    Span4Mux_v I__2536 (
            .O(N__13131),
            .I(N__13122));
    LocalMux I__2535 (
            .O(N__13128),
            .I(M_current_address_qZ0Z_1));
    LocalMux I__2534 (
            .O(N__13125),
            .I(M_current_address_qZ0Z_1));
    Odrv4 I__2533 (
            .O(N__13122),
            .I(M_current_address_qZ0Z_1));
    CascadeMux I__2532 (
            .O(N__13115),
            .I(m32_am_cascade_));
    InMux I__2531 (
            .O(N__13112),
            .I(N__13109));
    LocalMux I__2530 (
            .O(N__13109),
            .I(m7_bm));
    InMux I__2529 (
            .O(N__13106),
            .I(N__13103));
    LocalMux I__2528 (
            .O(N__13103),
            .I(m32_bm));
    InMux I__2527 (
            .O(N__13100),
            .I(N__13096));
    InMux I__2526 (
            .O(N__13099),
            .I(N__13093));
    LocalMux I__2525 (
            .O(N__13096),
            .I(N__13090));
    LocalMux I__2524 (
            .O(N__13093),
            .I(N__13087));
    Odrv4 I__2523 (
            .O(N__13090),
            .I(m32_ns));
    Odrv4 I__2522 (
            .O(N__13087),
            .I(m32_ns));
    InMux I__2521 (
            .O(N__13082),
            .I(N__13079));
    LocalMux I__2520 (
            .O(N__13079),
            .I(N__13076));
    Span4Mux_h I__2519 (
            .O(N__13076),
            .I(N__13073));
    Odrv4 I__2518 (
            .O(N__13073),
            .I(rgb_2_4));
    InMux I__2517 (
            .O(N__13070),
            .I(N__13067));
    LocalMux I__2516 (
            .O(N__13067),
            .I(N__13063));
    InMux I__2515 (
            .O(N__13066),
            .I(N__13060));
    Odrv12 I__2514 (
            .O(N__13063),
            .I(m29));
    LocalMux I__2513 (
            .O(N__13060),
            .I(m29));
    InMux I__2512 (
            .O(N__13055),
            .I(N__13052));
    LocalMux I__2511 (
            .O(N__13052),
            .I(N__13049));
    Span12Mux_h I__2510 (
            .O(N__13049),
            .I(N__13046));
    Odrv12 I__2509 (
            .O(N__13046),
            .I(\this_vga_signals.rgb_bmZ0Z_3 ));
    InMux I__2508 (
            .O(N__13043),
            .I(un1_M_current_address_q_cry_12));
    InMux I__2507 (
            .O(N__13040),
            .I(N__13033));
    InMux I__2506 (
            .O(N__13039),
            .I(N__13033));
    InMux I__2505 (
            .O(N__13038),
            .I(N__13029));
    LocalMux I__2504 (
            .O(N__13033),
            .I(N__13026));
    InMux I__2503 (
            .O(N__13032),
            .I(N__13023));
    LocalMux I__2502 (
            .O(N__13029),
            .I(N__13020));
    Span4Mux_h I__2501 (
            .O(N__13026),
            .I(N__13017));
    LocalMux I__2500 (
            .O(N__13023),
            .I(\this_pixel_clock.M_counter_qZ0Z_0 ));
    Odrv4 I__2499 (
            .O(N__13020),
            .I(\this_pixel_clock.M_counter_qZ0Z_0 ));
    Odrv4 I__2498 (
            .O(N__13017),
            .I(\this_pixel_clock.M_counter_qZ0Z_0 ));
    CascadeMux I__2497 (
            .O(N__13010),
            .I(N__13003));
    InMux I__2496 (
            .O(N__13009),
            .I(N__12998));
    InMux I__2495 (
            .O(N__13008),
            .I(N__12998));
    InMux I__2494 (
            .O(N__13007),
            .I(N__12995));
    InMux I__2493 (
            .O(N__13006),
            .I(N__12992));
    InMux I__2492 (
            .O(N__13003),
            .I(N__12989));
    LocalMux I__2491 (
            .O(N__12998),
            .I(N__12981));
    LocalMux I__2490 (
            .O(N__12995),
            .I(N__12981));
    LocalMux I__2489 (
            .O(N__12992),
            .I(N__12976));
    LocalMux I__2488 (
            .O(N__12989),
            .I(N__12976));
    CascadeMux I__2487 (
            .O(N__12988),
            .I(N__12973));
    InMux I__2486 (
            .O(N__12987),
            .I(N__12968));
    InMux I__2485 (
            .O(N__12986),
            .I(N__12968));
    Span4Mux_v I__2484 (
            .O(N__12981),
            .I(N__12963));
    Span4Mux_v I__2483 (
            .O(N__12976),
            .I(N__12963));
    InMux I__2482 (
            .O(N__12973),
            .I(N__12960));
    LocalMux I__2481 (
            .O(N__12968),
            .I(N__12955));
    Span4Mux_h I__2480 (
            .O(N__12963),
            .I(N__12952));
    LocalMux I__2479 (
            .O(N__12960),
            .I(N__12949));
    InMux I__2478 (
            .O(N__12959),
            .I(N__12946));
    InMux I__2477 (
            .O(N__12958),
            .I(N__12943));
    Span4Mux_v I__2476 (
            .O(N__12955),
            .I(N__12940));
    Sp12to4 I__2475 (
            .O(N__12952),
            .I(N__12931));
    Span12Mux_s8_h I__2474 (
            .O(N__12949),
            .I(N__12931));
    LocalMux I__2473 (
            .O(N__12946),
            .I(N__12931));
    LocalMux I__2472 (
            .O(N__12943),
            .I(N__12931));
    Odrv4 I__2471 (
            .O(N__12940),
            .I(M_this_vram_read_data_3));
    Odrv12 I__2470 (
            .O(N__12931),
            .I(M_this_vram_read_data_3));
    InMux I__2469 (
            .O(N__12926),
            .I(N__12923));
    LocalMux I__2468 (
            .O(N__12923),
            .I(N__12920));
    Span4Mux_v I__2467 (
            .O(N__12920),
            .I(N__12917));
    Span4Mux_h I__2466 (
            .O(N__12917),
            .I(N__12914));
    Span4Mux_h I__2465 (
            .O(N__12914),
            .I(N__12911));
    Odrv4 I__2464 (
            .O(N__12911),
            .I(\this_vga_signals.rgb_bmZ0Z_0 ));
    InMux I__2463 (
            .O(N__12908),
            .I(N__12905));
    LocalMux I__2462 (
            .O(N__12905),
            .I(N__12902));
    Odrv12 I__2461 (
            .O(N__12902),
            .I(\this_vga_signals.rgb_bmZ0Z_2 ));
    CascadeMux I__2460 (
            .O(N__12899),
            .I(m7_am_cascade_));
    InMux I__2459 (
            .O(N__12896),
            .I(N__12893));
    LocalMux I__2458 (
            .O(N__12893),
            .I(m7_ns));
    CascadeMux I__2457 (
            .O(N__12890),
            .I(m28_cascade_));
    InMux I__2456 (
            .O(N__12887),
            .I(un1_M_current_address_q_cry_3));
    InMux I__2455 (
            .O(N__12884),
            .I(un1_M_current_address_q_cry_4));
    InMux I__2454 (
            .O(N__12881),
            .I(un1_M_current_address_q_cry_5));
    InMux I__2453 (
            .O(N__12878),
            .I(un1_M_current_address_q_cry_6));
    InMux I__2452 (
            .O(N__12875),
            .I(bfn_15_22_0_));
    InMux I__2451 (
            .O(N__12872),
            .I(un1_M_current_address_q_cry_8));
    InMux I__2450 (
            .O(N__12869),
            .I(un1_M_current_address_q_cry_9));
    InMux I__2449 (
            .O(N__12866),
            .I(un1_M_current_address_q_cry_10));
    InMux I__2448 (
            .O(N__12863),
            .I(un1_M_current_address_q_cry_11));
    CascadeMux I__2447 (
            .O(N__12860),
            .I(N_349_0_cascade_));
    InMux I__2446 (
            .O(N__12857),
            .I(N__12852));
    InMux I__2445 (
            .O(N__12856),
            .I(N__12847));
    InMux I__2444 (
            .O(N__12855),
            .I(N__12847));
    LocalMux I__2443 (
            .O(N__12852),
            .I(N__12842));
    LocalMux I__2442 (
            .O(N__12847),
            .I(N__12842));
    Span4Mux_v I__2441 (
            .O(N__12842),
            .I(N__12838));
    InMux I__2440 (
            .O(N__12841),
            .I(N__12835));
    Sp12to4 I__2439 (
            .O(N__12838),
            .I(N__12830));
    LocalMux I__2438 (
            .O(N__12835),
            .I(N__12830));
    Span12Mux_h I__2437 (
            .O(N__12830),
            .I(N__12827));
    Odrv12 I__2436 (
            .O(N__12827),
            .I(port_enb_c));
    InMux I__2435 (
            .O(N__12824),
            .I(N__12818));
    InMux I__2434 (
            .O(N__12823),
            .I(N__12811));
    InMux I__2433 (
            .O(N__12822),
            .I(N__12811));
    InMux I__2432 (
            .O(N__12821),
            .I(N__12811));
    LocalMux I__2431 (
            .O(N__12818),
            .I(N__12808));
    LocalMux I__2430 (
            .O(N__12811),
            .I(N__12805));
    Odrv4 I__2429 (
            .O(N__12808),
            .I(\this_delay_clk.M_this_delay_clk_out_0 ));
    Odrv4 I__2428 (
            .O(N__12805),
            .I(\this_delay_clk.M_this_delay_clk_out_0 ));
    InMux I__2427 (
            .O(N__12800),
            .I(N__12797));
    LocalMux I__2426 (
            .O(N__12797),
            .I(debug_0));
    InMux I__2425 (
            .O(N__12794),
            .I(N__12791));
    LocalMux I__2424 (
            .O(N__12791),
            .I(N__12788));
    Span4Mux_v I__2423 (
            .O(N__12788),
            .I(N__12785));
    Sp12to4 I__2422 (
            .O(N__12785),
            .I(N__12782));
    Span12Mux_h I__2421 (
            .O(N__12782),
            .I(N__12778));
    InMux I__2420 (
            .O(N__12781),
            .I(N__12775));
    Odrv12 I__2419 (
            .O(N__12778),
            .I(port_rw_c));
    LocalMux I__2418 (
            .O(N__12775),
            .I(port_rw_c));
    InMux I__2417 (
            .O(N__12770),
            .I(N__12767));
    LocalMux I__2416 (
            .O(N__12767),
            .I(N__12764));
    Span4Mux_v I__2415 (
            .O(N__12764),
            .I(N__12761));
    Sp12to4 I__2414 (
            .O(N__12761),
            .I(N__12758));
    Span12Mux_h I__2413 (
            .O(N__12758),
            .I(N__12755));
    Span12Mux_v I__2412 (
            .O(N__12755),
            .I(N__12752));
    Odrv12 I__2411 (
            .O(N__12752),
            .I(port_address_c_7));
    CascadeMux I__2410 (
            .O(N__12749),
            .I(debug_0_cascade_));
    CascadeMux I__2409 (
            .O(N__12746),
            .I(N__12741));
    InMux I__2408 (
            .O(N__12745),
            .I(N__12734));
    InMux I__2407 (
            .O(N__12744),
            .I(N__12734));
    InMux I__2406 (
            .O(N__12741),
            .I(N__12734));
    LocalMux I__2405 (
            .O(N__12734),
            .I(this_start_data_delay_M_last_q));
    CascadeMux I__2404 (
            .O(N__12731),
            .I(N__12728));
    CascadeBuf I__2403 (
            .O(N__12728),
            .I(N__12725));
    CascadeMux I__2402 (
            .O(N__12725),
            .I(N__12722));
    CascadeBuf I__2401 (
            .O(N__12722),
            .I(N__12719));
    CascadeMux I__2400 (
            .O(N__12719),
            .I(N__12716));
    CascadeBuf I__2399 (
            .O(N__12716),
            .I(N__12713));
    CascadeMux I__2398 (
            .O(N__12713),
            .I(N__12710));
    CascadeBuf I__2397 (
            .O(N__12710),
            .I(N__12707));
    CascadeMux I__2396 (
            .O(N__12707),
            .I(N__12704));
    CascadeBuf I__2395 (
            .O(N__12704),
            .I(N__12701));
    CascadeMux I__2394 (
            .O(N__12701),
            .I(N__12698));
    CascadeBuf I__2393 (
            .O(N__12698),
            .I(N__12695));
    CascadeMux I__2392 (
            .O(N__12695),
            .I(N__12692));
    CascadeBuf I__2391 (
            .O(N__12692),
            .I(N__12689));
    CascadeMux I__2390 (
            .O(N__12689),
            .I(N__12686));
    CascadeBuf I__2389 (
            .O(N__12686),
            .I(N__12683));
    CascadeMux I__2388 (
            .O(N__12683),
            .I(N__12680));
    CascadeBuf I__2387 (
            .O(N__12680),
            .I(N__12677));
    CascadeMux I__2386 (
            .O(N__12677),
            .I(N__12674));
    CascadeBuf I__2385 (
            .O(N__12674),
            .I(N__12671));
    CascadeMux I__2384 (
            .O(N__12671),
            .I(N__12668));
    CascadeBuf I__2383 (
            .O(N__12668),
            .I(N__12665));
    CascadeMux I__2382 (
            .O(N__12665),
            .I(N__12662));
    CascadeBuf I__2381 (
            .O(N__12662),
            .I(N__12659));
    CascadeMux I__2380 (
            .O(N__12659),
            .I(N__12656));
    CascadeBuf I__2379 (
            .O(N__12656),
            .I(N__12653));
    CascadeMux I__2378 (
            .O(N__12653),
            .I(N__12650));
    CascadeBuf I__2377 (
            .O(N__12650),
            .I(N__12647));
    CascadeMux I__2376 (
            .O(N__12647),
            .I(N__12644));
    CascadeBuf I__2375 (
            .O(N__12644),
            .I(N__12641));
    CascadeMux I__2374 (
            .O(N__12641),
            .I(N__12638));
    InMux I__2373 (
            .O(N__12638),
            .I(N__12635));
    LocalMux I__2372 (
            .O(N__12635),
            .I(N__12632));
    Sp12to4 I__2371 (
            .O(N__12632),
            .I(N__12629));
    Span12Mux_s4_v I__2370 (
            .O(N__12629),
            .I(N__12624));
    InMux I__2369 (
            .O(N__12628),
            .I(N__12621));
    InMux I__2368 (
            .O(N__12627),
            .I(N__12618));
    Span12Mux_h I__2367 (
            .O(N__12624),
            .I(N__12615));
    LocalMux I__2366 (
            .O(N__12621),
            .I(M_current_address_qZ0Z_0));
    LocalMux I__2365 (
            .O(N__12618),
            .I(M_current_address_qZ0Z_0));
    Odrv12 I__2364 (
            .O(N__12615),
            .I(M_current_address_qZ0Z_0));
    CascadeMux I__2363 (
            .O(N__12608),
            .I(N__12604));
    InMux I__2362 (
            .O(N__12607),
            .I(N__12601));
    InMux I__2361 (
            .O(N__12604),
            .I(N__12598));
    LocalMux I__2360 (
            .O(N__12601),
            .I(N_312_0));
    LocalMux I__2359 (
            .O(N__12598),
            .I(N_312_0));
    InMux I__2358 (
            .O(N__12593),
            .I(N__12590));
    LocalMux I__2357 (
            .O(N__12590),
            .I(M_current_address_q_RNO_1Z0Z_0));
    InMux I__2356 (
            .O(N__12587),
            .I(un1_M_current_address_q_cry_0));
    InMux I__2355 (
            .O(N__12584),
            .I(un1_M_current_address_q_cry_1));
    InMux I__2354 (
            .O(N__12581),
            .I(un1_M_current_address_q_cry_2));
    InMux I__2353 (
            .O(N__12578),
            .I(N__12575));
    LocalMux I__2352 (
            .O(N__12575),
            .I(\this_vga_signals.if_N_16_i_0 ));
    InMux I__2351 (
            .O(N__12572),
            .I(N__12569));
    LocalMux I__2350 (
            .O(N__12569),
            .I(N__12566));
    Odrv12 I__2349 (
            .O(N__12566),
            .I(\this_vga_signals.g0_1_N_5L8 ));
    InMux I__2348 (
            .O(N__12563),
            .I(N__12559));
    InMux I__2347 (
            .O(N__12562),
            .I(N__12556));
    LocalMux I__2346 (
            .O(N__12559),
            .I(N__12553));
    LocalMux I__2345 (
            .O(N__12556),
            .I(N__12549));
    Span12Mux_h I__2344 (
            .O(N__12553),
            .I(N__12545));
    InMux I__2343 (
            .O(N__12552),
            .I(N__12542));
    Span4Mux_h I__2342 (
            .O(N__12549),
            .I(N__12539));
    InMux I__2341 (
            .O(N__12548),
            .I(N__12536));
    Odrv12 I__2340 (
            .O(N__12545),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2339 (
            .O(N__12542),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    Odrv4 I__2338 (
            .O(N__12539),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__2337 (
            .O(N__12536),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    InMux I__2336 (
            .O(N__12527),
            .I(N__12524));
    LocalMux I__2335 (
            .O(N__12524),
            .I(N__12520));
    CascadeMux I__2334 (
            .O(N__12523),
            .I(N__12517));
    Span4Mux_v I__2333 (
            .O(N__12520),
            .I(N__12513));
    InMux I__2332 (
            .O(N__12517),
            .I(N__12510));
    InMux I__2331 (
            .O(N__12516),
            .I(N__12505));
    Sp12to4 I__2330 (
            .O(N__12513),
            .I(N__12500));
    LocalMux I__2329 (
            .O(N__12510),
            .I(N__12500));
    InMux I__2328 (
            .O(N__12509),
            .I(N__12497));
    InMux I__2327 (
            .O(N__12508),
            .I(N__12494));
    LocalMux I__2326 (
            .O(N__12505),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    Odrv12 I__2325 (
            .O(N__12500),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2324 (
            .O(N__12497),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    LocalMux I__2323 (
            .O(N__12494),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_d ));
    InMux I__2322 (
            .O(N__12485),
            .I(N__12482));
    LocalMux I__2321 (
            .O(N__12482),
            .I(N__12479));
    Odrv12 I__2320 (
            .O(N__12479),
            .I(\this_vga_signals.g0_1_N_3L3 ));
    InMux I__2319 (
            .O(N__12476),
            .I(N__12470));
    InMux I__2318 (
            .O(N__12475),
            .I(N__12467));
    InMux I__2317 (
            .O(N__12474),
            .I(N__12464));
    InMux I__2316 (
            .O(N__12473),
            .I(N__12461));
    LocalMux I__2315 (
            .O(N__12470),
            .I(N__12456));
    LocalMux I__2314 (
            .O(N__12467),
            .I(N__12453));
    LocalMux I__2313 (
            .O(N__12464),
            .I(N__12448));
    LocalMux I__2312 (
            .O(N__12461),
            .I(N__12448));
    InMux I__2311 (
            .O(N__12460),
            .I(N__12445));
    InMux I__2310 (
            .O(N__12459),
            .I(N__12442));
    Span4Mux_v I__2309 (
            .O(N__12456),
            .I(N__12437));
    Span4Mux_v I__2308 (
            .O(N__12453),
            .I(N__12434));
    Span4Mux_v I__2307 (
            .O(N__12448),
            .I(N__12429));
    LocalMux I__2306 (
            .O(N__12445),
            .I(N__12429));
    LocalMux I__2305 (
            .O(N__12442),
            .I(N__12426));
    InMux I__2304 (
            .O(N__12441),
            .I(N__12423));
    InMux I__2303 (
            .O(N__12440),
            .I(N__12420));
    Span4Mux_v I__2302 (
            .O(N__12437),
            .I(N__12415));
    Span4Mux_v I__2301 (
            .O(N__12434),
            .I(N__12415));
    Span4Mux_h I__2300 (
            .O(N__12429),
            .I(N__12410));
    Span4Mux_v I__2299 (
            .O(N__12426),
            .I(N__12410));
    LocalMux I__2298 (
            .O(N__12423),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2297 (
            .O(N__12420),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__2296 (
            .O(N__12415),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__2295 (
            .O(N__12410),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    CascadeMux I__2294 (
            .O(N__12401),
            .I(\this_vga_signals.g0_1_N_6L11_cascade_ ));
    CascadeMux I__2293 (
            .O(N__12398),
            .I(N__12395));
    InMux I__2292 (
            .O(N__12395),
            .I(N__12391));
    InMux I__2291 (
            .O(N__12394),
            .I(N__12387));
    LocalMux I__2290 (
            .O(N__12391),
            .I(N__12384));
    InMux I__2289 (
            .O(N__12390),
            .I(N__12381));
    LocalMux I__2288 (
            .O(N__12387),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    Odrv4 I__2287 (
            .O(N__12384),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    LocalMux I__2286 (
            .O(N__12381),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    InMux I__2285 (
            .O(N__12374),
            .I(N__12371));
    LocalMux I__2284 (
            .O(N__12371),
            .I(\this_vga_signals.g0_1_N_7L13 ));
    CascadeMux I__2283 (
            .O(N__12368),
            .I(\this_vga_signals.g0_1_N_8L15_cascade_ ));
    CascadeMux I__2282 (
            .O(N__12365),
            .I(N__12360));
    CascadeMux I__2281 (
            .O(N__12364),
            .I(N__12357));
    CascadeMux I__2280 (
            .O(N__12363),
            .I(N__12344));
    InMux I__2279 (
            .O(N__12360),
            .I(N__12337));
    InMux I__2278 (
            .O(N__12357),
            .I(N__12337));
    InMux I__2277 (
            .O(N__12356),
            .I(N__12337));
    CascadeMux I__2276 (
            .O(N__12355),
            .I(N__12327));
    CascadeMux I__2275 (
            .O(N__12354),
            .I(N__12324));
    InMux I__2274 (
            .O(N__12353),
            .I(N__12321));
    InMux I__2273 (
            .O(N__12352),
            .I(N__12316));
    InMux I__2272 (
            .O(N__12351),
            .I(N__12316));
    InMux I__2271 (
            .O(N__12350),
            .I(N__12313));
    InMux I__2270 (
            .O(N__12349),
            .I(N__12306));
    InMux I__2269 (
            .O(N__12348),
            .I(N__12306));
    InMux I__2268 (
            .O(N__12347),
            .I(N__12306));
    InMux I__2267 (
            .O(N__12344),
            .I(N__12301));
    LocalMux I__2266 (
            .O(N__12337),
            .I(N__12298));
    InMux I__2265 (
            .O(N__12336),
            .I(N__12294));
    InMux I__2264 (
            .O(N__12335),
            .I(N__12291));
    InMux I__2263 (
            .O(N__12334),
            .I(N__12286));
    InMux I__2262 (
            .O(N__12333),
            .I(N__12286));
    InMux I__2261 (
            .O(N__12332),
            .I(N__12281));
    InMux I__2260 (
            .O(N__12331),
            .I(N__12281));
    InMux I__2259 (
            .O(N__12330),
            .I(N__12278));
    InMux I__2258 (
            .O(N__12327),
            .I(N__12273));
    InMux I__2257 (
            .O(N__12324),
            .I(N__12273));
    LocalMux I__2256 (
            .O(N__12321),
            .I(N__12264));
    LocalMux I__2255 (
            .O(N__12316),
            .I(N__12264));
    LocalMux I__2254 (
            .O(N__12313),
            .I(N__12264));
    LocalMux I__2253 (
            .O(N__12306),
            .I(N__12264));
    InMux I__2252 (
            .O(N__12305),
            .I(N__12259));
    InMux I__2251 (
            .O(N__12304),
            .I(N__12259));
    LocalMux I__2250 (
            .O(N__12301),
            .I(N__12254));
    Span4Mux_h I__2249 (
            .O(N__12298),
            .I(N__12251));
    InMux I__2248 (
            .O(N__12297),
            .I(N__12248));
    LocalMux I__2247 (
            .O(N__12294),
            .I(N__12242));
    LocalMux I__2246 (
            .O(N__12291),
            .I(N__12242));
    LocalMux I__2245 (
            .O(N__12286),
            .I(N__12237));
    LocalMux I__2244 (
            .O(N__12281),
            .I(N__12237));
    LocalMux I__2243 (
            .O(N__12278),
            .I(N__12234));
    LocalMux I__2242 (
            .O(N__12273),
            .I(N__12227));
    Span4Mux_v I__2241 (
            .O(N__12264),
            .I(N__12227));
    LocalMux I__2240 (
            .O(N__12259),
            .I(N__12227));
    InMux I__2239 (
            .O(N__12258),
            .I(N__12224));
    InMux I__2238 (
            .O(N__12257),
            .I(N__12221));
    Span4Mux_v I__2237 (
            .O(N__12254),
            .I(N__12218));
    Span4Mux_v I__2236 (
            .O(N__12251),
            .I(N__12215));
    LocalMux I__2235 (
            .O(N__12248),
            .I(N__12212));
    InMux I__2234 (
            .O(N__12247),
            .I(N__12209));
    Span4Mux_v I__2233 (
            .O(N__12242),
            .I(N__12204));
    Span4Mux_v I__2232 (
            .O(N__12237),
            .I(N__12204));
    Span4Mux_v I__2231 (
            .O(N__12234),
            .I(N__12199));
    Span4Mux_h I__2230 (
            .O(N__12227),
            .I(N__12199));
    LocalMux I__2229 (
            .O(N__12224),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2228 (
            .O(N__12221),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2227 (
            .O(N__12218),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2226 (
            .O(N__12215),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv12 I__2225 (
            .O(N__12212),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2224 (
            .O(N__12209),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2223 (
            .O(N__12204),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2222 (
            .O(N__12199),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    CascadeMux I__2221 (
            .O(N__12182),
            .I(N__12175));
    InMux I__2220 (
            .O(N__12181),
            .I(N__12165));
    InMux I__2219 (
            .O(N__12180),
            .I(N__12162));
    InMux I__2218 (
            .O(N__12179),
            .I(N__12157));
    InMux I__2217 (
            .O(N__12178),
            .I(N__12157));
    InMux I__2216 (
            .O(N__12175),
            .I(N__12152));
    InMux I__2215 (
            .O(N__12174),
            .I(N__12152));
    InMux I__2214 (
            .O(N__12173),
            .I(N__12149));
    InMux I__2213 (
            .O(N__12172),
            .I(N__12144));
    InMux I__2212 (
            .O(N__12171),
            .I(N__12144));
    CascadeMux I__2211 (
            .O(N__12170),
            .I(N__12141));
    InMux I__2210 (
            .O(N__12169),
            .I(N__12135));
    InMux I__2209 (
            .O(N__12168),
            .I(N__12132));
    LocalMux I__2208 (
            .O(N__12165),
            .I(N__12127));
    LocalMux I__2207 (
            .O(N__12162),
            .I(N__12127));
    LocalMux I__2206 (
            .O(N__12157),
            .I(N__12124));
    LocalMux I__2205 (
            .O(N__12152),
            .I(N__12117));
    LocalMux I__2204 (
            .O(N__12149),
            .I(N__12117));
    LocalMux I__2203 (
            .O(N__12144),
            .I(N__12117));
    InMux I__2202 (
            .O(N__12141),
            .I(N__12114));
    InMux I__2201 (
            .O(N__12140),
            .I(N__12109));
    InMux I__2200 (
            .O(N__12139),
            .I(N__12109));
    CascadeMux I__2199 (
            .O(N__12138),
            .I(N__12105));
    LocalMux I__2198 (
            .O(N__12135),
            .I(N__12102));
    LocalMux I__2197 (
            .O(N__12132),
            .I(N__12095));
    Span4Mux_h I__2196 (
            .O(N__12127),
            .I(N__12095));
    Span4Mux_h I__2195 (
            .O(N__12124),
            .I(N__12095));
    Span4Mux_h I__2194 (
            .O(N__12117),
            .I(N__12092));
    LocalMux I__2193 (
            .O(N__12114),
            .I(N__12087));
    LocalMux I__2192 (
            .O(N__12109),
            .I(N__12087));
    InMux I__2191 (
            .O(N__12108),
            .I(N__12084));
    InMux I__2190 (
            .O(N__12105),
            .I(N__12081));
    Span4Mux_h I__2189 (
            .O(N__12102),
            .I(N__12076));
    Span4Mux_v I__2188 (
            .O(N__12095),
            .I(N__12076));
    Span4Mux_h I__2187 (
            .O(N__12092),
            .I(N__12073));
    Span4Mux_v I__2186 (
            .O(N__12087),
            .I(N__12070));
    LocalMux I__2185 (
            .O(N__12084),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__2184 (
            .O(N__12081),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2183 (
            .O(N__12076),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2182 (
            .O(N__12073),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2181 (
            .O(N__12070),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    InMux I__2180 (
            .O(N__12059),
            .I(N__12052));
    InMux I__2179 (
            .O(N__12058),
            .I(N__12049));
    InMux I__2178 (
            .O(N__12057),
            .I(N__12046));
    InMux I__2177 (
            .O(N__12056),
            .I(N__12041));
    InMux I__2176 (
            .O(N__12055),
            .I(N__12041));
    LocalMux I__2175 (
            .O(N__12052),
            .I(\this_vga_signals.mult1_un68_sum_axb2_0 ));
    LocalMux I__2174 (
            .O(N__12049),
            .I(\this_vga_signals.mult1_un68_sum_axb2_0 ));
    LocalMux I__2173 (
            .O(N__12046),
            .I(\this_vga_signals.mult1_un68_sum_axb2_0 ));
    LocalMux I__2172 (
            .O(N__12041),
            .I(\this_vga_signals.mult1_un68_sum_axb2_0 ));
    CascadeMux I__2171 (
            .O(N__12032),
            .I(\this_vga_signals.mult1_un68_sum_c2_0_0_cascade_ ));
    InMux I__2170 (
            .O(N__12029),
            .I(N__12026));
    LocalMux I__2169 (
            .O(N__12026),
            .I(\this_vga_signals.if_N_6_3_0 ));
    CascadeMux I__2168 (
            .O(N__12023),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0_cascade_ ));
    CascadeMux I__2167 (
            .O(N__12020),
            .I(N__12017));
    CascadeBuf I__2166 (
            .O(N__12017),
            .I(N__12014));
    CascadeMux I__2165 (
            .O(N__12014),
            .I(N__12011));
    CascadeBuf I__2164 (
            .O(N__12011),
            .I(N__12008));
    CascadeMux I__2163 (
            .O(N__12008),
            .I(N__12005));
    CascadeBuf I__2162 (
            .O(N__12005),
            .I(N__12002));
    CascadeMux I__2161 (
            .O(N__12002),
            .I(N__11999));
    CascadeBuf I__2160 (
            .O(N__11999),
            .I(N__11996));
    CascadeMux I__2159 (
            .O(N__11996),
            .I(N__11993));
    CascadeBuf I__2158 (
            .O(N__11993),
            .I(N__11990));
    CascadeMux I__2157 (
            .O(N__11990),
            .I(N__11987));
    CascadeBuf I__2156 (
            .O(N__11987),
            .I(N__11984));
    CascadeMux I__2155 (
            .O(N__11984),
            .I(N__11981));
    CascadeBuf I__2154 (
            .O(N__11981),
            .I(N__11978));
    CascadeMux I__2153 (
            .O(N__11978),
            .I(N__11975));
    CascadeBuf I__2152 (
            .O(N__11975),
            .I(N__11972));
    CascadeMux I__2151 (
            .O(N__11972),
            .I(N__11969));
    CascadeBuf I__2150 (
            .O(N__11969),
            .I(N__11966));
    CascadeMux I__2149 (
            .O(N__11966),
            .I(N__11963));
    CascadeBuf I__2148 (
            .O(N__11963),
            .I(N__11960));
    CascadeMux I__2147 (
            .O(N__11960),
            .I(N__11957));
    CascadeBuf I__2146 (
            .O(N__11957),
            .I(N__11954));
    CascadeMux I__2145 (
            .O(N__11954),
            .I(N__11951));
    CascadeBuf I__2144 (
            .O(N__11951),
            .I(N__11948));
    CascadeMux I__2143 (
            .O(N__11948),
            .I(N__11945));
    CascadeBuf I__2142 (
            .O(N__11945),
            .I(N__11942));
    CascadeMux I__2141 (
            .O(N__11942),
            .I(N__11939));
    CascadeBuf I__2140 (
            .O(N__11939),
            .I(N__11936));
    CascadeMux I__2139 (
            .O(N__11936),
            .I(N__11933));
    CascadeBuf I__2138 (
            .O(N__11933),
            .I(N__11930));
    CascadeMux I__2137 (
            .O(N__11930),
            .I(N__11927));
    InMux I__2136 (
            .O(N__11927),
            .I(N__11924));
    LocalMux I__2135 (
            .O(N__11924),
            .I(N__11921));
    Sp12to4 I__2134 (
            .O(N__11921),
            .I(N__11918));
    Span12Mux_v I__2133 (
            .O(N__11918),
            .I(N__11915));
    Odrv12 I__2132 (
            .O(N__11915),
            .I(M_this_vga_signals_address_8));
    CascadeMux I__2131 (
            .O(N__11912),
            .I(N__11909));
    InMux I__2130 (
            .O(N__11909),
            .I(N__11906));
    LocalMux I__2129 (
            .O(N__11906),
            .I(N_401));
    CascadeMux I__2128 (
            .O(N__11903),
            .I(N__11898));
    InMux I__2127 (
            .O(N__11902),
            .I(N__11893));
    InMux I__2126 (
            .O(N__11901),
            .I(N__11888));
    InMux I__2125 (
            .O(N__11898),
            .I(N__11888));
    InMux I__2124 (
            .O(N__11897),
            .I(N__11885));
    InMux I__2123 (
            .O(N__11896),
            .I(N__11882));
    LocalMux I__2122 (
            .O(N__11893),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ));
    LocalMux I__2121 (
            .O(N__11888),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ));
    LocalMux I__2120 (
            .O(N__11885),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ));
    LocalMux I__2119 (
            .O(N__11882),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ));
    InMux I__2118 (
            .O(N__11873),
            .I(N__11867));
    InMux I__2117 (
            .O(N__11872),
            .I(N__11864));
    InMux I__2116 (
            .O(N__11871),
            .I(N__11859));
    InMux I__2115 (
            .O(N__11870),
            .I(N__11859));
    LocalMux I__2114 (
            .O(N__11867),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ));
    LocalMux I__2113 (
            .O(N__11864),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ));
    LocalMux I__2112 (
            .O(N__11859),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ));
    CascadeMux I__2111 (
            .O(N__11852),
            .I(N__11849));
    CascadeBuf I__2110 (
            .O(N__11849),
            .I(N__11846));
    CascadeMux I__2109 (
            .O(N__11846),
            .I(N__11843));
    CascadeBuf I__2108 (
            .O(N__11843),
            .I(N__11840));
    CascadeMux I__2107 (
            .O(N__11840),
            .I(N__11837));
    CascadeBuf I__2106 (
            .O(N__11837),
            .I(N__11834));
    CascadeMux I__2105 (
            .O(N__11834),
            .I(N__11831));
    CascadeBuf I__2104 (
            .O(N__11831),
            .I(N__11828));
    CascadeMux I__2103 (
            .O(N__11828),
            .I(N__11825));
    CascadeBuf I__2102 (
            .O(N__11825),
            .I(N__11822));
    CascadeMux I__2101 (
            .O(N__11822),
            .I(N__11819));
    CascadeBuf I__2100 (
            .O(N__11819),
            .I(N__11816));
    CascadeMux I__2099 (
            .O(N__11816),
            .I(N__11813));
    CascadeBuf I__2098 (
            .O(N__11813),
            .I(N__11810));
    CascadeMux I__2097 (
            .O(N__11810),
            .I(N__11807));
    CascadeBuf I__2096 (
            .O(N__11807),
            .I(N__11804));
    CascadeMux I__2095 (
            .O(N__11804),
            .I(N__11801));
    CascadeBuf I__2094 (
            .O(N__11801),
            .I(N__11798));
    CascadeMux I__2093 (
            .O(N__11798),
            .I(N__11795));
    CascadeBuf I__2092 (
            .O(N__11795),
            .I(N__11792));
    CascadeMux I__2091 (
            .O(N__11792),
            .I(N__11789));
    CascadeBuf I__2090 (
            .O(N__11789),
            .I(N__11786));
    CascadeMux I__2089 (
            .O(N__11786),
            .I(N__11783));
    CascadeBuf I__2088 (
            .O(N__11783),
            .I(N__11780));
    CascadeMux I__2087 (
            .O(N__11780),
            .I(N__11777));
    CascadeBuf I__2086 (
            .O(N__11777),
            .I(N__11774));
    CascadeMux I__2085 (
            .O(N__11774),
            .I(N__11771));
    CascadeBuf I__2084 (
            .O(N__11771),
            .I(N__11768));
    CascadeMux I__2083 (
            .O(N__11768),
            .I(N__11765));
    CascadeBuf I__2082 (
            .O(N__11765),
            .I(N__11762));
    CascadeMux I__2081 (
            .O(N__11762),
            .I(N__11759));
    InMux I__2080 (
            .O(N__11759),
            .I(N__11756));
    LocalMux I__2079 (
            .O(N__11756),
            .I(N__11753));
    Span12Mux_h I__2078 (
            .O(N__11753),
            .I(N__11750));
    Odrv12 I__2077 (
            .O(N__11750),
            .I(M_this_vga_signals_address_4));
    InMux I__2076 (
            .O(N__11747),
            .I(N__11742));
    InMux I__2075 (
            .O(N__11746),
            .I(N__11737));
    InMux I__2074 (
            .O(N__11745),
            .I(N__11737));
    LocalMux I__2073 (
            .O(N__11742),
            .I(N__11732));
    LocalMux I__2072 (
            .O(N__11737),
            .I(N__11729));
    InMux I__2071 (
            .O(N__11736),
            .I(N__11726));
    InMux I__2070 (
            .O(N__11735),
            .I(N__11723));
    Span4Mux_v I__2069 (
            .O(N__11732),
            .I(N__11720));
    Span4Mux_h I__2068 (
            .O(N__11729),
            .I(N__11715));
    LocalMux I__2067 (
            .O(N__11726),
            .I(N__11715));
    LocalMux I__2066 (
            .O(N__11723),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__2065 (
            .O(N__11720),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__2064 (
            .O(N__11715),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    InMux I__2063 (
            .O(N__11708),
            .I(N__11694));
    InMux I__2062 (
            .O(N__11707),
            .I(N__11694));
    InMux I__2061 (
            .O(N__11706),
            .I(N__11690));
    InMux I__2060 (
            .O(N__11705),
            .I(N__11677));
    InMux I__2059 (
            .O(N__11704),
            .I(N__11677));
    InMux I__2058 (
            .O(N__11703),
            .I(N__11677));
    InMux I__2057 (
            .O(N__11702),
            .I(N__11677));
    InMux I__2056 (
            .O(N__11701),
            .I(N__11670));
    InMux I__2055 (
            .O(N__11700),
            .I(N__11670));
    InMux I__2054 (
            .O(N__11699),
            .I(N__11670));
    LocalMux I__2053 (
            .O(N__11694),
            .I(N__11667));
    InMux I__2052 (
            .O(N__11693),
            .I(N__11664));
    LocalMux I__2051 (
            .O(N__11690),
            .I(N__11661));
    InMux I__2050 (
            .O(N__11689),
            .I(N__11655));
    InMux I__2049 (
            .O(N__11688),
            .I(N__11655));
    InMux I__2048 (
            .O(N__11687),
            .I(N__11650));
    InMux I__2047 (
            .O(N__11686),
            .I(N__11650));
    LocalMux I__2046 (
            .O(N__11677),
            .I(N__11647));
    LocalMux I__2045 (
            .O(N__11670),
            .I(N__11644));
    Span4Mux_h I__2044 (
            .O(N__11667),
            .I(N__11639));
    LocalMux I__2043 (
            .O(N__11664),
            .I(N__11639));
    Span12Mux_v I__2042 (
            .O(N__11661),
            .I(N__11636));
    InMux I__2041 (
            .O(N__11660),
            .I(N__11633));
    LocalMux I__2040 (
            .O(N__11655),
            .I(M_counter_q_RNIJR071_1));
    LocalMux I__2039 (
            .O(N__11650),
            .I(M_counter_q_RNIJR071_1));
    Odrv12 I__2038 (
            .O(N__11647),
            .I(M_counter_q_RNIJR071_1));
    Odrv4 I__2037 (
            .O(N__11644),
            .I(M_counter_q_RNIJR071_1));
    Odrv4 I__2036 (
            .O(N__11639),
            .I(M_counter_q_RNIJR071_1));
    Odrv12 I__2035 (
            .O(N__11636),
            .I(M_counter_q_RNIJR071_1));
    LocalMux I__2034 (
            .O(N__11633),
            .I(M_counter_q_RNIJR071_1));
    CascadeMux I__2033 (
            .O(N__11618),
            .I(N__11615));
    InMux I__2032 (
            .O(N__11615),
            .I(N__11611));
    CascadeMux I__2031 (
            .O(N__11614),
            .I(N__11607));
    LocalMux I__2030 (
            .O(N__11611),
            .I(N__11603));
    InMux I__2029 (
            .O(N__11610),
            .I(N__11600));
    InMux I__2028 (
            .O(N__11607),
            .I(N__11595));
    InMux I__2027 (
            .O(N__11606),
            .I(N__11595));
    Span4Mux_v I__2026 (
            .O(N__11603),
            .I(N__11592));
    LocalMux I__2025 (
            .O(N__11600),
            .I(N__11589));
    LocalMux I__2024 (
            .O(N__11595),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv4 I__2023 (
            .O(N__11592),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv4 I__2022 (
            .O(N__11589),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    SRMux I__2021 (
            .O(N__11582),
            .I(N__11579));
    LocalMux I__2020 (
            .O(N__11579),
            .I(N__11574));
    SRMux I__2019 (
            .O(N__11578),
            .I(N__11571));
    SRMux I__2018 (
            .O(N__11577),
            .I(N__11568));
    Span4Mux_v I__2017 (
            .O(N__11574),
            .I(N__11562));
    LocalMux I__2016 (
            .O(N__11571),
            .I(N__11562));
    LocalMux I__2015 (
            .O(N__11568),
            .I(N__11559));
    InMux I__2014 (
            .O(N__11567),
            .I(N__11556));
    Span4Mux_h I__2013 (
            .O(N__11562),
            .I(N__11553));
    Span4Mux_v I__2012 (
            .O(N__11559),
            .I(N__11550));
    LocalMux I__2011 (
            .O(N__11556),
            .I(N__11547));
    Odrv4 I__2010 (
            .O(N__11553),
            .I(M_counter_q_RNIQR4I2_1));
    Odrv4 I__2009 (
            .O(N__11550),
            .I(M_counter_q_RNIQR4I2_1));
    Odrv4 I__2008 (
            .O(N__11547),
            .I(M_counter_q_RNIQR4I2_1));
    InMux I__2007 (
            .O(N__11540),
            .I(N__11537));
    LocalMux I__2006 (
            .O(N__11537),
            .I(N__11534));
    Odrv12 I__2005 (
            .O(N__11534),
            .I(\this_vga_signals.rgb_bmZ0Z_1 ));
    InMux I__2004 (
            .O(N__11531),
            .I(N__11528));
    LocalMux I__2003 (
            .O(N__11528),
            .I(N__11525));
    Span4Mux_h I__2002 (
            .O(N__11525),
            .I(N__11522));
    Span4Mux_h I__2001 (
            .O(N__11522),
            .I(N__11519));
    Span4Mux_h I__2000 (
            .O(N__11519),
            .I(N__11516));
    Odrv4 I__1999 (
            .O(N__11516),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    InMux I__1998 (
            .O(N__11513),
            .I(N__11509));
    InMux I__1997 (
            .O(N__11512),
            .I(N__11506));
    LocalMux I__1996 (
            .O(N__11509),
            .I(N__11500));
    LocalMux I__1995 (
            .O(N__11506),
            .I(N__11497));
    InMux I__1994 (
            .O(N__11505),
            .I(N__11493));
    InMux I__1993 (
            .O(N__11504),
            .I(N__11488));
    InMux I__1992 (
            .O(N__11503),
            .I(N__11488));
    Span4Mux_h I__1991 (
            .O(N__11500),
            .I(N__11485));
    Span4Mux_h I__1990 (
            .O(N__11497),
            .I(N__11482));
    InMux I__1989 (
            .O(N__11496),
            .I(N__11479));
    LocalMux I__1988 (
            .O(N__11493),
            .I(N__11474));
    LocalMux I__1987 (
            .O(N__11488),
            .I(N__11474));
    Odrv4 I__1986 (
            .O(N__11485),
            .I(\this_vga_signals.mult1_un54_sum_axb1_5 ));
    Odrv4 I__1985 (
            .O(N__11482),
            .I(\this_vga_signals.mult1_un54_sum_axb1_5 ));
    LocalMux I__1984 (
            .O(N__11479),
            .I(\this_vga_signals.mult1_un54_sum_axb1_5 ));
    Odrv4 I__1983 (
            .O(N__11474),
            .I(\this_vga_signals.mult1_un54_sum_axb1_5 ));
    CascadeMux I__1982 (
            .O(N__11465),
            .I(N__11452));
    CascadeMux I__1981 (
            .O(N__11464),
            .I(N__11447));
    CascadeMux I__1980 (
            .O(N__11463),
            .I(N__11444));
    InMux I__1979 (
            .O(N__11462),
            .I(N__11439));
    CascadeMux I__1978 (
            .O(N__11461),
            .I(N__11432));
    CascadeMux I__1977 (
            .O(N__11460),
            .I(N__11429));
    CascadeMux I__1976 (
            .O(N__11459),
            .I(N__11423));
    CascadeMux I__1975 (
            .O(N__11458),
            .I(N__11419));
    CascadeMux I__1974 (
            .O(N__11457),
            .I(N__11414));
    CascadeMux I__1973 (
            .O(N__11456),
            .I(N__11410));
    InMux I__1972 (
            .O(N__11455),
            .I(N__11403));
    InMux I__1971 (
            .O(N__11452),
            .I(N__11396));
    InMux I__1970 (
            .O(N__11451),
            .I(N__11396));
    InMux I__1969 (
            .O(N__11450),
            .I(N__11396));
    InMux I__1968 (
            .O(N__11447),
            .I(N__11391));
    InMux I__1967 (
            .O(N__11444),
            .I(N__11388));
    InMux I__1966 (
            .O(N__11443),
            .I(N__11383));
    InMux I__1965 (
            .O(N__11442),
            .I(N__11383));
    LocalMux I__1964 (
            .O(N__11439),
            .I(N__11380));
    InMux I__1963 (
            .O(N__11438),
            .I(N__11377));
    InMux I__1962 (
            .O(N__11437),
            .I(N__11368));
    InMux I__1961 (
            .O(N__11436),
            .I(N__11368));
    InMux I__1960 (
            .O(N__11435),
            .I(N__11368));
    InMux I__1959 (
            .O(N__11432),
            .I(N__11368));
    InMux I__1958 (
            .O(N__11429),
            .I(N__11363));
    InMux I__1957 (
            .O(N__11428),
            .I(N__11363));
    InMux I__1956 (
            .O(N__11427),
            .I(N__11360));
    InMux I__1955 (
            .O(N__11426),
            .I(N__11357));
    InMux I__1954 (
            .O(N__11423),
            .I(N__11354));
    InMux I__1953 (
            .O(N__11422),
            .I(N__11349));
    InMux I__1952 (
            .O(N__11419),
            .I(N__11349));
    CascadeMux I__1951 (
            .O(N__11418),
            .I(N__11345));
    InMux I__1950 (
            .O(N__11417),
            .I(N__11342));
    InMux I__1949 (
            .O(N__11414),
            .I(N__11337));
    InMux I__1948 (
            .O(N__11413),
            .I(N__11337));
    InMux I__1947 (
            .O(N__11410),
            .I(N__11332));
    InMux I__1946 (
            .O(N__11409),
            .I(N__11332));
    CascadeMux I__1945 (
            .O(N__11408),
            .I(N__11328));
    InMux I__1944 (
            .O(N__11407),
            .I(N__11323));
    InMux I__1943 (
            .O(N__11406),
            .I(N__11323));
    LocalMux I__1942 (
            .O(N__11403),
            .I(N__11318));
    LocalMux I__1941 (
            .O(N__11396),
            .I(N__11318));
    InMux I__1940 (
            .O(N__11395),
            .I(N__11313));
    InMux I__1939 (
            .O(N__11394),
            .I(N__11313));
    LocalMux I__1938 (
            .O(N__11391),
            .I(N__11310));
    LocalMux I__1937 (
            .O(N__11388),
            .I(N__11307));
    LocalMux I__1936 (
            .O(N__11383),
            .I(N__11298));
    Span4Mux_v I__1935 (
            .O(N__11380),
            .I(N__11298));
    LocalMux I__1934 (
            .O(N__11377),
            .I(N__11298));
    LocalMux I__1933 (
            .O(N__11368),
            .I(N__11298));
    LocalMux I__1932 (
            .O(N__11363),
            .I(N__11295));
    LocalMux I__1931 (
            .O(N__11360),
            .I(N__11290));
    LocalMux I__1930 (
            .O(N__11357),
            .I(N__11290));
    LocalMux I__1929 (
            .O(N__11354),
            .I(N__11284));
    LocalMux I__1928 (
            .O(N__11349),
            .I(N__11284));
    InMux I__1927 (
            .O(N__11348),
            .I(N__11281));
    InMux I__1926 (
            .O(N__11345),
            .I(N__11278));
    LocalMux I__1925 (
            .O(N__11342),
            .I(N__11271));
    LocalMux I__1924 (
            .O(N__11337),
            .I(N__11271));
    LocalMux I__1923 (
            .O(N__11332),
            .I(N__11271));
    InMux I__1922 (
            .O(N__11331),
            .I(N__11265));
    InMux I__1921 (
            .O(N__11328),
            .I(N__11265));
    LocalMux I__1920 (
            .O(N__11323),
            .I(N__11262));
    Span4Mux_v I__1919 (
            .O(N__11318),
            .I(N__11259));
    LocalMux I__1918 (
            .O(N__11313),
            .I(N__11254));
    Span4Mux_v I__1917 (
            .O(N__11310),
            .I(N__11254));
    Span4Mux_h I__1916 (
            .O(N__11307),
            .I(N__11245));
    Span4Mux_h I__1915 (
            .O(N__11298),
            .I(N__11245));
    Span4Mux_v I__1914 (
            .O(N__11295),
            .I(N__11245));
    Span4Mux_h I__1913 (
            .O(N__11290),
            .I(N__11245));
    InMux I__1912 (
            .O(N__11289),
            .I(N__11242));
    Span4Mux_v I__1911 (
            .O(N__11284),
            .I(N__11235));
    LocalMux I__1910 (
            .O(N__11281),
            .I(N__11235));
    LocalMux I__1909 (
            .O(N__11278),
            .I(N__11235));
    Span4Mux_v I__1908 (
            .O(N__11271),
            .I(N__11232));
    InMux I__1907 (
            .O(N__11270),
            .I(N__11229));
    LocalMux I__1906 (
            .O(N__11265),
            .I(N__11226));
    Span4Mux_v I__1905 (
            .O(N__11262),
            .I(N__11219));
    Span4Mux_v I__1904 (
            .O(N__11259),
            .I(N__11219));
    Span4Mux_v I__1903 (
            .O(N__11254),
            .I(N__11219));
    Span4Mux_v I__1902 (
            .O(N__11245),
            .I(N__11216));
    LocalMux I__1901 (
            .O(N__11242),
            .I(N__11209));
    Span4Mux_h I__1900 (
            .O(N__11235),
            .I(N__11209));
    Span4Mux_h I__1899 (
            .O(N__11232),
            .I(N__11209));
    LocalMux I__1898 (
            .O(N__11229),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv12 I__1897 (
            .O(N__11226),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__1896 (
            .O(N__11219),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__1895 (
            .O(N__11216),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__1894 (
            .O(N__11209),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    CascadeMux I__1893 (
            .O(N__11198),
            .I(\this_vga_signals.if_N_13_i_i_0_cascade_ ));
    InMux I__1892 (
            .O(N__11195),
            .I(N__11187));
    InMux I__1891 (
            .O(N__11194),
            .I(N__11184));
    InMux I__1890 (
            .O(N__11193),
            .I(N__11180));
    InMux I__1889 (
            .O(N__11192),
            .I(N__11175));
    InMux I__1888 (
            .O(N__11191),
            .I(N__11175));
    InMux I__1887 (
            .O(N__11190),
            .I(N__11170));
    LocalMux I__1886 (
            .O(N__11187),
            .I(N__11166));
    LocalMux I__1885 (
            .O(N__11184),
            .I(N__11163));
    InMux I__1884 (
            .O(N__11183),
            .I(N__11160));
    LocalMux I__1883 (
            .O(N__11180),
            .I(N__11155));
    LocalMux I__1882 (
            .O(N__11175),
            .I(N__11155));
    InMux I__1881 (
            .O(N__11174),
            .I(N__11150));
    InMux I__1880 (
            .O(N__11173),
            .I(N__11150));
    LocalMux I__1879 (
            .O(N__11170),
            .I(N__11140));
    InMux I__1878 (
            .O(N__11169),
            .I(N__11137));
    Span4Mux_h I__1877 (
            .O(N__11166),
            .I(N__11126));
    Span4Mux_h I__1876 (
            .O(N__11163),
            .I(N__11126));
    LocalMux I__1875 (
            .O(N__11160),
            .I(N__11126));
    Span4Mux_v I__1874 (
            .O(N__11155),
            .I(N__11126));
    LocalMux I__1873 (
            .O(N__11150),
            .I(N__11126));
    InMux I__1872 (
            .O(N__11149),
            .I(N__11119));
    InMux I__1871 (
            .O(N__11148),
            .I(N__11119));
    InMux I__1870 (
            .O(N__11147),
            .I(N__11119));
    InMux I__1869 (
            .O(N__11146),
            .I(N__11114));
    InMux I__1868 (
            .O(N__11145),
            .I(N__11114));
    InMux I__1867 (
            .O(N__11144),
            .I(N__11109));
    InMux I__1866 (
            .O(N__11143),
            .I(N__11109));
    Odrv4 I__1865 (
            .O(N__11140),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0 ));
    LocalMux I__1864 (
            .O(N__11137),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0 ));
    Odrv4 I__1863 (
            .O(N__11126),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0 ));
    LocalMux I__1862 (
            .O(N__11119),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0 ));
    LocalMux I__1861 (
            .O(N__11114),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0 ));
    LocalMux I__1860 (
            .O(N__11109),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0 ));
    CascadeMux I__1859 (
            .O(N__11096),
            .I(\this_vga_signals.g0_1_0_0_cascade_ ));
    InMux I__1858 (
            .O(N__11093),
            .I(N__11090));
    LocalMux I__1857 (
            .O(N__11090),
            .I(N__11087));
    Odrv12 I__1856 (
            .O(N__11087),
            .I(\this_vga_signals.g4_0 ));
    CascadeMux I__1855 (
            .O(N__11084),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_d_0_cascade_ ));
    InMux I__1854 (
            .O(N__11081),
            .I(N__11078));
    LocalMux I__1853 (
            .O(N__11078),
            .I(N__11073));
    InMux I__1852 (
            .O(N__11077),
            .I(N__11070));
    InMux I__1851 (
            .O(N__11076),
            .I(N__11067));
    Odrv4 I__1850 (
            .O(N__11073),
            .I(\this_vga_signals.mult1_un68_sum_ac0_4 ));
    LocalMux I__1849 (
            .O(N__11070),
            .I(\this_vga_signals.mult1_un68_sum_ac0_4 ));
    LocalMux I__1848 (
            .O(N__11067),
            .I(\this_vga_signals.mult1_un68_sum_ac0_4 ));
    CascadeMux I__1847 (
            .O(N__11060),
            .I(\this_vga_signals.g0_i_o2_0_0_x2_0_cascade_ ));
    InMux I__1846 (
            .O(N__11057),
            .I(N__11054));
    LocalMux I__1845 (
            .O(N__11054),
            .I(\this_vga_signals.N_16 ));
    CascadeMux I__1844 (
            .O(N__11051),
            .I(N__11048));
    InMux I__1843 (
            .O(N__11048),
            .I(N__11045));
    LocalMux I__1842 (
            .O(N__11045),
            .I(N__11040));
    InMux I__1841 (
            .O(N__11044),
            .I(N__11037));
    InMux I__1840 (
            .O(N__11043),
            .I(N__11034));
    Span4Mux_v I__1839 (
            .O(N__11040),
            .I(N__11029));
    LocalMux I__1838 (
            .O(N__11037),
            .I(N__11029));
    LocalMux I__1837 (
            .O(N__11034),
            .I(N__11024));
    Span4Mux_h I__1836 (
            .O(N__11029),
            .I(N__11021));
    InMux I__1835 (
            .O(N__11028),
            .I(N__11018));
    InMux I__1834 (
            .O(N__11027),
            .I(N__11015));
    Odrv12 I__1833 (
            .O(N__11024),
            .I(\this_vga_signals.mult1_un54_sum_i_1 ));
    Odrv4 I__1832 (
            .O(N__11021),
            .I(\this_vga_signals.mult1_un54_sum_i_1 ));
    LocalMux I__1831 (
            .O(N__11018),
            .I(\this_vga_signals.mult1_un54_sum_i_1 ));
    LocalMux I__1830 (
            .O(N__11015),
            .I(\this_vga_signals.mult1_un54_sum_i_1 ));
    InMux I__1829 (
            .O(N__11006),
            .I(N__11002));
    CascadeMux I__1828 (
            .O(N__11005),
            .I(N__10999));
    LocalMux I__1827 (
            .O(N__11002),
            .I(N__10996));
    InMux I__1826 (
            .O(N__10999),
            .I(N__10993));
    Odrv4 I__1825 (
            .O(N__10996),
            .I(\this_vga_signals.if_N_1_i_0 ));
    LocalMux I__1824 (
            .O(N__10993),
            .I(\this_vga_signals.if_N_1_i_0 ));
    InMux I__1823 (
            .O(N__10988),
            .I(N__10982));
    InMux I__1822 (
            .O(N__10987),
            .I(N__10982));
    LocalMux I__1821 (
            .O(N__10982),
            .I(N__10977));
    InMux I__1820 (
            .O(N__10981),
            .I(N__10972));
    InMux I__1819 (
            .O(N__10980),
            .I(N__10972));
    Span4Mux_v I__1818 (
            .O(N__10977),
            .I(N__10959));
    LocalMux I__1817 (
            .O(N__10972),
            .I(N__10959));
    CascadeMux I__1816 (
            .O(N__10971),
            .I(N__10956));
    CascadeMux I__1815 (
            .O(N__10970),
            .I(N__10953));
    CascadeMux I__1814 (
            .O(N__10969),
            .I(N__10950));
    InMux I__1813 (
            .O(N__10968),
            .I(N__10944));
    InMux I__1812 (
            .O(N__10967),
            .I(N__10944));
    InMux I__1811 (
            .O(N__10966),
            .I(N__10937));
    InMux I__1810 (
            .O(N__10965),
            .I(N__10937));
    InMux I__1809 (
            .O(N__10964),
            .I(N__10937));
    Span4Mux_h I__1808 (
            .O(N__10959),
            .I(N__10934));
    InMux I__1807 (
            .O(N__10956),
            .I(N__10925));
    InMux I__1806 (
            .O(N__10953),
            .I(N__10925));
    InMux I__1805 (
            .O(N__10950),
            .I(N__10925));
    InMux I__1804 (
            .O(N__10949),
            .I(N__10925));
    LocalMux I__1803 (
            .O(N__10944),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1802 (
            .O(N__10937),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    Odrv4 I__1801 (
            .O(N__10934),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1800 (
            .O(N__10925),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    InMux I__1799 (
            .O(N__10916),
            .I(N__10907));
    InMux I__1798 (
            .O(N__10915),
            .I(N__10907));
    CascadeMux I__1797 (
            .O(N__10914),
            .I(N__10903));
    InMux I__1796 (
            .O(N__10913),
            .I(N__10894));
    InMux I__1795 (
            .O(N__10912),
            .I(N__10894));
    LocalMux I__1794 (
            .O(N__10907),
            .I(N__10891));
    InMux I__1793 (
            .O(N__10906),
            .I(N__10884));
    InMux I__1792 (
            .O(N__10903),
            .I(N__10884));
    InMux I__1791 (
            .O(N__10902),
            .I(N__10884));
    InMux I__1790 (
            .O(N__10901),
            .I(N__10877));
    InMux I__1789 (
            .O(N__10900),
            .I(N__10874));
    InMux I__1788 (
            .O(N__10899),
            .I(N__10871));
    LocalMux I__1787 (
            .O(N__10894),
            .I(N__10868));
    Span4Mux_h I__1786 (
            .O(N__10891),
            .I(N__10865));
    LocalMux I__1785 (
            .O(N__10884),
            .I(N__10862));
    InMux I__1784 (
            .O(N__10883),
            .I(N__10853));
    InMux I__1783 (
            .O(N__10882),
            .I(N__10853));
    InMux I__1782 (
            .O(N__10881),
            .I(N__10853));
    InMux I__1781 (
            .O(N__10880),
            .I(N__10853));
    LocalMux I__1780 (
            .O(N__10877),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1779 (
            .O(N__10874),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1778 (
            .O(N__10871),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv12 I__1777 (
            .O(N__10868),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__1776 (
            .O(N__10865),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__1775 (
            .O(N__10862),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1774 (
            .O(N__10853),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    InMux I__1773 (
            .O(N__10838),
            .I(N__10835));
    LocalMux I__1772 (
            .O(N__10835),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_0 ));
    InMux I__1771 (
            .O(N__10832),
            .I(N__10829));
    LocalMux I__1770 (
            .O(N__10829),
            .I(N__10826));
    Span4Mux_h I__1769 (
            .O(N__10826),
            .I(N__10823));
    Odrv4 I__1768 (
            .O(N__10823),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    CascadeMux I__1767 (
            .O(N__10820),
            .I(\this_vga_signals.if_m3_5_cascade_ ));
    InMux I__1766 (
            .O(N__10817),
            .I(N__10814));
    LocalMux I__1765 (
            .O(N__10814),
            .I(\this_vga_signals.if_N_3_i ));
    CascadeMux I__1764 (
            .O(N__10811),
            .I(\this_vga_signals.if_m5_4_cascade_ ));
    InMux I__1763 (
            .O(N__10808),
            .I(N__10805));
    LocalMux I__1762 (
            .O(N__10805),
            .I(\this_vga_signals.g1_1_4 ));
    InMux I__1761 (
            .O(N__10802),
            .I(N__10799));
    LocalMux I__1760 (
            .O(N__10799),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_1 ));
    CascadeMux I__1759 (
            .O(N__10796),
            .I(\this_vga_signals.mult1_un68_sum_axb2_0_1_cascade_ ));
    InMux I__1758 (
            .O(N__10793),
            .I(N__10790));
    LocalMux I__1757 (
            .O(N__10790),
            .I(\this_vga_signals.g1_1_1 ));
    InMux I__1756 (
            .O(N__10787),
            .I(N__10784));
    LocalMux I__1755 (
            .O(N__10784),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    CascadeMux I__1754 (
            .O(N__10781),
            .I(\this_vga_signals.SUM_3_cascade_ ));
    CascadeMux I__1753 (
            .O(N__10778),
            .I(N__10775));
    InMux I__1752 (
            .O(N__10775),
            .I(N__10766));
    InMux I__1751 (
            .O(N__10774),
            .I(N__10763));
    InMux I__1750 (
            .O(N__10773),
            .I(N__10758));
    InMux I__1749 (
            .O(N__10772),
            .I(N__10758));
    InMux I__1748 (
            .O(N__10771),
            .I(N__10751));
    InMux I__1747 (
            .O(N__10770),
            .I(N__10751));
    InMux I__1746 (
            .O(N__10769),
            .I(N__10751));
    LocalMux I__1745 (
            .O(N__10766),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1744 (
            .O(N__10763),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1743 (
            .O(N__10758),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1742 (
            .O(N__10751),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    CascadeMux I__1741 (
            .O(N__10742),
            .I(N__10734));
    InMux I__1740 (
            .O(N__10741),
            .I(N__10730));
    InMux I__1739 (
            .O(N__10740),
            .I(N__10727));
    InMux I__1738 (
            .O(N__10739),
            .I(N__10722));
    InMux I__1737 (
            .O(N__10738),
            .I(N__10722));
    InMux I__1736 (
            .O(N__10737),
            .I(N__10715));
    InMux I__1735 (
            .O(N__10734),
            .I(N__10715));
    InMux I__1734 (
            .O(N__10733),
            .I(N__10715));
    LocalMux I__1733 (
            .O(N__10730),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1732 (
            .O(N__10727),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1731 (
            .O(N__10722),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1730 (
            .O(N__10715),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__1729 (
            .O(N__10706),
            .I(N__10696));
    InMux I__1728 (
            .O(N__10705),
            .I(N__10696));
    CascadeMux I__1727 (
            .O(N__10704),
            .I(N__10693));
    CascadeMux I__1726 (
            .O(N__10703),
            .I(N__10690));
    InMux I__1725 (
            .O(N__10702),
            .I(N__10686));
    InMux I__1724 (
            .O(N__10701),
            .I(N__10683));
    LocalMux I__1723 (
            .O(N__10696),
            .I(N__10680));
    InMux I__1722 (
            .O(N__10693),
            .I(N__10673));
    InMux I__1721 (
            .O(N__10690),
            .I(N__10673));
    InMux I__1720 (
            .O(N__10689),
            .I(N__10673));
    LocalMux I__1719 (
            .O(N__10686),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1718 (
            .O(N__10683),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__1717 (
            .O(N__10680),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1716 (
            .O(N__10673),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    InMux I__1715 (
            .O(N__10664),
            .I(N__10661));
    LocalMux I__1714 (
            .O(N__10661),
            .I(\this_vga_signals.N_34 ));
    CascadeMux I__1713 (
            .O(N__10658),
            .I(\this_vga_signals.N_34_cascade_ ));
    InMux I__1712 (
            .O(N__10655),
            .I(N__10650));
    InMux I__1711 (
            .O(N__10654),
            .I(N__10645));
    InMux I__1710 (
            .O(N__10653),
            .I(N__10645));
    LocalMux I__1709 (
            .O(N__10650),
            .I(\this_vga_signals.SUM_3 ));
    LocalMux I__1708 (
            .O(N__10645),
            .I(\this_vga_signals.SUM_3 ));
    CascadeMux I__1707 (
            .O(N__10640),
            .I(N__10633));
    InMux I__1706 (
            .O(N__10639),
            .I(N__10627));
    InMux I__1705 (
            .O(N__10638),
            .I(N__10624));
    InMux I__1704 (
            .O(N__10637),
            .I(N__10621));
    InMux I__1703 (
            .O(N__10636),
            .I(N__10616));
    InMux I__1702 (
            .O(N__10633),
            .I(N__10616));
    InMux I__1701 (
            .O(N__10632),
            .I(N__10609));
    InMux I__1700 (
            .O(N__10631),
            .I(N__10609));
    InMux I__1699 (
            .O(N__10630),
            .I(N__10609));
    LocalMux I__1698 (
            .O(N__10627),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1697 (
            .O(N__10624),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1696 (
            .O(N__10621),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1695 (
            .O(N__10616),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1694 (
            .O(N__10609),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    CascadeMux I__1693 (
            .O(N__10598),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0_cascade_ ));
    InMux I__1692 (
            .O(N__10595),
            .I(N__10584));
    InMux I__1691 (
            .O(N__10594),
            .I(N__10581));
    InMux I__1690 (
            .O(N__10593),
            .I(N__10578));
    InMux I__1689 (
            .O(N__10592),
            .I(N__10575));
    InMux I__1688 (
            .O(N__10591),
            .I(N__10564));
    InMux I__1687 (
            .O(N__10590),
            .I(N__10564));
    InMux I__1686 (
            .O(N__10589),
            .I(N__10564));
    InMux I__1685 (
            .O(N__10588),
            .I(N__10564));
    InMux I__1684 (
            .O(N__10587),
            .I(N__10564));
    LocalMux I__1683 (
            .O(N__10584),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1682 (
            .O(N__10581),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1681 (
            .O(N__10578),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1680 (
            .O(N__10575),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1679 (
            .O(N__10564),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    InMux I__1678 (
            .O(N__10553),
            .I(N__10545));
    InMux I__1677 (
            .O(N__10552),
            .I(N__10536));
    InMux I__1676 (
            .O(N__10551),
            .I(N__10536));
    InMux I__1675 (
            .O(N__10550),
            .I(N__10536));
    InMux I__1674 (
            .O(N__10549),
            .I(N__10536));
    InMux I__1673 (
            .O(N__10548),
            .I(N__10531));
    LocalMux I__1672 (
            .O(N__10545),
            .I(N__10526));
    LocalMux I__1671 (
            .O(N__10536),
            .I(N__10526));
    InMux I__1670 (
            .O(N__10535),
            .I(N__10523));
    InMux I__1669 (
            .O(N__10534),
            .I(N__10520));
    LocalMux I__1668 (
            .O(N__10531),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1667 (
            .O(N__10526),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1666 (
            .O(N__10523),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1665 (
            .O(N__10520),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__1664 (
            .O(N__10511),
            .I(N__10502));
    InMux I__1663 (
            .O(N__10510),
            .I(N__10499));
    InMux I__1662 (
            .O(N__10509),
            .I(N__10494));
    InMux I__1661 (
            .O(N__10508),
            .I(N__10494));
    InMux I__1660 (
            .O(N__10507),
            .I(N__10487));
    InMux I__1659 (
            .O(N__10506),
            .I(N__10487));
    InMux I__1658 (
            .O(N__10505),
            .I(N__10487));
    LocalMux I__1657 (
            .O(N__10502),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1656 (
            .O(N__10499),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1655 (
            .O(N__10494),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1654 (
            .O(N__10487),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    CascadeMux I__1653 (
            .O(N__10478),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_ ));
    InMux I__1652 (
            .O(N__10475),
            .I(N__10469));
    InMux I__1651 (
            .O(N__10474),
            .I(N__10469));
    LocalMux I__1650 (
            .O(N__10469),
            .I(\this_vga_signals.mult1_un68_sum_c2_0 ));
    CEMux I__1649 (
            .O(N__10466),
            .I(N__10463));
    LocalMux I__1648 (
            .O(N__10463),
            .I(N__10460));
    Odrv4 I__1647 (
            .O(N__10460),
            .I(\this_vga_signals.N_469_1 ));
    IoInMux I__1646 (
            .O(N__10457),
            .I(N__10454));
    LocalMux I__1645 (
            .O(N__10454),
            .I(N__10451));
    IoSpan4Mux I__1644 (
            .O(N__10451),
            .I(N__10448));
    Span4Mux_s3_v I__1643 (
            .O(N__10448),
            .I(N__10445));
    Sp12to4 I__1642 (
            .O(N__10445),
            .I(N__10442));
    Span12Mux_v I__1641 (
            .O(N__10442),
            .I(N__10439));
    Odrv12 I__1640 (
            .O(N__10439),
            .I(debug_0_i));
    InMux I__1639 (
            .O(N__10436),
            .I(N__10433));
    LocalMux I__1638 (
            .O(N__10433),
            .I(N__10430));
    Span4Mux_h I__1637 (
            .O(N__10430),
            .I(N__10427));
    Span4Mux_h I__1636 (
            .O(N__10427),
            .I(N__10424));
    Odrv4 I__1635 (
            .O(N__10424),
            .I(\this_vga_signals.rgb_cnst_i_a5_0_0Z0Z_3 ));
    InMux I__1634 (
            .O(N__10421),
            .I(N__10417));
    InMux I__1633 (
            .O(N__10420),
            .I(N__10414));
    LocalMux I__1632 (
            .O(N__10417),
            .I(N__10405));
    LocalMux I__1631 (
            .O(N__10414),
            .I(N__10405));
    InMux I__1630 (
            .O(N__10413),
            .I(N__10402));
    InMux I__1629 (
            .O(N__10412),
            .I(N__10399));
    InMux I__1628 (
            .O(N__10411),
            .I(N__10396));
    CascadeMux I__1627 (
            .O(N__10410),
            .I(N__10393));
    Span4Mux_v I__1626 (
            .O(N__10405),
            .I(N__10387));
    LocalMux I__1625 (
            .O(N__10402),
            .I(N__10387));
    LocalMux I__1624 (
            .O(N__10399),
            .I(N__10382));
    LocalMux I__1623 (
            .O(N__10396),
            .I(N__10382));
    InMux I__1622 (
            .O(N__10393),
            .I(N__10377));
    InMux I__1621 (
            .O(N__10392),
            .I(N__10377));
    Span4Mux_h I__1620 (
            .O(N__10387),
            .I(N__10373));
    Span4Mux_v I__1619 (
            .O(N__10382),
            .I(N__10370));
    LocalMux I__1618 (
            .O(N__10377),
            .I(N__10367));
    InMux I__1617 (
            .O(N__10376),
            .I(N__10364));
    Span4Mux_h I__1616 (
            .O(N__10373),
            .I(N__10361));
    Span4Mux_h I__1615 (
            .O(N__10370),
            .I(N__10354));
    Span4Mux_v I__1614 (
            .O(N__10367),
            .I(N__10354));
    LocalMux I__1613 (
            .O(N__10364),
            .I(N__10354));
    Odrv4 I__1612 (
            .O(N__10361),
            .I(M_this_vram_read_data_0));
    Odrv4 I__1611 (
            .O(N__10354),
            .I(M_this_vram_read_data_0));
    CascadeMux I__1610 (
            .O(N__10349),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ));
    CascadeMux I__1609 (
            .O(N__10346),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1_cascade_ ));
    CascadeMux I__1608 (
            .O(N__10343),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_cascade_ ));
    InMux I__1607 (
            .O(N__10340),
            .I(N__10337));
    LocalMux I__1606 (
            .O(N__10337),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1 ));
    CascadeMux I__1605 (
            .O(N__10334),
            .I(N__10327));
    InMux I__1604 (
            .O(N__10333),
            .I(N__10318));
    InMux I__1603 (
            .O(N__10332),
            .I(N__10318));
    InMux I__1602 (
            .O(N__10331),
            .I(N__10318));
    InMux I__1601 (
            .O(N__10330),
            .I(N__10313));
    InMux I__1600 (
            .O(N__10327),
            .I(N__10313));
    CascadeMux I__1599 (
            .O(N__10326),
            .I(N__10310));
    InMux I__1598 (
            .O(N__10325),
            .I(N__10305));
    LocalMux I__1597 (
            .O(N__10318),
            .I(N__10300));
    LocalMux I__1596 (
            .O(N__10313),
            .I(N__10300));
    InMux I__1595 (
            .O(N__10310),
            .I(N__10293));
    InMux I__1594 (
            .O(N__10309),
            .I(N__10293));
    InMux I__1593 (
            .O(N__10308),
            .I(N__10293));
    LocalMux I__1592 (
            .O(N__10305),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1591 (
            .O(N__10300),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__1590 (
            .O(N__10293),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    CascadeMux I__1589 (
            .O(N__10286),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0_0_cascade_ ));
    InMux I__1588 (
            .O(N__10283),
            .I(N__10280));
    LocalMux I__1587 (
            .O(N__10280),
            .I(\this_vga_signals.if_N_9_0_0 ));
    InMux I__1586 (
            .O(N__10277),
            .I(N__10269));
    InMux I__1585 (
            .O(N__10276),
            .I(N__10269));
    InMux I__1584 (
            .O(N__10275),
            .I(N__10264));
    InMux I__1583 (
            .O(N__10274),
            .I(N__10264));
    LocalMux I__1582 (
            .O(N__10269),
            .I(\this_vga_signals.mult1_un68_sum_axb1 ));
    LocalMux I__1581 (
            .O(N__10264),
            .I(\this_vga_signals.mult1_un68_sum_axb1 ));
    CascadeMux I__1580 (
            .O(N__10259),
            .I(N__10256));
    CascadeBuf I__1579 (
            .O(N__10256),
            .I(N__10253));
    CascadeMux I__1578 (
            .O(N__10253),
            .I(N__10250));
    CascadeBuf I__1577 (
            .O(N__10250),
            .I(N__10247));
    CascadeMux I__1576 (
            .O(N__10247),
            .I(N__10244));
    CascadeBuf I__1575 (
            .O(N__10244),
            .I(N__10241));
    CascadeMux I__1574 (
            .O(N__10241),
            .I(N__10238));
    CascadeBuf I__1573 (
            .O(N__10238),
            .I(N__10235));
    CascadeMux I__1572 (
            .O(N__10235),
            .I(N__10232));
    CascadeBuf I__1571 (
            .O(N__10232),
            .I(N__10229));
    CascadeMux I__1570 (
            .O(N__10229),
            .I(N__10226));
    CascadeBuf I__1569 (
            .O(N__10226),
            .I(N__10223));
    CascadeMux I__1568 (
            .O(N__10223),
            .I(N__10220));
    CascadeBuf I__1567 (
            .O(N__10220),
            .I(N__10217));
    CascadeMux I__1566 (
            .O(N__10217),
            .I(N__10214));
    CascadeBuf I__1565 (
            .O(N__10214),
            .I(N__10211));
    CascadeMux I__1564 (
            .O(N__10211),
            .I(N__10208));
    CascadeBuf I__1563 (
            .O(N__10208),
            .I(N__10205));
    CascadeMux I__1562 (
            .O(N__10205),
            .I(N__10202));
    CascadeBuf I__1561 (
            .O(N__10202),
            .I(N__10199));
    CascadeMux I__1560 (
            .O(N__10199),
            .I(N__10196));
    CascadeBuf I__1559 (
            .O(N__10196),
            .I(N__10193));
    CascadeMux I__1558 (
            .O(N__10193),
            .I(N__10190));
    CascadeBuf I__1557 (
            .O(N__10190),
            .I(N__10187));
    CascadeMux I__1556 (
            .O(N__10187),
            .I(N__10184));
    CascadeBuf I__1555 (
            .O(N__10184),
            .I(N__10181));
    CascadeMux I__1554 (
            .O(N__10181),
            .I(N__10178));
    CascadeBuf I__1553 (
            .O(N__10178),
            .I(N__10175));
    CascadeMux I__1552 (
            .O(N__10175),
            .I(N__10172));
    CascadeBuf I__1551 (
            .O(N__10172),
            .I(N__10169));
    CascadeMux I__1550 (
            .O(N__10169),
            .I(N__10166));
    InMux I__1549 (
            .O(N__10166),
            .I(N__10163));
    LocalMux I__1548 (
            .O(N__10163),
            .I(N__10160));
    Span12Mux_s2_v I__1547 (
            .O(N__10160),
            .I(N__10157));
    Span12Mux_h I__1546 (
            .O(N__10157),
            .I(N__10154));
    Odrv12 I__1545 (
            .O(N__10154),
            .I(M_this_vga_signals_address_0));
    CascadeMux I__1544 (
            .O(N__10151),
            .I(\this_vga_signals.if_N_8_i_cascade_ ));
    InMux I__1543 (
            .O(N__10148),
            .I(N__10145));
    LocalMux I__1542 (
            .O(N__10145),
            .I(\this_vga_signals.mult1_un82_sum_axb1 ));
    InMux I__1541 (
            .O(N__10142),
            .I(N__10139));
    LocalMux I__1540 (
            .O(N__10139),
            .I(\this_vga_signals.mult1_un89_sum_c3 ));
    CascadeMux I__1539 (
            .O(N__10136),
            .I(\this_vga_signals.mult1_un82_sum_c3_cascade_ ));
    CascadeMux I__1538 (
            .O(N__10133),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_ ));
    InMux I__1537 (
            .O(N__10130),
            .I(N__10127));
    LocalMux I__1536 (
            .O(N__10127),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_2 ));
    InMux I__1535 (
            .O(N__10124),
            .I(N__10121));
    LocalMux I__1534 (
            .O(N__10121),
            .I(\this_vga_signals.mult1_un82_sum_c2_0 ));
    InMux I__1533 (
            .O(N__10118),
            .I(N__10115));
    LocalMux I__1532 (
            .O(N__10115),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0 ));
    InMux I__1531 (
            .O(N__10112),
            .I(N__10109));
    LocalMux I__1530 (
            .O(N__10109),
            .I(\this_vga_signals.g0_i_x2_5 ));
    CascadeMux I__1529 (
            .O(N__10106),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_cascade_ ));
    InMux I__1528 (
            .O(N__10103),
            .I(N__10100));
    LocalMux I__1527 (
            .O(N__10100),
            .I(\this_vga_signals.N_9_1_0 ));
    CascadeMux I__1526 (
            .O(N__10097),
            .I(N__10094));
    InMux I__1525 (
            .O(N__10094),
            .I(N__10091));
    LocalMux I__1524 (
            .O(N__10091),
            .I(N__10088));
    Odrv4 I__1523 (
            .O(N__10088),
            .I(\this_vga_signals.g1_5 ));
    InMux I__1522 (
            .O(N__10085),
            .I(N__10082));
    LocalMux I__1521 (
            .O(N__10082),
            .I(\this_vga_signals.N_6 ));
    CascadeMux I__1520 (
            .O(N__10079),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_0_0_1_cascade_ ));
    CascadeMux I__1519 (
            .O(N__10076),
            .I(N__10073));
    CascadeBuf I__1518 (
            .O(N__10073),
            .I(N__10070));
    CascadeMux I__1517 (
            .O(N__10070),
            .I(N__10067));
    CascadeBuf I__1516 (
            .O(N__10067),
            .I(N__10064));
    CascadeMux I__1515 (
            .O(N__10064),
            .I(N__10061));
    CascadeBuf I__1514 (
            .O(N__10061),
            .I(N__10058));
    CascadeMux I__1513 (
            .O(N__10058),
            .I(N__10055));
    CascadeBuf I__1512 (
            .O(N__10055),
            .I(N__10052));
    CascadeMux I__1511 (
            .O(N__10052),
            .I(N__10049));
    CascadeBuf I__1510 (
            .O(N__10049),
            .I(N__10046));
    CascadeMux I__1509 (
            .O(N__10046),
            .I(N__10043));
    CascadeBuf I__1508 (
            .O(N__10043),
            .I(N__10040));
    CascadeMux I__1507 (
            .O(N__10040),
            .I(N__10037));
    CascadeBuf I__1506 (
            .O(N__10037),
            .I(N__10034));
    CascadeMux I__1505 (
            .O(N__10034),
            .I(N__10031));
    CascadeBuf I__1504 (
            .O(N__10031),
            .I(N__10028));
    CascadeMux I__1503 (
            .O(N__10028),
            .I(N__10025));
    CascadeBuf I__1502 (
            .O(N__10025),
            .I(N__10022));
    CascadeMux I__1501 (
            .O(N__10022),
            .I(N__10019));
    CascadeBuf I__1500 (
            .O(N__10019),
            .I(N__10016));
    CascadeMux I__1499 (
            .O(N__10016),
            .I(N__10013));
    CascadeBuf I__1498 (
            .O(N__10013),
            .I(N__10010));
    CascadeMux I__1497 (
            .O(N__10010),
            .I(N__10007));
    CascadeBuf I__1496 (
            .O(N__10007),
            .I(N__10004));
    CascadeMux I__1495 (
            .O(N__10004),
            .I(N__10001));
    CascadeBuf I__1494 (
            .O(N__10001),
            .I(N__9998));
    CascadeMux I__1493 (
            .O(N__9998),
            .I(N__9995));
    CascadeBuf I__1492 (
            .O(N__9995),
            .I(N__9992));
    CascadeMux I__1491 (
            .O(N__9992),
            .I(N__9989));
    CascadeBuf I__1490 (
            .O(N__9989),
            .I(N__9986));
    CascadeMux I__1489 (
            .O(N__9986),
            .I(N__9983));
    InMux I__1488 (
            .O(N__9983),
            .I(N__9980));
    LocalMux I__1487 (
            .O(N__9980),
            .I(N__9977));
    Span4Mux_v I__1486 (
            .O(N__9977),
            .I(N__9974));
    Span4Mux_v I__1485 (
            .O(N__9974),
            .I(N__9971));
    Span4Mux_v I__1484 (
            .O(N__9971),
            .I(N__9968));
    Span4Mux_h I__1483 (
            .O(N__9968),
            .I(N__9965));
    Span4Mux_h I__1482 (
            .O(N__9965),
            .I(N__9962));
    Odrv4 I__1481 (
            .O(N__9962),
            .I(M_this_vga_signals_address_7));
    InMux I__1480 (
            .O(N__9959),
            .I(N__9956));
    LocalMux I__1479 (
            .O(N__9956),
            .I(\this_vga_signals.g2_0_1_0 ));
    InMux I__1478 (
            .O(N__9953),
            .I(N__9950));
    LocalMux I__1477 (
            .O(N__9950),
            .I(\this_vga_signals.g0_i_x2_2 ));
    CascadeMux I__1476 (
            .O(N__9947),
            .I(\this_vga_signals.g0_i_0_N_4L5_cascade_ ));
    InMux I__1475 (
            .O(N__9944),
            .I(N__9941));
    LocalMux I__1474 (
            .O(N__9941),
            .I(\this_vga_signals.g0_i_0_N_5L7 ));
    InMux I__1473 (
            .O(N__9938),
            .I(N__9935));
    LocalMux I__1472 (
            .O(N__9935),
            .I(\this_vga_signals.if_i4_mux_0_0_0_1 ));
    InMux I__1471 (
            .O(N__9932),
            .I(N__9929));
    LocalMux I__1470 (
            .O(N__9929),
            .I(\this_vga_signals.N_6_i ));
    CascadeMux I__1469 (
            .O(N__9926),
            .I(N__9923));
    InMux I__1468 (
            .O(N__9923),
            .I(N__9920));
    LocalMux I__1467 (
            .O(N__9920),
            .I(N__9917));
    Span4Mux_v I__1466 (
            .O(N__9917),
            .I(N__9914));
    Odrv4 I__1465 (
            .O(N__9914),
            .I(\this_vga_signals.g1_1_2 ));
    InMux I__1464 (
            .O(N__9911),
            .I(N__9908));
    LocalMux I__1463 (
            .O(N__9908),
            .I(\this_vga_signals.g1_4_1 ));
    InMux I__1462 (
            .O(N__9905),
            .I(N__9902));
    LocalMux I__1461 (
            .O(N__9902),
            .I(N__9898));
    InMux I__1460 (
            .O(N__9901),
            .I(N__9894));
    Span4Mux_h I__1459 (
            .O(N__9898),
            .I(N__9891));
    InMux I__1458 (
            .O(N__9897),
            .I(N__9888));
    LocalMux I__1457 (
            .O(N__9894),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__1456 (
            .O(N__9891),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__1455 (
            .O(N__9888),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    InMux I__1454 (
            .O(N__9881),
            .I(N__9878));
    LocalMux I__1453 (
            .O(N__9878),
            .I(\this_vga_signals.g0_i_0_N_2L1 ));
    InMux I__1452 (
            .O(N__9875),
            .I(N__9868));
    InMux I__1451 (
            .O(N__9874),
            .I(N__9868));
    CascadeMux I__1450 (
            .O(N__9873),
            .I(N__9864));
    LocalMux I__1449 (
            .O(N__9868),
            .I(N__9856));
    InMux I__1448 (
            .O(N__9867),
            .I(N__9853));
    InMux I__1447 (
            .O(N__9864),
            .I(N__9849));
    InMux I__1446 (
            .O(N__9863),
            .I(N__9844));
    InMux I__1445 (
            .O(N__9862),
            .I(N__9844));
    InMux I__1444 (
            .O(N__9861),
            .I(N__9841));
    InMux I__1443 (
            .O(N__9860),
            .I(N__9836));
    InMux I__1442 (
            .O(N__9859),
            .I(N__9836));
    Span4Mux_v I__1441 (
            .O(N__9856),
            .I(N__9825));
    LocalMux I__1440 (
            .O(N__9853),
            .I(N__9825));
    InMux I__1439 (
            .O(N__9852),
            .I(N__9822));
    LocalMux I__1438 (
            .O(N__9849),
            .I(N__9814));
    LocalMux I__1437 (
            .O(N__9844),
            .I(N__9814));
    LocalMux I__1436 (
            .O(N__9841),
            .I(N__9814));
    LocalMux I__1435 (
            .O(N__9836),
            .I(N__9811));
    InMux I__1434 (
            .O(N__9835),
            .I(N__9808));
    InMux I__1433 (
            .O(N__9834),
            .I(N__9801));
    InMux I__1432 (
            .O(N__9833),
            .I(N__9801));
    InMux I__1431 (
            .O(N__9832),
            .I(N__9801));
    InMux I__1430 (
            .O(N__9831),
            .I(N__9796));
    InMux I__1429 (
            .O(N__9830),
            .I(N__9796));
    Span4Mux_h I__1428 (
            .O(N__9825),
            .I(N__9785));
    LocalMux I__1427 (
            .O(N__9822),
            .I(N__9785));
    InMux I__1426 (
            .O(N__9821),
            .I(N__9782));
    Span4Mux_v I__1425 (
            .O(N__9814),
            .I(N__9775));
    Span4Mux_v I__1424 (
            .O(N__9811),
            .I(N__9775));
    LocalMux I__1423 (
            .O(N__9808),
            .I(N__9775));
    LocalMux I__1422 (
            .O(N__9801),
            .I(N__9770));
    LocalMux I__1421 (
            .O(N__9796),
            .I(N__9770));
    InMux I__1420 (
            .O(N__9795),
            .I(N__9763));
    InMux I__1419 (
            .O(N__9794),
            .I(N__9763));
    InMux I__1418 (
            .O(N__9793),
            .I(N__9763));
    InMux I__1417 (
            .O(N__9792),
            .I(N__9756));
    InMux I__1416 (
            .O(N__9791),
            .I(N__9756));
    InMux I__1415 (
            .O(N__9790),
            .I(N__9756));
    Odrv4 I__1414 (
            .O(N__9785),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__1413 (
            .O(N__9782),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__1412 (
            .O(N__9775),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__1411 (
            .O(N__9770),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__1410 (
            .O(N__9763),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__1409 (
            .O(N__9756),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__1408 (
            .O(N__9743),
            .I(N__9736));
    InMux I__1407 (
            .O(N__9742),
            .I(N__9733));
    InMux I__1406 (
            .O(N__9741),
            .I(N__9729));
    InMux I__1405 (
            .O(N__9740),
            .I(N__9722));
    InMux I__1404 (
            .O(N__9739),
            .I(N__9722));
    LocalMux I__1403 (
            .O(N__9736),
            .I(N__9718));
    LocalMux I__1402 (
            .O(N__9733),
            .I(N__9715));
    InMux I__1401 (
            .O(N__9732),
            .I(N__9712));
    LocalMux I__1400 (
            .O(N__9729),
            .I(N__9706));
    InMux I__1399 (
            .O(N__9728),
            .I(N__9701));
    InMux I__1398 (
            .O(N__9727),
            .I(N__9701));
    LocalMux I__1397 (
            .O(N__9722),
            .I(N__9698));
    InMux I__1396 (
            .O(N__9721),
            .I(N__9694));
    Span4Mux_h I__1395 (
            .O(N__9718),
            .I(N__9691));
    Span4Mux_h I__1394 (
            .O(N__9715),
            .I(N__9688));
    LocalMux I__1393 (
            .O(N__9712),
            .I(N__9685));
    InMux I__1392 (
            .O(N__9711),
            .I(N__9680));
    InMux I__1391 (
            .O(N__9710),
            .I(N__9680));
    InMux I__1390 (
            .O(N__9709),
            .I(N__9677));
    Span4Mux_h I__1389 (
            .O(N__9706),
            .I(N__9670));
    LocalMux I__1388 (
            .O(N__9701),
            .I(N__9670));
    Span4Mux_h I__1387 (
            .O(N__9698),
            .I(N__9670));
    InMux I__1386 (
            .O(N__9697),
            .I(N__9667));
    LocalMux I__1385 (
            .O(N__9694),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__1384 (
            .O(N__9691),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__1383 (
            .O(N__9688),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv12 I__1382 (
            .O(N__9685),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__1381 (
            .O(N__9680),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__1380 (
            .O(N__9677),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__1379 (
            .O(N__9670),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__1378 (
            .O(N__9667),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    InMux I__1377 (
            .O(N__9650),
            .I(N__9647));
    LocalMux I__1376 (
            .O(N__9647),
            .I(N__9644));
    Span4Mux_v I__1375 (
            .O(N__9644),
            .I(N__9641));
    Odrv4 I__1374 (
            .O(N__9641),
            .I(\this_vga_signals.M_vcounter_d_1_sqmuxa_i_a3_1 ));
    InMux I__1373 (
            .O(N__9638),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__1372 (
            .O(N__9635),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__1371 (
            .O(N__9632),
            .I(bfn_12_25_0_));
    InMux I__1370 (
            .O(N__9629),
            .I(N__9626));
    LocalMux I__1369 (
            .O(N__9626),
            .I(N__9623));
    Odrv4 I__1368 (
            .O(N__9623),
            .I(\this_vga_signals.N_22 ));
    CascadeMux I__1367 (
            .O(N__9620),
            .I(\this_vga_signals.g1_0_0_2_cascade_ ));
    InMux I__1366 (
            .O(N__9617),
            .I(N__9614));
    LocalMux I__1365 (
            .O(N__9614),
            .I(\this_vga_signals.N_21 ));
    InMux I__1364 (
            .O(N__9611),
            .I(N__9608));
    LocalMux I__1363 (
            .O(N__9608),
            .I(N__9605));
    Odrv12 I__1362 (
            .O(N__9605),
            .I(\this_vga_signals.g0_i_x2_1 ));
    InMux I__1361 (
            .O(N__9602),
            .I(N__9599));
    LocalMux I__1360 (
            .O(N__9599),
            .I(\this_vga_signals.g4_1 ));
    CascadeMux I__1359 (
            .O(N__9596),
            .I(\this_vga_signals.g0_1_0_cascade_ ));
    InMux I__1358 (
            .O(N__9593),
            .I(N__9590));
    LocalMux I__1357 (
            .O(N__9590),
            .I(N__9586));
    InMux I__1356 (
            .O(N__9589),
            .I(N__9583));
    Odrv12 I__1355 (
            .O(N__9586),
            .I(\this_vga_signals.CO0_i_i ));
    LocalMux I__1354 (
            .O(N__9583),
            .I(\this_vga_signals.CO0_i_i ));
    CascadeMux I__1353 (
            .O(N__9578),
            .I(\this_vga_signals.N_45_cascade_ ));
    CascadeMux I__1352 (
            .O(N__9575),
            .I(N__9571));
    InMux I__1351 (
            .O(N__9574),
            .I(N__9567));
    InMux I__1350 (
            .O(N__9571),
            .I(N__9564));
    InMux I__1349 (
            .O(N__9570),
            .I(N__9561));
    LocalMux I__1348 (
            .O(N__9567),
            .I(N_23_0));
    LocalMux I__1347 (
            .O(N__9564),
            .I(N_23_0));
    LocalMux I__1346 (
            .O(N__9561),
            .I(N_23_0));
    CascadeMux I__1345 (
            .O(N__9554),
            .I(N_23_0_cascade_));
    InMux I__1344 (
            .O(N__9551),
            .I(N__9546));
    InMux I__1343 (
            .O(N__9550),
            .I(N__9541));
    InMux I__1342 (
            .O(N__9549),
            .I(N__9541));
    LocalMux I__1341 (
            .O(N__9546),
            .I(\this_pixel_clock.M_counter_q_i_1 ));
    LocalMux I__1340 (
            .O(N__9541),
            .I(\this_pixel_clock.M_counter_q_i_1 ));
    InMux I__1339 (
            .O(N__9536),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__1338 (
            .O(N__9533),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__1337 (
            .O(N__9530),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__1336 (
            .O(N__9527),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__1335 (
            .O(N__9524),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    CascadeMux I__1334 (
            .O(N__9521),
            .I(\this_vga_signals.N_28_0_cascade_ ));
    CascadeMux I__1333 (
            .O(N__9518),
            .I(\this_vga_signals.N_42_cascade_ ));
    IoInMux I__1332 (
            .O(N__9515),
            .I(N__9512));
    LocalMux I__1331 (
            .O(N__9512),
            .I(N__9509));
    Span4Mux_s2_v I__1330 (
            .O(N__9509),
            .I(N__9506));
    Span4Mux_v I__1329 (
            .O(N__9506),
            .I(N__9503));
    Span4Mux_v I__1328 (
            .O(N__9503),
            .I(N__9500));
    Odrv4 I__1327 (
            .O(N__9500),
            .I(\this_vga_signals.M_vcounter_q_esr_RNIVV6F6Z0Z_9 ));
    InMux I__1326 (
            .O(N__9497),
            .I(N__9492));
    InMux I__1325 (
            .O(N__9496),
            .I(N__9489));
    InMux I__1324 (
            .O(N__9495),
            .I(N__9486));
    LocalMux I__1323 (
            .O(N__9492),
            .I(N__9481));
    LocalMux I__1322 (
            .O(N__9489),
            .I(N__9476));
    LocalMux I__1321 (
            .O(N__9486),
            .I(N__9476));
    CascadeMux I__1320 (
            .O(N__9485),
            .I(N__9466));
    CascadeMux I__1319 (
            .O(N__9484),
            .I(N__9462));
    Span4Mux_v I__1318 (
            .O(N__9481),
            .I(N__9459));
    Span4Mux_h I__1317 (
            .O(N__9476),
            .I(N__9456));
    InMux I__1316 (
            .O(N__9475),
            .I(N__9453));
    InMux I__1315 (
            .O(N__9474),
            .I(N__9448));
    InMux I__1314 (
            .O(N__9473),
            .I(N__9448));
    InMux I__1313 (
            .O(N__9472),
            .I(N__9445));
    InMux I__1312 (
            .O(N__9471),
            .I(N__9440));
    InMux I__1311 (
            .O(N__9470),
            .I(N__9440));
    InMux I__1310 (
            .O(N__9469),
            .I(N__9435));
    InMux I__1309 (
            .O(N__9466),
            .I(N__9435));
    InMux I__1308 (
            .O(N__9465),
            .I(N__9430));
    InMux I__1307 (
            .O(N__9462),
            .I(N__9430));
    Odrv4 I__1306 (
            .O(N__9459),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__1305 (
            .O(N__9456),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__1304 (
            .O(N__9453),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__1303 (
            .O(N__9448),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__1302 (
            .O(N__9445),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__1301 (
            .O(N__9440),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__1300 (
            .O(N__9435),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__1299 (
            .O(N__9430),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    CascadeMux I__1298 (
            .O(N__9413),
            .I(\this_vga_signals.rgb297_i_a3_0_cascade_ ));
    CascadeMux I__1297 (
            .O(N__9410),
            .I(N__9407));
    InMux I__1296 (
            .O(N__9407),
            .I(N__9399));
    InMux I__1295 (
            .O(N__9406),
            .I(N__9396));
    InMux I__1294 (
            .O(N__9405),
            .I(N__9393));
    InMux I__1293 (
            .O(N__9404),
            .I(N__9385));
    InMux I__1292 (
            .O(N__9403),
            .I(N__9385));
    CascadeMux I__1291 (
            .O(N__9402),
            .I(N__9382));
    LocalMux I__1290 (
            .O(N__9399),
            .I(N__9375));
    LocalMux I__1289 (
            .O(N__9396),
            .I(N__9372));
    LocalMux I__1288 (
            .O(N__9393),
            .I(N__9369));
    CascadeMux I__1287 (
            .O(N__9392),
            .I(N__9366));
    CascadeMux I__1286 (
            .O(N__9391),
            .I(N__9361));
    InMux I__1285 (
            .O(N__9390),
            .I(N__9354));
    LocalMux I__1284 (
            .O(N__9385),
            .I(N__9351));
    InMux I__1283 (
            .O(N__9382),
            .I(N__9344));
    InMux I__1282 (
            .O(N__9381),
            .I(N__9344));
    InMux I__1281 (
            .O(N__9380),
            .I(N__9344));
    InMux I__1280 (
            .O(N__9379),
            .I(N__9339));
    InMux I__1279 (
            .O(N__9378),
            .I(N__9339));
    Span4Mux_v I__1278 (
            .O(N__9375),
            .I(N__9336));
    Span4Mux_h I__1277 (
            .O(N__9372),
            .I(N__9331));
    Span4Mux_h I__1276 (
            .O(N__9369),
            .I(N__9331));
    InMux I__1275 (
            .O(N__9366),
            .I(N__9324));
    InMux I__1274 (
            .O(N__9365),
            .I(N__9324));
    InMux I__1273 (
            .O(N__9364),
            .I(N__9324));
    InMux I__1272 (
            .O(N__9361),
            .I(N__9321));
    InMux I__1271 (
            .O(N__9360),
            .I(N__9312));
    InMux I__1270 (
            .O(N__9359),
            .I(N__9312));
    InMux I__1269 (
            .O(N__9358),
            .I(N__9312));
    InMux I__1268 (
            .O(N__9357),
            .I(N__9312));
    LocalMux I__1267 (
            .O(N__9354),
            .I(N__9309));
    Span4Mux_h I__1266 (
            .O(N__9351),
            .I(N__9302));
    LocalMux I__1265 (
            .O(N__9344),
            .I(N__9302));
    LocalMux I__1264 (
            .O(N__9339),
            .I(N__9302));
    Odrv4 I__1263 (
            .O(N__9336),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__1262 (
            .O(N__9331),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__1261 (
            .O(N__9324),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__1260 (
            .O(N__9321),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__1259 (
            .O(N__9312),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__1258 (
            .O(N__9309),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__1257 (
            .O(N__9302),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    InMux I__1256 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__1255 (
            .O(N__9284),
            .I(\this_vga_signals.SUM_2_i_a4_0_a0_2_3 ));
    InMux I__1254 (
            .O(N__9281),
            .I(N__9278));
    LocalMux I__1253 (
            .O(N__9278),
            .I(N__9275));
    Span4Mux_v I__1252 (
            .O(N__9275),
            .I(N__9272));
    Span4Mux_h I__1251 (
            .O(N__9272),
            .I(N__9269));
    Span4Mux_h I__1250 (
            .O(N__9269),
            .I(N__9266));
    Odrv4 I__1249 (
            .O(N__9266),
            .I(\this_vga_signals.N_33_0 ));
    InMux I__1248 (
            .O(N__9263),
            .I(N__9254));
    InMux I__1247 (
            .O(N__9262),
            .I(N__9251));
    InMux I__1246 (
            .O(N__9261),
            .I(N__9247));
    InMux I__1245 (
            .O(N__9260),
            .I(N__9244));
    InMux I__1244 (
            .O(N__9259),
            .I(N__9241));
    InMux I__1243 (
            .O(N__9258),
            .I(N__9236));
    InMux I__1242 (
            .O(N__9257),
            .I(N__9236));
    LocalMux I__1241 (
            .O(N__9254),
            .I(N__9233));
    LocalMux I__1240 (
            .O(N__9251),
            .I(N__9230));
    CascadeMux I__1239 (
            .O(N__9250),
            .I(N__9224));
    LocalMux I__1238 (
            .O(N__9247),
            .I(N__9220));
    LocalMux I__1237 (
            .O(N__9244),
            .I(N__9217));
    LocalMux I__1236 (
            .O(N__9241),
            .I(N__9212));
    LocalMux I__1235 (
            .O(N__9236),
            .I(N__9212));
    Span4Mux_h I__1234 (
            .O(N__9233),
            .I(N__9208));
    Span4Mux_h I__1233 (
            .O(N__9230),
            .I(N__9205));
    InMux I__1232 (
            .O(N__9229),
            .I(N__9200));
    InMux I__1231 (
            .O(N__9228),
            .I(N__9200));
    InMux I__1230 (
            .O(N__9227),
            .I(N__9197));
    InMux I__1229 (
            .O(N__9224),
            .I(N__9192));
    InMux I__1228 (
            .O(N__9223),
            .I(N__9192));
    Span4Mux_v I__1227 (
            .O(N__9220),
            .I(N__9185));
    Span4Mux_v I__1226 (
            .O(N__9217),
            .I(N__9185));
    Span4Mux_v I__1225 (
            .O(N__9212),
            .I(N__9185));
    InMux I__1224 (
            .O(N__9211),
            .I(N__9182));
    Odrv4 I__1223 (
            .O(N__9208),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__1222 (
            .O(N__9205),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__1221 (
            .O(N__9200),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__1220 (
            .O(N__9197),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__1219 (
            .O(N__9192),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__1218 (
            .O(N__9185),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__1217 (
            .O(N__9182),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    InMux I__1216 (
            .O(N__9167),
            .I(N__9164));
    LocalMux I__1215 (
            .O(N__9164),
            .I(N__9160));
    InMux I__1214 (
            .O(N__9163),
            .I(N__9157));
    Odrv12 I__1213 (
            .O(N__9160),
            .I(\this_vga_signals.N_49 ));
    LocalMux I__1212 (
            .O(N__9157),
            .I(\this_vga_signals.N_49 ));
    CascadeMux I__1211 (
            .O(N__9152),
            .I(\this_vga_signals.N_33_0_cascade_ ));
    InMux I__1210 (
            .O(N__9149),
            .I(N__9146));
    LocalMux I__1209 (
            .O(N__9146),
            .I(\this_vga_signals.N_11_i ));
    InMux I__1208 (
            .O(N__9143),
            .I(N__9139));
    InMux I__1207 (
            .O(N__9142),
            .I(N__9132));
    LocalMux I__1206 (
            .O(N__9139),
            .I(N__9129));
    InMux I__1205 (
            .O(N__9138),
            .I(N__9122));
    InMux I__1204 (
            .O(N__9137),
            .I(N__9122));
    InMux I__1203 (
            .O(N__9136),
            .I(N__9122));
    InMux I__1202 (
            .O(N__9135),
            .I(N__9119));
    LocalMux I__1201 (
            .O(N__9132),
            .I(\this_vga_signals.mult1_un40_sum_axb1 ));
    Odrv4 I__1200 (
            .O(N__9129),
            .I(\this_vga_signals.mult1_un40_sum_axb1 ));
    LocalMux I__1199 (
            .O(N__9122),
            .I(\this_vga_signals.mult1_un40_sum_axb1 ));
    LocalMux I__1198 (
            .O(N__9119),
            .I(\this_vga_signals.mult1_un40_sum_axb1 ));
    CascadeMux I__1197 (
            .O(N__9110),
            .I(N__9107));
    InMux I__1196 (
            .O(N__9107),
            .I(N__9104));
    LocalMux I__1195 (
            .O(N__9104),
            .I(\this_vga_signals.g0_5_0_0 ));
    InMux I__1194 (
            .O(N__9101),
            .I(N__9098));
    LocalMux I__1193 (
            .O(N__9098),
            .I(\this_vga_signals.mult1_un54_sum_axb1_5_4 ));
    CascadeMux I__1192 (
            .O(N__9095),
            .I(\this_vga_signals.g0_25_1_cascade_ ));
    InMux I__1191 (
            .O(N__9092),
            .I(N__9086));
    InMux I__1190 (
            .O(N__9091),
            .I(N__9083));
    InMux I__1189 (
            .O(N__9090),
            .I(N__9078));
    InMux I__1188 (
            .O(N__9089),
            .I(N__9078));
    LocalMux I__1187 (
            .O(N__9086),
            .I(N__9075));
    LocalMux I__1186 (
            .O(N__9083),
            .I(N__9072));
    LocalMux I__1185 (
            .O(N__9078),
            .I(N__9069));
    Span4Mux_v I__1184 (
            .O(N__9075),
            .I(N__9066));
    Span4Mux_h I__1183 (
            .O(N__9072),
            .I(N__9063));
    Span4Mux_h I__1182 (
            .O(N__9069),
            .I(N__9060));
    Odrv4 I__1181 (
            .O(N__9066),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c ));
    Odrv4 I__1180 (
            .O(N__9063),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c ));
    Odrv4 I__1179 (
            .O(N__9060),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c ));
    CascadeMux I__1178 (
            .O(N__9053),
            .I(\this_vga_signals.if_N_13_i_i_1_0_0_cascade_ ));
    InMux I__1177 (
            .O(N__9050),
            .I(N__9047));
    LocalMux I__1176 (
            .O(N__9047),
            .I(\this_vga_signals.g2_0_0_0 ));
    InMux I__1175 (
            .O(N__9044),
            .I(N__9041));
    LocalMux I__1174 (
            .O(N__9041),
            .I(N__9038));
    Span4Mux_v I__1173 (
            .O(N__9038),
            .I(N__9035));
    Odrv4 I__1172 (
            .O(N__9035),
            .I(\this_vga_signals.N_371_0 ));
    IoInMux I__1171 (
            .O(N__9032),
            .I(N__9029));
    LocalMux I__1170 (
            .O(N__9029),
            .I(N__9026));
    Span12Mux_s11_h I__1169 (
            .O(N__9026),
            .I(N__9023));
    Odrv12 I__1168 (
            .O(N__9023),
            .I(rgb_c_4));
    CascadeMux I__1167 (
            .O(N__9020),
            .I(N__9007));
    InMux I__1166 (
            .O(N__9019),
            .I(N__9004));
    CascadeMux I__1165 (
            .O(N__9018),
            .I(N__9001));
    CascadeMux I__1164 (
            .O(N__9017),
            .I(N__8997));
    CascadeMux I__1163 (
            .O(N__9016),
            .I(N__8994));
    CascadeMux I__1162 (
            .O(N__9015),
            .I(N__8991));
    InMux I__1161 (
            .O(N__9014),
            .I(N__8987));
    InMux I__1160 (
            .O(N__9013),
            .I(N__8983));
    InMux I__1159 (
            .O(N__9012),
            .I(N__8980));
    InMux I__1158 (
            .O(N__9011),
            .I(N__8975));
    InMux I__1157 (
            .O(N__9010),
            .I(N__8975));
    InMux I__1156 (
            .O(N__9007),
            .I(N__8972));
    LocalMux I__1155 (
            .O(N__9004),
            .I(N__8969));
    InMux I__1154 (
            .O(N__9001),
            .I(N__8962));
    InMux I__1153 (
            .O(N__9000),
            .I(N__8962));
    InMux I__1152 (
            .O(N__8997),
            .I(N__8962));
    InMux I__1151 (
            .O(N__8994),
            .I(N__8957));
    InMux I__1150 (
            .O(N__8991),
            .I(N__8957));
    InMux I__1149 (
            .O(N__8990),
            .I(N__8954));
    LocalMux I__1148 (
            .O(N__8987),
            .I(N__8951));
    InMux I__1147 (
            .O(N__8986),
            .I(N__8948));
    LocalMux I__1146 (
            .O(N__8983),
            .I(N__8945));
    LocalMux I__1145 (
            .O(N__8980),
            .I(N__8936));
    LocalMux I__1144 (
            .O(N__8975),
            .I(N__8936));
    LocalMux I__1143 (
            .O(N__8972),
            .I(N__8936));
    Span4Mux_h I__1142 (
            .O(N__8969),
            .I(N__8929));
    LocalMux I__1141 (
            .O(N__8962),
            .I(N__8929));
    LocalMux I__1140 (
            .O(N__8957),
            .I(N__8929));
    LocalMux I__1139 (
            .O(N__8954),
            .I(N__8926));
    Span4Mux_h I__1138 (
            .O(N__8951),
            .I(N__8919));
    LocalMux I__1137 (
            .O(N__8948),
            .I(N__8919));
    Span4Mux_v I__1136 (
            .O(N__8945),
            .I(N__8919));
    InMux I__1135 (
            .O(N__8944),
            .I(N__8914));
    InMux I__1134 (
            .O(N__8943),
            .I(N__8914));
    Span4Mux_h I__1133 (
            .O(N__8936),
            .I(N__8911));
    Span4Mux_v I__1132 (
            .O(N__8929),
            .I(N__8908));
    Odrv4 I__1131 (
            .O(N__8926),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0 ));
    Odrv4 I__1130 (
            .O(N__8919),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0 ));
    LocalMux I__1129 (
            .O(N__8914),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0 ));
    Odrv4 I__1128 (
            .O(N__8911),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0 ));
    Odrv4 I__1127 (
            .O(N__8908),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0 ));
    CascadeMux I__1126 (
            .O(N__8897),
            .I(\this_vga_signals.un11_address_0_7_cascade_ ));
    InMux I__1125 (
            .O(N__8894),
            .I(N__8888));
    InMux I__1124 (
            .O(N__8893),
            .I(N__8885));
    InMux I__1123 (
            .O(N__8892),
            .I(N__8880));
    InMux I__1122 (
            .O(N__8891),
            .I(N__8880));
    LocalMux I__1121 (
            .O(N__8888),
            .I(N__8877));
    LocalMux I__1120 (
            .O(N__8885),
            .I(\this_vga_signals.SUM_2 ));
    LocalMux I__1119 (
            .O(N__8880),
            .I(\this_vga_signals.SUM_2 ));
    Odrv4 I__1118 (
            .O(N__8877),
            .I(\this_vga_signals.SUM_2 ));
    InMux I__1117 (
            .O(N__8870),
            .I(N__8867));
    LocalMux I__1116 (
            .O(N__8867),
            .I(N__8864));
    Odrv4 I__1115 (
            .O(N__8864),
            .I(\this_vga_signals.g0_3_0 ));
    CascadeMux I__1114 (
            .O(N__8861),
            .I(this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_cascade_));
    InMux I__1113 (
            .O(N__8858),
            .I(N__8855));
    LocalMux I__1112 (
            .O(N__8855),
            .I(\this_vga_signals.g0_i_x2_1_1 ));
    InMux I__1111 (
            .O(N__8852),
            .I(N__8849));
    LocalMux I__1110 (
            .O(N__8849),
            .I(\this_vga_signals.g0_i_x1 ));
    CascadeMux I__1109 (
            .O(N__8846),
            .I(\this_vga_signals.g0_i_x0_cascade_ ));
    CascadeMux I__1108 (
            .O(N__8843),
            .I(this_vga_signals_un16_address_if_i1_mux_0_cascade_));
    CascadeMux I__1107 (
            .O(N__8840),
            .I(\this_vga_signals.N_6_i_cascade_ ));
    InMux I__1106 (
            .O(N__8837),
            .I(N__8834));
    LocalMux I__1105 (
            .O(N__8834),
            .I(\this_vga_signals.g1_1_0 ));
    CascadeMux I__1104 (
            .O(N__8831),
            .I(\this_vga_signals.M_vcounter_q_esr_RNIO6OD01Z0Z_9_cascade_ ));
    IoInMux I__1103 (
            .O(N__8828),
            .I(N__8825));
    LocalMux I__1102 (
            .O(N__8825),
            .I(N__8822));
    Span12Mux_s5_h I__1101 (
            .O(N__8822),
            .I(N__8819));
    Odrv12 I__1100 (
            .O(N__8819),
            .I(rgb_c_2));
    CascadeMux I__1099 (
            .O(N__8816),
            .I(N__8813));
    InMux I__1098 (
            .O(N__8813),
            .I(N__8810));
    LocalMux I__1097 (
            .O(N__8810),
            .I(N__8807));
    Odrv12 I__1096 (
            .O(N__8807),
            .I(\this_vga_signals.g0_i_x2_1_0 ));
    InMux I__1095 (
            .O(N__8804),
            .I(N__8801));
    LocalMux I__1094 (
            .O(N__8801),
            .I(\this_vga_signals.N_10_i ));
    CascadeMux I__1093 (
            .O(N__8798),
            .I(\this_vga_signals.N_10_i_cascade_ ));
    InMux I__1092 (
            .O(N__8795),
            .I(N__8792));
    LocalMux I__1091 (
            .O(N__8792),
            .I(\this_vga_signals.g0_i_x2_5_1 ));
    InMux I__1090 (
            .O(N__8789),
            .I(N__8786));
    LocalMux I__1089 (
            .O(N__8786),
            .I(N__8783));
    Odrv4 I__1088 (
            .O(N__8783),
            .I(\this_vga_signals.if_N_13_i_i_1 ));
    CascadeMux I__1087 (
            .O(N__8780),
            .I(\this_vga_signals.g4_0_0_cascade_ ));
    InMux I__1086 (
            .O(N__8777),
            .I(N__8774));
    LocalMux I__1085 (
            .O(N__8774),
            .I(N__8771));
    Odrv4 I__1084 (
            .O(N__8771),
            .I(\this_vga_signals.g0_i_0_N_3L3 ));
    InMux I__1083 (
            .O(N__8768),
            .I(N__8765));
    LocalMux I__1082 (
            .O(N__8765),
            .I(N__8762));
    Odrv4 I__1081 (
            .O(N__8762),
            .I(\this_vga_signals.N_3_1_0_1 ));
    CascadeMux I__1080 (
            .O(N__8759),
            .I(\this_vga_signals.g0_i_x2_1_1_cascade_ ));
    InMux I__1079 (
            .O(N__8756),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    InMux I__1078 (
            .O(N__8753),
            .I(N__8749));
    InMux I__1077 (
            .O(N__8752),
            .I(N__8746));
    LocalMux I__1076 (
            .O(N__8749),
            .I(N__8740));
    LocalMux I__1075 (
            .O(N__8746),
            .I(N__8740));
    InMux I__1074 (
            .O(N__8745),
            .I(N__8737));
    Span4Mux_h I__1073 (
            .O(N__8740),
            .I(N__8734));
    LocalMux I__1072 (
            .O(N__8737),
            .I(N__8731));
    Odrv4 I__1071 (
            .O(N__8734),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    Odrv4 I__1070 (
            .O(N__8731),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    IoInMux I__1069 (
            .O(N__8726),
            .I(N__8723));
    LocalMux I__1068 (
            .O(N__8723),
            .I(N__8720));
    Span4Mux_s2_v I__1067 (
            .O(N__8720),
            .I(N__8717));
    Sp12to4 I__1066 (
            .O(N__8717),
            .I(N__8714));
    Span12Mux_s10_h I__1065 (
            .O(N__8714),
            .I(N__8711));
    Odrv12 I__1064 (
            .O(N__8711),
            .I(N_18));
    InMux I__1063 (
            .O(N__8708),
            .I(N__8705));
    LocalMux I__1062 (
            .O(N__8705),
            .I(\this_vga_signals.hsync_1_i_0_1 ));
    InMux I__1061 (
            .O(N__8702),
            .I(N__8697));
    InMux I__1060 (
            .O(N__8701),
            .I(N__8692));
    InMux I__1059 (
            .O(N__8700),
            .I(N__8692));
    LocalMux I__1058 (
            .O(N__8697),
            .I(N__8689));
    LocalMux I__1057 (
            .O(N__8692),
            .I(N__8686));
    Odrv4 I__1056 (
            .O(N__8689),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    Odrv12 I__1055 (
            .O(N__8686),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    CEMux I__1054 (
            .O(N__8681),
            .I(N__8657));
    CEMux I__1053 (
            .O(N__8680),
            .I(N__8657));
    CEMux I__1052 (
            .O(N__8679),
            .I(N__8657));
    CEMux I__1051 (
            .O(N__8678),
            .I(N__8657));
    CEMux I__1050 (
            .O(N__8677),
            .I(N__8657));
    CEMux I__1049 (
            .O(N__8676),
            .I(N__8657));
    CEMux I__1048 (
            .O(N__8675),
            .I(N__8657));
    CEMux I__1047 (
            .O(N__8674),
            .I(N__8657));
    GlobalMux I__1046 (
            .O(N__8657),
            .I(N__8654));
    gio2CtrlBuf I__1045 (
            .O(N__8654),
            .I(\this_vga_signals.N_469_0_g ));
    InMux I__1044 (
            .O(N__8651),
            .I(N__8648));
    LocalMux I__1043 (
            .O(N__8648),
            .I(N__8636));
    SRMux I__1042 (
            .O(N__8647),
            .I(N__8615));
    SRMux I__1041 (
            .O(N__8646),
            .I(N__8615));
    SRMux I__1040 (
            .O(N__8645),
            .I(N__8615));
    SRMux I__1039 (
            .O(N__8644),
            .I(N__8615));
    SRMux I__1038 (
            .O(N__8643),
            .I(N__8615));
    SRMux I__1037 (
            .O(N__8642),
            .I(N__8615));
    SRMux I__1036 (
            .O(N__8641),
            .I(N__8615));
    SRMux I__1035 (
            .O(N__8640),
            .I(N__8615));
    SRMux I__1034 (
            .O(N__8639),
            .I(N__8615));
    Glb2LocalMux I__1033 (
            .O(N__8636),
            .I(N__8615));
    GlobalMux I__1032 (
            .O(N__8615),
            .I(N__8612));
    gio2CtrlBuf I__1031 (
            .O(N__8612),
            .I(\this_vga_signals.N_608_g ));
    InMux I__1030 (
            .O(N__8609),
            .I(N__8606));
    LocalMux I__1029 (
            .O(N__8606),
            .I(\this_vga_signals.N_381_0 ));
    CascadeMux I__1028 (
            .O(N__8603),
            .I(\this_vga_signals.N_390_cascade_ ));
    CascadeMux I__1027 (
            .O(N__8600),
            .I(\this_vga_signals.rgb_cnst_i_0_2_cascade_ ));
    InMux I__1026 (
            .O(N__8597),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__1025 (
            .O(N__8594),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__1024 (
            .O(N__8591),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__1023 (
            .O(N__8588),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__1022 (
            .O(N__8585),
            .I(N__8582));
    LocalMux I__1021 (
            .O(N__8582),
            .I(N__8578));
    InMux I__1020 (
            .O(N__8581),
            .I(N__8575));
    Span4Mux_h I__1019 (
            .O(N__8578),
            .I(N__8569));
    LocalMux I__1018 (
            .O(N__8575),
            .I(N__8569));
    InMux I__1017 (
            .O(N__8574),
            .I(N__8566));
    Odrv4 I__1016 (
            .O(N__8569),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    LocalMux I__1015 (
            .O(N__8566),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    InMux I__1014 (
            .O(N__8561),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__1013 (
            .O(N__8558),
            .I(N__8555));
    LocalMux I__1012 (
            .O(N__8555),
            .I(N__8552));
    Span12Mux_v I__1011 (
            .O(N__8552),
            .I(N__8547));
    InMux I__1010 (
            .O(N__8551),
            .I(N__8542));
    InMux I__1009 (
            .O(N__8550),
            .I(N__8542));
    Odrv12 I__1008 (
            .O(N__8547),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    LocalMux I__1007 (
            .O(N__8542),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    InMux I__1006 (
            .O(N__8537),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__1005 (
            .O(N__8534),
            .I(N__8531));
    LocalMux I__1004 (
            .O(N__8531),
            .I(N__8526));
    InMux I__1003 (
            .O(N__8530),
            .I(N__8521));
    InMux I__1002 (
            .O(N__8529),
            .I(N__8521));
    Odrv4 I__1001 (
            .O(N__8526),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    LocalMux I__1000 (
            .O(N__8521),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    InMux I__999 (
            .O(N__8516),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__998 (
            .O(N__8513),
            .I(N__8509));
    InMux I__997 (
            .O(N__8512),
            .I(N__8506));
    LocalMux I__996 (
            .O(N__8509),
            .I(N__8502));
    LocalMux I__995 (
            .O(N__8506),
            .I(N__8499));
    InMux I__994 (
            .O(N__8505),
            .I(N__8496));
    Odrv4 I__993 (
            .O(N__8502),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    Odrv4 I__992 (
            .O(N__8499),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__991 (
            .O(N__8496),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    InMux I__990 (
            .O(N__8489),
            .I(bfn_11_24_0_));
    InMux I__989 (
            .O(N__8486),
            .I(N__8483));
    LocalMux I__988 (
            .O(N__8483),
            .I(\this_vga_signals.un11_address_c4_i ));
    CascadeMux I__987 (
            .O(N__8480),
            .I(\this_vga_signals.SUM_2_i_a4_1_0_3_cascade_ ));
    CascadeMux I__986 (
            .O(N__8477),
            .I(\this_vga_signals.un11_address_c5_a0_0_cascade_ ));
    InMux I__985 (
            .O(N__8474),
            .I(N__8470));
    InMux I__984 (
            .O(N__8473),
            .I(N__8467));
    LocalMux I__983 (
            .O(N__8470),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPMZ0Z1 ));
    LocalMux I__982 (
            .O(N__8467),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPMZ0Z1 ));
    InMux I__981 (
            .O(N__8462),
            .I(N__8455));
    InMux I__980 (
            .O(N__8461),
            .I(N__8455));
    InMux I__979 (
            .O(N__8460),
            .I(N__8449));
    LocalMux I__978 (
            .O(N__8455),
            .I(N__8443));
    InMux I__977 (
            .O(N__8454),
            .I(N__8440));
    InMux I__976 (
            .O(N__8453),
            .I(N__8435));
    InMux I__975 (
            .O(N__8452),
            .I(N__8435));
    LocalMux I__974 (
            .O(N__8449),
            .I(N__8432));
    InMux I__973 (
            .O(N__8448),
            .I(N__8425));
    InMux I__972 (
            .O(N__8447),
            .I(N__8425));
    InMux I__971 (
            .O(N__8446),
            .I(N__8425));
    Odrv4 I__970 (
            .O(N__8443),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__969 (
            .O(N__8440),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__968 (
            .O(N__8435),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv4 I__967 (
            .O(N__8432),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__966 (
            .O(N__8425),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    CascadeMux I__965 (
            .O(N__8414),
            .I(N__8406));
    InMux I__964 (
            .O(N__8413),
            .I(N__8401));
    InMux I__963 (
            .O(N__8412),
            .I(N__8401));
    InMux I__962 (
            .O(N__8411),
            .I(N__8396));
    InMux I__961 (
            .O(N__8410),
            .I(N__8396));
    InMux I__960 (
            .O(N__8409),
            .I(N__8391));
    InMux I__959 (
            .O(N__8406),
            .I(N__8391));
    LocalMux I__958 (
            .O(N__8401),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__957 (
            .O(N__8396),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__956 (
            .O(N__8391),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    InMux I__955 (
            .O(N__8384),
            .I(N__8381));
    LocalMux I__954 (
            .O(N__8381),
            .I(N__8375));
    CascadeMux I__953 (
            .O(N__8380),
            .I(N__8372));
    CascadeMux I__952 (
            .O(N__8379),
            .I(N__8368));
    CascadeMux I__951 (
            .O(N__8378),
            .I(N__8364));
    Span4Mux_h I__950 (
            .O(N__8375),
            .I(N__8359));
    InMux I__949 (
            .O(N__8372),
            .I(N__8356));
    InMux I__948 (
            .O(N__8371),
            .I(N__8353));
    InMux I__947 (
            .O(N__8368),
            .I(N__8346));
    InMux I__946 (
            .O(N__8367),
            .I(N__8346));
    InMux I__945 (
            .O(N__8364),
            .I(N__8346));
    InMux I__944 (
            .O(N__8363),
            .I(N__8343));
    InMux I__943 (
            .O(N__8362),
            .I(N__8340));
    Odrv4 I__942 (
            .O(N__8359),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__941 (
            .O(N__8356),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__940 (
            .O(N__8353),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__939 (
            .O(N__8346),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__938 (
            .O(N__8343),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__937 (
            .O(N__8340),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    InMux I__936 (
            .O(N__8327),
            .I(N__8315));
    InMux I__935 (
            .O(N__8326),
            .I(N__8315));
    InMux I__934 (
            .O(N__8325),
            .I(N__8312));
    InMux I__933 (
            .O(N__8324),
            .I(N__8305));
    InMux I__932 (
            .O(N__8323),
            .I(N__8305));
    InMux I__931 (
            .O(N__8322),
            .I(N__8305));
    InMux I__930 (
            .O(N__8321),
            .I(N__8300));
    InMux I__929 (
            .O(N__8320),
            .I(N__8300));
    LocalMux I__928 (
            .O(N__8315),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__927 (
            .O(N__8312),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__926 (
            .O(N__8305),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__925 (
            .O(N__8300),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    CascadeMux I__924 (
            .O(N__8291),
            .I(N__8285));
    CascadeMux I__923 (
            .O(N__8290),
            .I(N__8277));
    InMux I__922 (
            .O(N__8289),
            .I(N__8274));
    InMux I__921 (
            .O(N__8288),
            .I(N__8271));
    InMux I__920 (
            .O(N__8285),
            .I(N__8268));
    InMux I__919 (
            .O(N__8284),
            .I(N__8263));
    InMux I__918 (
            .O(N__8283),
            .I(N__8263));
    InMux I__917 (
            .O(N__8282),
            .I(N__8258));
    InMux I__916 (
            .O(N__8281),
            .I(N__8258));
    InMux I__915 (
            .O(N__8280),
            .I(N__8253));
    InMux I__914 (
            .O(N__8277),
            .I(N__8253));
    LocalMux I__913 (
            .O(N__8274),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__912 (
            .O(N__8271),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__911 (
            .O(N__8268),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__910 (
            .O(N__8263),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__909 (
            .O(N__8258),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__908 (
            .O(N__8253),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    InMux I__907 (
            .O(N__8240),
            .I(N__8230));
    InMux I__906 (
            .O(N__8239),
            .I(N__8230));
    InMux I__905 (
            .O(N__8238),
            .I(N__8230));
    InMux I__904 (
            .O(N__8237),
            .I(N__8225));
    LocalMux I__903 (
            .O(N__8230),
            .I(N__8215));
    InMux I__902 (
            .O(N__8229),
            .I(N__8210));
    InMux I__901 (
            .O(N__8228),
            .I(N__8210));
    LocalMux I__900 (
            .O(N__8225),
            .I(N__8207));
    InMux I__899 (
            .O(N__8224),
            .I(N__8198));
    InMux I__898 (
            .O(N__8223),
            .I(N__8198));
    InMux I__897 (
            .O(N__8222),
            .I(N__8198));
    InMux I__896 (
            .O(N__8221),
            .I(N__8198));
    InMux I__895 (
            .O(N__8220),
            .I(N__8193));
    InMux I__894 (
            .O(N__8219),
            .I(N__8193));
    InMux I__893 (
            .O(N__8218),
            .I(N__8190));
    Span4Mux_v I__892 (
            .O(N__8215),
            .I(N__8185));
    LocalMux I__891 (
            .O(N__8210),
            .I(N__8185));
    Odrv4 I__890 (
            .O(N__8207),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__889 (
            .O(N__8198),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__888 (
            .O(N__8193),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__887 (
            .O(N__8190),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__886 (
            .O(N__8185),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    CascadeMux I__885 (
            .O(N__8174),
            .I(\this_vga_signals.SUM_2_i_a4_0_a0_2_3_cascade_ ));
    InMux I__884 (
            .O(N__8171),
            .I(N__8168));
    LocalMux I__883 (
            .O(N__8168),
            .I(\this_vga_signals.SUM_2_i_a4_a0_2_3 ));
    InMux I__882 (
            .O(N__8165),
            .I(N__8162));
    LocalMux I__881 (
            .O(N__8162),
            .I(\this_vga_signals.SUM_2_i_1_0_3 ));
    InMux I__880 (
            .O(N__8159),
            .I(N__8156));
    LocalMux I__879 (
            .O(N__8156),
            .I(\this_vga_signals.SUM_2_i_0_1_3 ));
    InMux I__878 (
            .O(N__8153),
            .I(N__8150));
    LocalMux I__877 (
            .O(N__8150),
            .I(\this_vga_signals.SUM_2_i_0_3 ));
    CascadeMux I__876 (
            .O(N__8147),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ));
    InMux I__875 (
            .O(N__8144),
            .I(N__8141));
    LocalMux I__874 (
            .O(N__8141),
            .I(N__8138));
    Span4Mux_h I__873 (
            .O(N__8138),
            .I(N__8135));
    Odrv4 I__872 (
            .O(N__8135),
            .I(\this_vga_signals.g0_1 ));
    CascadeMux I__871 (
            .O(N__8132),
            .I(\this_vga_signals.un11_address_c4_i_cascade_ ));
    CascadeMux I__870 (
            .O(N__8129),
            .I(\this_vga_signals.mult1_un54_sum_axb1_5_4_1_cascade_ ));
    InMux I__869 (
            .O(N__8126),
            .I(N__8120));
    InMux I__868 (
            .O(N__8125),
            .I(N__8120));
    LocalMux I__867 (
            .O(N__8120),
            .I(N__8116));
    InMux I__866 (
            .O(N__8119),
            .I(N__8113));
    Odrv4 I__865 (
            .O(N__8116),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABCZ0Z21 ));
    LocalMux I__864 (
            .O(N__8113),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABCZ0Z21 ));
    CascadeMux I__863 (
            .O(N__8108),
            .I(\this_vga_signals.mult1_un54_sum_axb1_5_4_cascade_ ));
    InMux I__862 (
            .O(N__8105),
            .I(N__8095));
    InMux I__861 (
            .O(N__8104),
            .I(N__8095));
    InMux I__860 (
            .O(N__8103),
            .I(N__8095));
    InMux I__859 (
            .O(N__8102),
            .I(N__8092));
    LocalMux I__858 (
            .O(N__8095),
            .I(N__8087));
    LocalMux I__857 (
            .O(N__8092),
            .I(N__8084));
    InMux I__856 (
            .O(N__8091),
            .I(N__8081));
    InMux I__855 (
            .O(N__8090),
            .I(N__8078));
    Span4Mux_h I__854 (
            .O(N__8087),
            .I(N__8075));
    Odrv4 I__853 (
            .O(N__8084),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0 ));
    LocalMux I__852 (
            .O(N__8081),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0 ));
    LocalMux I__851 (
            .O(N__8078),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0 ));
    Odrv4 I__850 (
            .O(N__8075),
            .I(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0 ));
    InMux I__849 (
            .O(N__8066),
            .I(N__8058));
    InMux I__848 (
            .O(N__8065),
            .I(N__8058));
    InMux I__847 (
            .O(N__8064),
            .I(N__8053));
    InMux I__846 (
            .O(N__8063),
            .I(N__8053));
    LocalMux I__845 (
            .O(N__8058),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__844 (
            .O(N__8053),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    CascadeMux I__843 (
            .O(N__8048),
            .I(N__8043));
    CascadeMux I__842 (
            .O(N__8047),
            .I(N__8040));
    CascadeMux I__841 (
            .O(N__8046),
            .I(N__8037));
    InMux I__840 (
            .O(N__8043),
            .I(N__8034));
    InMux I__839 (
            .O(N__8040),
            .I(N__8029));
    InMux I__838 (
            .O(N__8037),
            .I(N__8029));
    LocalMux I__837 (
            .O(N__8034),
            .I(N__8026));
    LocalMux I__836 (
            .O(N__8029),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    Odrv4 I__835 (
            .O(N__8026),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    InMux I__834 (
            .O(N__8021),
            .I(N__8016));
    InMux I__833 (
            .O(N__8020),
            .I(N__8011));
    InMux I__832 (
            .O(N__8019),
            .I(N__8011));
    LocalMux I__831 (
            .O(N__8016),
            .I(N__8008));
    LocalMux I__830 (
            .O(N__8011),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    Odrv4 I__829 (
            .O(N__8008),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    InMux I__828 (
            .O(N__8003),
            .I(N__7998));
    InMux I__827 (
            .O(N__8002),
            .I(N__7995));
    InMux I__826 (
            .O(N__8001),
            .I(N__7992));
    LocalMux I__825 (
            .O(N__7998),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3 ));
    LocalMux I__824 (
            .O(N__7995),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3 ));
    LocalMux I__823 (
            .O(N__7992),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3 ));
    CascadeMux I__822 (
            .O(N__7985),
            .I(N__7981));
    InMux I__821 (
            .O(N__7984),
            .I(N__7976));
    InMux I__820 (
            .O(N__7981),
            .I(N__7976));
    LocalMux I__819 (
            .O(N__7976),
            .I(N__7973));
    Span4Mux_h I__818 (
            .O(N__7973),
            .I(N__7970));
    Odrv4 I__817 (
            .O(N__7970),
            .I(\this_vga_signals.if_N_3_0_i ));
    CascadeMux I__816 (
            .O(N__7967),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_c_cascade_ ));
    InMux I__815 (
            .O(N__7964),
            .I(N__7958));
    InMux I__814 (
            .O(N__7963),
            .I(N__7953));
    InMux I__813 (
            .O(N__7962),
            .I(N__7953));
    InMux I__812 (
            .O(N__7961),
            .I(N__7950));
    LocalMux I__811 (
            .O(N__7958),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1 ));
    LocalMux I__810 (
            .O(N__7953),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1 ));
    LocalMux I__809 (
            .O(N__7950),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1 ));
    InMux I__808 (
            .O(N__7943),
            .I(N__7937));
    InMux I__807 (
            .O(N__7942),
            .I(N__7937));
    LocalMux I__806 (
            .O(N__7937),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_c ));
    InMux I__805 (
            .O(N__7934),
            .I(N__7931));
    LocalMux I__804 (
            .O(N__7931),
            .I(N__7928));
    Span4Mux_v I__803 (
            .O(N__7928),
            .I(N__7925));
    Odrv4 I__802 (
            .O(N__7925),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1_0 ));
    CascadeMux I__801 (
            .O(N__7922),
            .I(N__7919));
    InMux I__800 (
            .O(N__7919),
            .I(N__7916));
    LocalMux I__799 (
            .O(N__7916),
            .I(N__7913));
    Span4Mux_h I__798 (
            .O(N__7913),
            .I(N__7910));
    Odrv4 I__797 (
            .O(N__7910),
            .I(\this_vga_signals.if_N_3_0_i_0 ));
    InMux I__796 (
            .O(N__7907),
            .I(N__7903));
    InMux I__795 (
            .O(N__7906),
            .I(N__7900));
    LocalMux I__794 (
            .O(N__7903),
            .I(N__7895));
    LocalMux I__793 (
            .O(N__7900),
            .I(N__7891));
    InMux I__792 (
            .O(N__7899),
            .I(N__7888));
    InMux I__791 (
            .O(N__7898),
            .I(N__7884));
    Span4Mux_v I__790 (
            .O(N__7895),
            .I(N__7879));
    InMux I__789 (
            .O(N__7894),
            .I(N__7876));
    Span4Mux_h I__788 (
            .O(N__7891),
            .I(N__7873));
    LocalMux I__787 (
            .O(N__7888),
            .I(N__7870));
    InMux I__786 (
            .O(N__7887),
            .I(N__7867));
    LocalMux I__785 (
            .O(N__7884),
            .I(N__7864));
    InMux I__784 (
            .O(N__7883),
            .I(N__7859));
    InMux I__783 (
            .O(N__7882),
            .I(N__7859));
    Odrv4 I__782 (
            .O(N__7879),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    LocalMux I__781 (
            .O(N__7876),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    Odrv4 I__780 (
            .O(N__7873),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    Odrv4 I__779 (
            .O(N__7870),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    LocalMux I__778 (
            .O(N__7867),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    Odrv4 I__777 (
            .O(N__7864),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    LocalMux I__776 (
            .O(N__7859),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    InMux I__775 (
            .O(N__7844),
            .I(N__7838));
    InMux I__774 (
            .O(N__7843),
            .I(N__7835));
    InMux I__773 (
            .O(N__7842),
            .I(N__7827));
    InMux I__772 (
            .O(N__7841),
            .I(N__7824));
    LocalMux I__771 (
            .O(N__7838),
            .I(N__7821));
    LocalMux I__770 (
            .O(N__7835),
            .I(N__7818));
    InMux I__769 (
            .O(N__7834),
            .I(N__7815));
    InMux I__768 (
            .O(N__7833),
            .I(N__7810));
    InMux I__767 (
            .O(N__7832),
            .I(N__7810));
    InMux I__766 (
            .O(N__7831),
            .I(N__7805));
    InMux I__765 (
            .O(N__7830),
            .I(N__7805));
    LocalMux I__764 (
            .O(N__7827),
            .I(N__7802));
    LocalMux I__763 (
            .O(N__7824),
            .I(N__7799));
    Span4Mux_h I__762 (
            .O(N__7821),
            .I(N__7791));
    Span4Mux_v I__761 (
            .O(N__7818),
            .I(N__7791));
    LocalMux I__760 (
            .O(N__7815),
            .I(N__7791));
    LocalMux I__759 (
            .O(N__7810),
            .I(N__7788));
    LocalMux I__758 (
            .O(N__7805),
            .I(N__7781));
    Span4Mux_v I__757 (
            .O(N__7802),
            .I(N__7781));
    Span4Mux_h I__756 (
            .O(N__7799),
            .I(N__7781));
    InMux I__755 (
            .O(N__7798),
            .I(N__7778));
    Odrv4 I__754 (
            .O(N__7791),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_2 ));
    Odrv12 I__753 (
            .O(N__7788),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_2 ));
    Odrv4 I__752 (
            .O(N__7781),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_2 ));
    LocalMux I__751 (
            .O(N__7778),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_2 ));
    InMux I__750 (
            .O(N__7769),
            .I(N__7766));
    LocalMux I__749 (
            .O(N__7766),
            .I(N__7762));
    InMux I__748 (
            .O(N__7765),
            .I(N__7759));
    Odrv4 I__747 (
            .O(N__7762),
            .I(\this_vga_signals.mult1_un54_sum_axb2_0 ));
    LocalMux I__746 (
            .O(N__7759),
            .I(\this_vga_signals.mult1_un54_sum_axb2_0 ));
    CascadeMux I__745 (
            .O(N__7754),
            .I(\this_vga_signals.mult1_un40_sum_axb1_cascade_ ));
    InMux I__744 (
            .O(N__7751),
            .I(N__7747));
    InMux I__743 (
            .O(N__7750),
            .I(N__7744));
    LocalMux I__742 (
            .O(N__7747),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_0 ));
    LocalMux I__741 (
            .O(N__7744),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_0 ));
    InMux I__740 (
            .O(N__7739),
            .I(N__7736));
    LocalMux I__739 (
            .O(N__7736),
            .I(N__7733));
    Odrv4 I__738 (
            .O(N__7733),
            .I(\this_vga_signals.g0_5_1 ));
    InMux I__737 (
            .O(N__7730),
            .I(N__7724));
    InMux I__736 (
            .O(N__7729),
            .I(N__7724));
    LocalMux I__735 (
            .O(N__7724),
            .I(N__7720));
    InMux I__734 (
            .O(N__7723),
            .I(N__7717));
    Odrv4 I__733 (
            .O(N__7720),
            .I(\this_vga_signals.mult1_un47_sum_c2_0 ));
    LocalMux I__732 (
            .O(N__7717),
            .I(\this_vga_signals.mult1_un47_sum_c2_0 ));
    InMux I__731 (
            .O(N__7712),
            .I(N__7709));
    LocalMux I__730 (
            .O(N__7709),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_x1 ));
    CascadeMux I__729 (
            .O(N__7706),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_x0_cascade_ ));
    InMux I__728 (
            .O(N__7703),
            .I(N__7700));
    LocalMux I__727 (
            .O(N__7700),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    CascadeMux I__726 (
            .O(N__7697),
            .I(\this_vga_signals.mult1_un54_sum_i_1_cascade_ ));
    CascadeMux I__725 (
            .O(N__7694),
            .I(\this_vga_signals.un11_address_2_5_cascade_ ));
    CascadeMux I__724 (
            .O(N__7691),
            .I(\this_vga_signals.mult1_un54_sum_i_x0_3_cascade_ ));
    CascadeMux I__723 (
            .O(N__7688),
            .I(N__7685));
    InMux I__722 (
            .O(N__7685),
            .I(N__7681));
    InMux I__721 (
            .O(N__7684),
            .I(N__7678));
    LocalMux I__720 (
            .O(N__7681),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    LocalMux I__719 (
            .O(N__7678),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    InMux I__718 (
            .O(N__7673),
            .I(N__7669));
    InMux I__717 (
            .O(N__7672),
            .I(N__7666));
    LocalMux I__716 (
            .O(N__7669),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    LocalMux I__715 (
            .O(N__7666),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    InMux I__714 (
            .O(N__7661),
            .I(N__7655));
    InMux I__713 (
            .O(N__7660),
            .I(N__7655));
    LocalMux I__712 (
            .O(N__7655),
            .I(N__7651));
    InMux I__711 (
            .O(N__7654),
            .I(N__7648));
    Span4Mux_h I__710 (
            .O(N__7651),
            .I(N__7645));
    LocalMux I__709 (
            .O(N__7648),
            .I(N__7642));
    Odrv4 I__708 (
            .O(N__7645),
            .I(\this_vga_signals.d_N_8_0 ));
    Odrv12 I__707 (
            .O(N__7642),
            .I(\this_vga_signals.d_N_8_0 ));
    CascadeMux I__706 (
            .O(N__7637),
            .I(\this_vga_signals.un11_address_1_5_cascade_ ));
    InMux I__705 (
            .O(N__7634),
            .I(N__7631));
    LocalMux I__704 (
            .O(N__7631),
            .I(\this_vga_signals.g0_11_1 ));
    CascadeMux I__703 (
            .O(N__7628),
            .I(N__7625));
    InMux I__702 (
            .O(N__7625),
            .I(N__7622));
    LocalMux I__701 (
            .O(N__7622),
            .I(\this_vga_signals.g0_6_0 ));
    CascadeMux I__700 (
            .O(N__7619),
            .I(\this_vga_signals.g2_1_0_cascade_ ));
    CascadeMux I__699 (
            .O(N__7616),
            .I(\this_vga_signals.g3_cascade_ ));
    InMux I__698 (
            .O(N__7613),
            .I(N__7610));
    LocalMux I__697 (
            .O(N__7610),
            .I(\this_vga_signals.g2_4_0 ));
    CascadeMux I__696 (
            .O(N__7607),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_2_N_2L1_cascade_ ));
    InMux I__695 (
            .O(N__7604),
            .I(N__7598));
    InMux I__694 (
            .O(N__7603),
            .I(N__7598));
    LocalMux I__693 (
            .O(N__7598),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    InMux I__692 (
            .O(N__7595),
            .I(N__7592));
    LocalMux I__691 (
            .O(N__7592),
            .I(N__7589));
    Span4Mux_h I__690 (
            .O(N__7589),
            .I(N__7586));
    Odrv4 I__689 (
            .O(N__7586),
            .I(\this_vga_signals.un11_address_0_5 ));
    InMux I__688 (
            .O(N__7583),
            .I(N__7580));
    LocalMux I__687 (
            .O(N__7580),
            .I(N__7577));
    Odrv4 I__686 (
            .O(N__7577),
            .I(\this_vga_signals.vsync_1_0_a3_4 ));
    CascadeMux I__685 (
            .O(N__7574),
            .I(N__7571));
    InMux I__684 (
            .O(N__7571),
            .I(N__7568));
    LocalMux I__683 (
            .O(N__7568),
            .I(N__7565));
    Odrv4 I__682 (
            .O(N__7565),
            .I(\this_vga_signals.if_N_15_mux ));
    CascadeMux I__681 (
            .O(N__7562),
            .I(\this_vga_signals.if_m13_ns_1_cascade_ ));
    InMux I__680 (
            .O(N__7559),
            .I(N__7556));
    LocalMux I__679 (
            .O(N__7556),
            .I(N__7552));
    CascadeMux I__678 (
            .O(N__7555),
            .I(N__7549));
    Span4Mux_h I__677 (
            .O(N__7552),
            .I(N__7545));
    InMux I__676 (
            .O(N__7549),
            .I(N__7540));
    InMux I__675 (
            .O(N__7548),
            .I(N__7540));
    Odrv4 I__674 (
            .O(N__7545),
            .I(\this_vga_signals.if_m13_ns ));
    LocalMux I__673 (
            .O(N__7540),
            .I(\this_vga_signals.if_m13_ns ));
    InMux I__672 (
            .O(N__7535),
            .I(N__7532));
    LocalMux I__671 (
            .O(N__7532),
            .I(\this_vga_signals.if_N_7 ));
    InMux I__670 (
            .O(N__7529),
            .I(N__7526));
    LocalMux I__669 (
            .O(N__7526),
            .I(\this_vga_signals.d_N_9_0 ));
    CascadeMux I__668 (
            .O(N__7523),
            .I(\this_vga_signals.rgb_1_4_cascade_ ));
    InMux I__667 (
            .O(N__7520),
            .I(N__7516));
    CascadeMux I__666 (
            .O(N__7519),
            .I(N__7513));
    LocalMux I__665 (
            .O(N__7516),
            .I(N__7509));
    InMux I__664 (
            .O(N__7513),
            .I(N__7504));
    InMux I__663 (
            .O(N__7512),
            .I(N__7504));
    Span4Mux_v I__662 (
            .O(N__7509),
            .I(N__7499));
    LocalMux I__661 (
            .O(N__7504),
            .I(N__7499));
    Odrv4 I__660 (
            .O(N__7499),
            .I(\this_vga_signals.M_vcounter_q_9_rep1_esr_RNIETZ0Z844 ));
    InMux I__659 (
            .O(N__7496),
            .I(N__7493));
    LocalMux I__658 (
            .O(N__7493),
            .I(\this_vga_signals.d_N_5_0 ));
    CascadeMux I__657 (
            .O(N__7490),
            .I(N__7487));
    InMux I__656 (
            .O(N__7487),
            .I(N__7484));
    LocalMux I__655 (
            .O(N__7484),
            .I(N__7481));
    Odrv4 I__654 (
            .O(N__7481),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1 ));
    CascadeMux I__653 (
            .O(N__7478),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ));
    CascadeMux I__652 (
            .O(N__7475),
            .I(N__7472));
    InMux I__651 (
            .O(N__7472),
            .I(N__7469));
    LocalMux I__650 (
            .O(N__7469),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_i_x1 ));
    InMux I__649 (
            .O(N__7466),
            .I(N__7463));
    LocalMux I__648 (
            .O(N__7463),
            .I(N__7460));
    Odrv4 I__647 (
            .O(N__7460),
            .I(\this_vga_signals.g1 ));
    CascadeMux I__646 (
            .O(N__7457),
            .I(\this_vga_signals.g3_0_2_cascade_ ));
    InMux I__645 (
            .O(N__7454),
            .I(N__7451));
    LocalMux I__644 (
            .O(N__7451),
            .I(\this_vga_signals.if_N_3_0_i_1 ));
    CascadeMux I__643 (
            .O(N__7448),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_c_0_cascade_ ));
    InMux I__642 (
            .O(N__7445),
            .I(N__7442));
    LocalMux I__641 (
            .O(N__7442),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_1 ));
    CascadeMux I__640 (
            .O(N__7439),
            .I(\this_vga_signals.mult1_un47_sum_ac0_1_cascade_ ));
    CascadeMux I__639 (
            .O(N__7436),
            .I(\this_vga_signals.rgb_1_2_cascade_ ));
    InMux I__638 (
            .O(N__7433),
            .I(N__7430));
    LocalMux I__637 (
            .O(N__7430),
            .I(N__7427));
    Odrv4 I__636 (
            .O(N__7427),
            .I(\this_vga_signals.if_i3_mux_0_0 ));
    InMux I__635 (
            .O(N__7424),
            .I(N__7420));
    CascadeMux I__634 (
            .O(N__7423),
            .I(N__7417));
    LocalMux I__633 (
            .O(N__7420),
            .I(N__7414));
    InMux I__632 (
            .O(N__7417),
            .I(N__7411));
    Odrv4 I__631 (
            .O(N__7414),
            .I(\this_vga_signals.if_i3_mux_2 ));
    LocalMux I__630 (
            .O(N__7411),
            .I(\this_vga_signals.if_i3_mux_2 ));
    CascadeMux I__629 (
            .O(N__7406),
            .I(\this_vga_signals.g2_1_cascade_ ));
    InMux I__628 (
            .O(N__7403),
            .I(N__7400));
    LocalMux I__627 (
            .O(N__7400),
            .I(\this_vga_signals.g2_1 ));
    InMux I__626 (
            .O(N__7397),
            .I(N__7394));
    LocalMux I__625 (
            .O(N__7394),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1_1_0 ));
    CascadeMux I__624 (
            .O(N__7391),
            .I(N__7388));
    InMux I__623 (
            .O(N__7388),
            .I(N__7385));
    LocalMux I__622 (
            .O(N__7385),
            .I(\this_vga_signals.g0_5_0_1 ));
    InMux I__621 (
            .O(N__7382),
            .I(N__7379));
    LocalMux I__620 (
            .O(N__7379),
            .I(\this_vga_signals.g3_0_2_0 ));
    CascadeMux I__619 (
            .O(N__7376),
            .I(\this_vga_signals.g2_cascade_ ));
    InMux I__618 (
            .O(N__7373),
            .I(N__7370));
    LocalMux I__617 (
            .O(N__7370),
            .I(\this_vga_signals.g0_3_0_0 ));
    CascadeMux I__616 (
            .O(N__7367),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_2_0_cascade_ ));
    CascadeMux I__615 (
            .O(N__7364),
            .I(N__7361));
    InMux I__614 (
            .O(N__7361),
            .I(N__7358));
    LocalMux I__613 (
            .O(N__7358),
            .I(\this_vga_signals.if_m1_3 ));
    InMux I__612 (
            .O(N__7355),
            .I(N__7352));
    LocalMux I__611 (
            .O(N__7352),
            .I(\this_vga_signals.if_N_4_2 ));
    CascadeMux I__610 (
            .O(N__7349),
            .I(\this_vga_signals.if_i4_mux_0_1_cascade_ ));
    CascadeMux I__609 (
            .O(N__7346),
            .I(\this_vga_signals.vsync_1_0_a3_5_cascade_ ));
    IoInMux I__608 (
            .O(N__7343),
            .I(N__7340));
    LocalMux I__607 (
            .O(N__7340),
            .I(N__7337));
    Span12Mux_s10_v I__606 (
            .O(N__7337),
            .I(N__7334));
    Odrv12 I__605 (
            .O(N__7334),
            .I(this_vga_signals_vsync_1_i));
    CascadeMux I__604 (
            .O(N__7331),
            .I(\this_vga_signals.if_m13_0_ns_1_cascade_ ));
    CascadeMux I__603 (
            .O(N__7328),
            .I(\this_vga_signals.if_i3_mux_0_0_cascade_ ));
    CascadeMux I__602 (
            .O(N__7325),
            .I(N__7322));
    InMux I__601 (
            .O(N__7322),
            .I(N__7319));
    LocalMux I__600 (
            .O(N__7319),
            .I(\this_vga_signals.if_m13_0_ns_1 ));
    InMux I__599 (
            .O(N__7316),
            .I(N__7313));
    LocalMux I__598 (
            .O(N__7313),
            .I(N__7310));
    Odrv12 I__597 (
            .O(N__7310),
            .I(\this_vga_signals.if_i3_mux_0_0_0 ));
    CascadeMux I__596 (
            .O(N__7307),
            .I(\this_vga_signals.if_m8_0_ns_1_cascade_ ));
    CascadeMux I__595 (
            .O(N__7304),
            .I(\this_vga_signals.g1_1_cascade_ ));
    CascadeMux I__594 (
            .O(N__7301),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ));
    CascadeMux I__593 (
            .O(N__7298),
            .I(\this_vga_signals.g1_cascade_ ));
    CascadeMux I__592 (
            .O(N__7295),
            .I(\this_vga_signals.if_m1_3_cascade_ ));
    InMux I__591 (
            .O(N__7292),
            .I(N__7280));
    InMux I__590 (
            .O(N__7291),
            .I(N__7280));
    InMux I__589 (
            .O(N__7290),
            .I(N__7280));
    InMux I__588 (
            .O(N__7289),
            .I(N__7280));
    LocalMux I__587 (
            .O(N__7280),
            .I(N__7277));
    Span4Mux_v I__586 (
            .O(N__7277),
            .I(N__7274));
    Sp12to4 I__585 (
            .O(N__7274),
            .I(N__7271));
    Span12Mux_h I__584 (
            .O(N__7271),
            .I(N__7268));
    Span12Mux_v I__583 (
            .O(N__7268),
            .I(N__7265));
    Odrv12 I__582 (
            .O(N__7265),
            .I(rst_n_c));
    InMux I__581 (
            .O(N__7262),
            .I(N__7259));
    LocalMux I__580 (
            .O(N__7259),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    CascadeMux I__579 (
            .O(N__7256),
            .I(\this_vga_signals.if_i3_mux_2_0_cascade_ ));
    CascadeMux I__578 (
            .O(N__7253),
            .I(\this_vga_signals.if_m2_8_0_cascade_ ));
    InMux I__577 (
            .O(N__7250),
            .I(N__7247));
    LocalMux I__576 (
            .O(N__7247),
            .I(\this_vga_signals.if_m8_0_ns_1 ));
    InMux I__575 (
            .O(N__7244),
            .I(N__7241));
    LocalMux I__574 (
            .O(N__7241),
            .I(\this_vga_signals.rgb_cnst_i_1Z0Z_5 ));
    IoInMux I__573 (
            .O(N__7238),
            .I(N__7235));
    LocalMux I__572 (
            .O(N__7235),
            .I(N__7232));
    Span4Mux_s1_h I__571 (
            .O(N__7232),
            .I(N__7229));
    Span4Mux_h I__570 (
            .O(N__7229),
            .I(N__7226));
    Span4Mux_v I__569 (
            .O(N__7226),
            .I(N__7223));
    Odrv4 I__568 (
            .O(N__7223),
            .I(rgb_c_5));
    InMux I__567 (
            .O(N__7220),
            .I(N__7217));
    LocalMux I__566 (
            .O(N__7217),
            .I(N__7214));
    Odrv4 I__565 (
            .O(N__7214),
            .I(\this_vga_signals.M_vcounter_q_esr_RNIAV48E1Z0Z_9 ));
    IoInMux I__564 (
            .O(N__7211),
            .I(N__7208));
    LocalMux I__563 (
            .O(N__7208),
            .I(N__7205));
    IoSpan4Mux I__562 (
            .O(N__7205),
            .I(N__7202));
    IoSpan4Mux I__561 (
            .O(N__7202),
            .I(N__7199));
    Span4Mux_s2_h I__560 (
            .O(N__7199),
            .I(N__7196));
    Odrv4 I__559 (
            .O(N__7196),
            .I(rgb_c_3));
    InMux I__558 (
            .O(N__7193),
            .I(N__7189));
    InMux I__557 (
            .O(N__7192),
            .I(N__7186));
    LocalMux I__556 (
            .O(N__7189),
            .I(\this_vga_signals.N_379_0 ));
    LocalMux I__555 (
            .O(N__7186),
            .I(\this_vga_signals.N_379_0 ));
    CascadeMux I__554 (
            .O(N__7181),
            .I(\this_vga_signals.M_vcounter_q_esr_RNIA99QRZ0Z_9_cascade_ ));
    IoInMux I__553 (
            .O(N__7178),
            .I(N__7175));
    LocalMux I__552 (
            .O(N__7175),
            .I(N__7172));
    Span4Mux_s3_h I__551 (
            .O(N__7172),
            .I(N__7169));
    Odrv4 I__550 (
            .O(N__7169),
            .I(rgb_c_1));
    InMux I__549 (
            .O(N__7166),
            .I(N__7163));
    LocalMux I__548 (
            .O(N__7163),
            .I(\this_vga_signals.rgb_cnst_i_0_5 ));
    IoInMux I__547 (
            .O(N__7160),
            .I(N__7157));
    LocalMux I__546 (
            .O(N__7157),
            .I(N__7153));
    InMux I__545 (
            .O(N__7156),
            .I(N__7150));
    IoSpan4Mux I__544 (
            .O(N__7153),
            .I(N__7147));
    LocalMux I__543 (
            .O(N__7150),
            .I(N__7144));
    Sp12to4 I__542 (
            .O(N__7147),
            .I(N__7141));
    Span4Mux_v I__541 (
            .O(N__7144),
            .I(N__7138));
    Span12Mux_s6_h I__540 (
            .O(N__7141),
            .I(N__7135));
    Span4Mux_v I__539 (
            .O(N__7138),
            .I(N__7132));
    Odrv12 I__538 (
            .O(N__7135),
            .I(N_11_0));
    Odrv4 I__537 (
            .O(N__7132),
            .I(N_11_0));
    InMux I__536 (
            .O(N__7127),
            .I(N__7124));
    LocalMux I__535 (
            .O(N__7124),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__534 (
            .O(N__7121),
            .I(N__7118));
    LocalMux I__533 (
            .O(N__7118),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__532 (
            .O(N__7115),
            .I(N__7112));
    LocalMux I__531 (
            .O(N__7112),
            .I(N__7109));
    Odrv4 I__530 (
            .O(N__7109),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    InMux I__529 (
            .O(N__7106),
            .I(N__7103));
    LocalMux I__528 (
            .O(N__7103),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    IoInMux I__527 (
            .O(N__7100),
            .I(N__7097));
    LocalMux I__526 (
            .O(N__7097),
            .I(N__7094));
    Odrv12 I__525 (
            .O(N__7094),
            .I(N_33));
    IoInMux I__524 (
            .O(N__7091),
            .I(N__7088));
    LocalMux I__523 (
            .O(N__7088),
            .I(N__7085));
    Odrv12 I__522 (
            .O(N__7085),
            .I(N_11));
    IoInMux I__521 (
            .O(N__7082),
            .I(N__7079));
    LocalMux I__520 (
            .O(N__7079),
            .I(N__7076));
    Span4Mux_s1_h I__519 (
            .O(N__7076),
            .I(N__7073));
    Span4Mux_v I__518 (
            .O(N__7073),
            .I(N__7070));
    Span4Mux_v I__517 (
            .O(N__7070),
            .I(N__7067));
    Span4Mux_h I__516 (
            .O(N__7067),
            .I(N__7064));
    Odrv4 I__515 (
            .O(N__7064),
            .I(rgb_c_0));
    InMux I__514 (
            .O(N__7061),
            .I(N__7058));
    LocalMux I__513 (
            .O(N__7058),
            .I(\this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1Z0Z_9 ));
    CascadeMux I__512 (
            .O(N__7055),
            .I(\this_vga_signals.rgb_cnst_i_1Z0Z_3_cascade_ ));
    InMux I__511 (
            .O(N__7052),
            .I(N__7049));
    LocalMux I__510 (
            .O(N__7049),
            .I(port_clk_c));
    IoInMux I__509 (
            .O(N__7046),
            .I(N__7043));
    LocalMux I__508 (
            .O(N__7043),
            .I(N__7040));
    Span4Mux_s0_h I__507 (
            .O(N__7040),
            .I(N__7037));
    Odrv4 I__506 (
            .O(N__7037),
            .I(\this_vga_signals.N_469_0 ));
    IoInMux I__505 (
            .O(N__7034),
            .I(N__7031));
    LocalMux I__504 (
            .O(N__7031),
            .I(port_rw_c_i));
    InMux I__503 (
            .O(N__7028),
            .I(N__7025));
    LocalMux I__502 (
            .O(N__7025),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    defparam IN_MUX_bfv_12_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_24_0_));
    defparam IN_MUX_bfv_12_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_25_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_12_25_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(un1_M_current_address_q_cry_7),
            .carryinitout(bfn_15_22_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNIVV6F6_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__9515),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_608_g ));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNIIR7M7_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__7046),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_469_0_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_1_19_1 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_1_19_1 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_1_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7052),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18231),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIR7M7_9_LC_1_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIR7M7_9_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIR7M7_9_LC_1_19_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIR7M7_9_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(N__11706),
            .in2(_gnd_net_),
            .in3(N__8651),
            .lcout(\this_vga_signals.N_469_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_rw_obuf_RNO_LC_1_21_0.C_ON=1'b0;
    defparam port_data_rw_obuf_RNO_LC_1_21_0.SEQ_MODE=4'b0000;
    defparam port_data_rw_obuf_RNO_LC_1_21_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 port_data_rw_obuf_RNO_LC_1_21_0 (
            .in0(N__12781),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(port_rw_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_3_19_2 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_3_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7106),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18230),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_3_19_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_3_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7028),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18230),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_3_19_7 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_3_19_7 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_3_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7115),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18230),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_3_28_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_3_28_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_3_28_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_3_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9281),
            .lcout(N_33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEC104_0_9_LC_5_27_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEC104_0_9_LC_5_27_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEC104_0_9_LC_5_27_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIEC104_0_9_LC_5_27_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7156),
            .lcout(N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI18GF6U3_9_LC_6_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI18GF6U3_9_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI18GF6U3_9_LC_6_15_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI18GF6U3_9_LC_6_15_2  (
            .in0(N__14091),
            .in1(N__7061),
            .in2(_gnd_net_),
            .in3(N__12926),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1_9_LC_6_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1_9_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1_9_LC_6_16_0 .LUT_INIT=16'b0001101000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1_9_LC_6_16_0  (
            .in0(N__10413),
            .in1(N__13774),
            .in2(N__12988),
            .in3(N__20309),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.rgb_cnst_i_1_3_LC_6_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.rgb_cnst_i_1_3_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.rgb_cnst_i_1_3_LC_6_18_5 .LUT_INIT=16'b1101111011101111;
    LogicCell40 \this_vga_signals.rgb_cnst_i_1_3_LC_6_18_5  (
            .in0(N__15904),
            .in1(N__10420),
            .in2(N__13787),
            .in3(N__13007),
            .lcout(),
            .ltout(\this_vga_signals.rgb_cnst_i_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIAV48E1_9_LC_6_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIAV48E1_9_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIAV48E1_9_LC_6_18_6 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIAV48E1_9_LC_6_18_6  (
            .in0(N__10436),
            .in1(N__7192),
            .in2(N__7055),
            .in3(N__13775),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNIAV48E1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGGSVD_9_LC_6_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGGSVD_9_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGGSVD_9_LC_6_19_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGGSVD_9_LC_6_19_0  (
            .in0(N__13008),
            .in1(N__13788),
            .in2(_gnd_net_),
            .in3(N__20331),
            .lcout(\this_vga_signals.N_379_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.rgb_cnst_i_1_5_LC_6_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.rgb_cnst_i_1_5_LC_6_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.rgb_cnst_i_1_5_LC_6_19_5 .LUT_INIT=16'b1101101111001111;
    LogicCell40 \this_vga_signals.rgb_cnst_i_1_5_LC_6_19_5  (
            .in0(N__10421),
            .in1(N__15905),
            .in2(N__13793),
            .in3(N__13009),
            .lcout(\this_vga_signals.rgb_cnst_i_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9UBTOU3_9_LC_6_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9UBTOU3_9_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9UBTOU3_9_LC_6_20_2 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI9UBTOU3_9_LC_6_20_2  (
            .in0(N__7244),
            .in1(N__14092),
            .in2(N__14849),
            .in3(N__7166),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIDP942V3_9_LC_6_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIDP942V3_9_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIDP942V3_9_LC_6_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIDP942V3_9_LC_6_20_3  (
            .in0(N__14093),
            .in1(N__7220),
            .in2(_gnd_net_),
            .in3(N__13055),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA99QR_9_LC_7_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA99QR_9_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA99QR_9_LC_7_18_1 .LUT_INIT=16'b1010101000000010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIA99QR_9_LC_7_18_1  (
            .in0(N__7193),
            .in1(N__10411),
            .in2(N__13010),
            .in3(N__15903),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_esr_RNIA99QRZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNID3EMFU3_9_LC_7_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNID3EMFU3_9_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNID3EMFU3_9_LC_7_18_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNID3EMFU3_9_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(N__14084),
            .in2(N__7181),
            .in3(N__11540),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_9_LC_7_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_9_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_9_LC_7_19_0 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_9_LC_7_19_0  (
            .in0(N__10412),
            .in1(N__13006),
            .in2(N__13792),
            .in3(N__20330),
            .lcout(\this_vga_signals.rgb_cnst_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_7_22_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_7_22_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_7_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7289),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18226),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEC104_9_LC_7_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEC104_9_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEC104_9_LC_7_22_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIEC104_9_LC_7_22_2  (
            .in0(N__9167),
            .in1(N__9593),
            .in2(_gnd_net_),
            .in3(N__9260),
            .lcout(N_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_7_22_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_7_22_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_7_22_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_7_22_5  (
            .in0(N__7290),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7127),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18226),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_7_22_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_7_22_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_7_22_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_7_22_6  (
            .in0(_gnd_net_),
            .in1(N__7291),
            .in2(_gnd_net_),
            .in3(N__7121),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18226),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_7_22_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_7_22_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_7_22_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_7_22_7  (
            .in0(N__7292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7262),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18226),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_3_1_LC_9_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_3_1_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_3_1_LC_9_18_1 .LUT_INIT=16'b1000010010100101;
    LogicCell40 \this_vga_signals.un16_address_g0_3_1_LC_9_18_1  (
            .in0(N__9821),
            .in1(N__7559),
            .in2(N__11464),
            .in3(N__7520),
            .lcout(\this_vga_signals.g0_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_26_LC_9_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_26_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_26_LC_9_19_1 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \this_vga_signals.un16_address_g0_26_LC_9_19_1  (
            .in0(N__9365),
            .in1(N__7250),
            .in2(_gnd_net_),
            .in3(N__9794),
            .lcout(),
            .ltout(\this_vga_signals.if_i3_mux_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_24_LC_9_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_24_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_24_LC_9_19_2 .LUT_INIT=16'b0001000100110000;
    LogicCell40 \this_vga_signals.un16_address_g0_24_LC_9_19_2  (
            .in0(N__7316),
            .in1(N__8240),
            .in2(N__7256),
            .in3(N__18342),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_5_2_LC_9_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_5_2_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_5_2_LC_9_19_3 .LUT_INIT=16'b0000111101011010;
    LogicCell40 \this_vga_signals.un16_address_g0_5_2_LC_9_19_3  (
            .in0(N__8239),
            .in1(_gnd_net_),
            .in2(N__9392),
            .in3(N__9795),
            .lcout(\this_vga_signals.g0_5_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m2_8_0_LC_9_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m2_8_0_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m2_8_0_LC_9_19_4 .LUT_INIT=16'b0011001101100110;
    LogicCell40 \this_vga_signals.un16_address_if_m2_8_0_LC_9_19_4  (
            .in0(N__9793),
            .in1(N__9364),
            .in2(_gnd_net_),
            .in3(N__8238),
            .lcout(),
            .ltout(\this_vga_signals.if_m2_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m2_8_LC_9_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m2_8_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m2_8_LC_9_19_5 .LUT_INIT=16'b1100001100001111;
    LogicCell40 \this_vga_signals.un16_address_if_m2_8_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__7887),
            .in2(N__7253),
            .in3(N__7841),
            .lcout(\this_vga_signals.if_N_3_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_9_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_9_19_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_9_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8585),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18212),
            .ce(N__8674),
            .sr(N__8647));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_9_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_9_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8558),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18212),
            .ce(N__8674),
            .sr(N__8647));
    defparam \this_vga_signals.un16_address_if_m8_0_ns_1_LC_9_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m8_0_ns_1_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m8_0_ns_1_LC_9_20_0 .LUT_INIT=16'b0101101100100100;
    LogicCell40 \this_vga_signals.un16_address_if_m8_0_ns_1_LC_9_20_0  (
            .in0(N__9740),
            .in1(N__9357),
            .in2(N__9250),
            .in3(N__9472),
            .lcout(\this_vga_signals.if_m8_0_ns_1 ),
            .ltout(\this_vga_signals.if_m8_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m8_0_ns_LC_9_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m8_0_ns_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m8_0_ns_LC_9_20_1 .LUT_INIT=16'b1010000001011010;
    LogicCell40 \this_vga_signals.un16_address_if_m8_0_ns_LC_9_20_1  (
            .in0(N__9358),
            .in1(_gnd_net_),
            .in2(N__7307),
            .in3(N__9832),
            .lcout(\this_vga_signals.if_i3_mux_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g1_1_LC_9_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g1_1_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g1_1_LC_9_20_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.un16_address_g1_1_LC_9_20_2  (
            .in0(N__9833),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11426),
            .lcout(),
            .ltout(\this_vga_signals.g1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_14_LC_9_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_14_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_14_LC_9_20_3 .LUT_INIT=16'b0110100110100101;
    LogicCell40 \this_vga_signals.un16_address_g0_14_LC_9_20_3  (
            .in0(N__9359),
            .in1(N__7894),
            .in2(N__7304),
            .in3(N__7831),
            .lcout(\this_vga_signals.if_N_3_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_20_5 .LUT_INIT=16'b0000101100011101;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_20_5  (
            .in0(N__8384),
            .in1(N__9223),
            .in2(N__7490),
            .in3(N__9739),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1 ),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g1_LC_9_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g1_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g1_LC_9_20_6 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \this_vga_signals.un16_address_g1_LC_9_20_6  (
            .in0(N__7830),
            .in1(_gnd_net_),
            .in2(N__7301),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.g1 ),
            .ltout(\this_vga_signals.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_22_LC_9_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_22_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_22_LC_9_20_7 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \this_vga_signals.un16_address_g0_22_LC_9_20_7  (
            .in0(N__9360),
            .in1(N__11427),
            .in2(N__7298),
            .in3(N__9834),
            .lcout(\this_vga_signals.if_N_3_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m1_3_LC_9_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m1_3_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m1_3_LC_9_21_1 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.un16_address_if_m1_3_LC_9_21_1  (
            .in0(N__9379),
            .in1(N__8229),
            .in2(_gnd_net_),
            .in3(N__8284),
            .lcout(\this_vga_signals.if_m1_3 ),
            .ltout(\this_vga_signals.if_m1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m3_1_LC_9_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m3_1_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m3_1_LC_9_21_2 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \this_vga_signals.un16_address_if_m3_1_LC_9_21_2  (
            .in0(N__9727),
            .in1(_gnd_net_),
            .in2(N__7295),
            .in3(N__9228),
            .lcout(\this_vga_signals.if_N_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_9_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_9_21_3 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_9_21_3  (
            .in0(N__9378),
            .in1(N__8228),
            .in2(_gnd_net_),
            .in3(N__8283),
            .lcout(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m7_1_LC_9_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m7_1_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m7_1_LC_9_21_4 .LUT_INIT=16'b0000100000000001;
    LogicCell40 \this_vga_signals.un16_address_if_m7_1_LC_9_21_4  (
            .in0(N__9728),
            .in1(N__9473),
            .in2(N__7364),
            .in3(N__9229),
            .lcout(),
            .ltout(\this_vga_signals.if_i4_mux_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m8_1_LC_9_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m8_1_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m8_1_LC_9_21_5 .LUT_INIT=16'b1101100011100100;
    LogicCell40 \this_vga_signals.un16_address_if_m8_1_LC_9_21_5  (
            .in0(N__9474),
            .in1(N__7355),
            .in2(N__7349),
            .in3(N__18297),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_9_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_9_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8753),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18220),
            .ce(N__8675),
            .sr(N__8646));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI2GCG1_7_LC_9_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI2GCG1_7_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI2GCG1_7_LC_9_22_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI2GCG1_7_LC_9_22_1  (
            .in0(N__11395),
            .in1(N__12169),
            .in2(N__9402),
            .in3(N__9711),
            .lcout(),
            .ltout(\this_vga_signals.vsync_1_0_a3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_9_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_9_22_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_9_22_2  (
            .in0(N__7583),
            .in1(N__9471),
            .in2(N__7346),
            .in3(N__12476),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m13_0_ns_1_LC_9_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m13_0_ns_1_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m13_0_ns_1_LC_9_22_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.un16_address_if_m13_0_ns_1_LC_9_22_3  (
            .in0(N__9470),
            .in1(N__9227),
            .in2(_gnd_net_),
            .in3(N__9710),
            .lcout(\this_vga_signals.if_m13_0_ns_1 ),
            .ltout(\this_vga_signals.if_m13_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m13_0_ns_LC_9_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m13_0_ns_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m13_0_ns_LC_9_22_4 .LUT_INIT=16'b1110110101100101;
    LogicCell40 \this_vga_signals.un16_address_if_m13_0_ns_LC_9_22_4  (
            .in0(N__9830),
            .in1(N__9380),
            .in2(N__7331),
            .in3(N__7660),
            .lcout(\this_vga_signals.if_i3_mux_0_0 ),
            .ltout(\this_vga_signals.if_i3_mux_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_15_LC_9_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_15_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_15_LC_9_22_5 .LUT_INIT=16'b0000010101000100;
    LogicCell40 \this_vga_signals.un16_address_g0_15_LC_9_22_5  (
            .in0(N__11394),
            .in1(N__7424),
            .in2(N__7328),
            .in3(N__18322),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_34_LC_9_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_34_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_34_LC_9_22_6 .LUT_INIT=16'b1110110101100101;
    LogicCell40 \this_vga_signals.un16_address_g0_34_LC_9_22_6  (
            .in0(N__9831),
            .in1(N__9381),
            .in2(N__7325),
            .in3(N__7661),
            .lcout(\this_vga_signals.if_i3_mux_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m11_1_LC_9_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m11_1_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m11_1_LC_9_23_0 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \this_vga_signals.un16_address_if_m11_1_LC_9_23_0  (
            .in0(N__7673),
            .in1(N__8371),
            .in2(N__7688),
            .in3(N__8454),
            .lcout(\this_vga_signals.if_N_15_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_9_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_9_24_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_9_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_9_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8745),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18227),
            .ce(N__8680),
            .sr(N__8642));
    defparam \this_vga_signals.un16_address_g2_3_LC_10_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g2_3_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g2_3_LC_10_18_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \this_vga_signals.un16_address_g2_3_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__7899),
            .in2(_gnd_net_),
            .in3(N__7842),
            .lcout(\this_vga_signals.g2_1 ),
            .ltout(\this_vga_signals.g2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g3_0_LC_10_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g3_0_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g3_0_LC_10_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_g3_0_LC_10_18_1  (
            .in0(N__11409),
            .in1(N__9852),
            .in2(N__7406),
            .in3(N__8990),
            .lcout(\this_vga_signals.g3_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g2_LC_10_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g2_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g2_LC_10_18_2 .LUT_INIT=16'b0001001001111011;
    LogicCell40 \this_vga_signals.un16_address_g2_LC_10_18_2  (
            .in0(N__7403),
            .in1(N__7397),
            .in2(N__7391),
            .in3(N__17321),
            .lcout(),
            .ltout(\this_vga_signals.g2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_13_LC_10_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_13_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_13_LC_10_18_3 .LUT_INIT=16'b1001000011110000;
    LogicCell40 \this_vga_signals.un16_address_g0_13_LC_10_18_3  (
            .in0(N__17322),
            .in1(N__7382),
            .in2(N__7376),
            .in3(N__7373),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_12_LC_10_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_12_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_12_LC_10_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_g0_12_LC_10_18_4  (
            .in0(N__17111),
            .in1(N__8144),
            .in2(N__7367),
            .in3(N__11146),
            .lcout(\this_vga_signals.N_3_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_0_N_3L3_LC_10_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_0_N_3L3_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_0_N_3L3_LC_10_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un16_address_g0_i_0_N_3L3_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__12330),
            .in2(N__17160),
            .in3(N__11145),
            .lcout(\this_vga_signals.g0_i_0_N_3L3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_x2_2_LC_10_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_x2_2_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_x2_2_LC_10_18_7 .LUT_INIT=16'b0110100101011010;
    LogicCell40 \this_vga_signals.un16_address_g0_i_x2_2_LC_10_18_7  (
            .in0(N__11512),
            .in1(N__12516),
            .in2(N__11456),
            .in3(N__12552),
            .lcout(\this_vga_signals.g0_i_x2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g4_0_LC_10_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g4_0_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g4_0_LC_10_19_0 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \this_vga_signals.un16_address_g4_0_LC_10_19_0  (
            .in0(N__11417),
            .in1(N__7445),
            .in2(N__12363),
            .in3(N__10901),
            .lcout(\this_vga_signals.g4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_5_1_0_LC_10_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_5_1_0_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_5_1_0_LC_10_19_1 .LUT_INIT=16'b0100000101010101;
    LogicCell40 \this_vga_signals.un16_address_g0_5_1_0_LC_10_19_1  (
            .in0(N__9090),
            .in1(N__9138),
            .in2(N__9018),
            .in3(N__18341),
            .lcout(\this_vga_signals.g0_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_c2_LC_10_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_c2_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_c2_LC_10_19_2 .LUT_INIT=16'b0111000111110101;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_c2_LC_10_19_2  (
            .in0(N__8103),
            .in1(N__7882),
            .in2(N__9015),
            .in3(N__7832),
            .lcout(\this_vga_signals.mult1_un47_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_0_0_LC_10_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_0_0_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_0_0_LC_10_19_3 .LUT_INIT=16'b0100000101010101;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_0_0_LC_10_19_3  (
            .in0(N__9089),
            .in1(N__9136),
            .in2(N__9017),
            .in3(N__18340),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_c2_LC_10_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_c2_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_c2_LC_10_19_4 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_c2_LC_10_19_4  (
            .in0(N__8105),
            .in1(N__7961),
            .in2(_gnd_net_),
            .in3(N__8001),
            .lcout(\this_vga_signals.mult1_un54_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_19_6 .LUT_INIT=16'b1000001000001010;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_19_6  (
            .in0(N__8104),
            .in1(N__7883),
            .in2(N__9016),
            .in3(N__7833),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_10_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_10_19_7 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_10_19_7  (
            .in0(N__9000),
            .in1(N__9137),
            .in2(N__7439),
            .in3(N__18339),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_i_3_LC_10_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_i_3_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_i_3_LC_10_20_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_i_3_LC_10_20_0  (
            .in0(N__8222),
            .in1(N__9790),
            .in2(N__7555),
            .in3(N__7512),
            .lcout(\this_vga_signals.rgb_1_2 ),
            .ltout(\this_vga_signals.rgb_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_10_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_10_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_10_20_1  (
            .in0(N__18336),
            .in1(N__8943),
            .in2(N__7436),
            .in3(N__7723),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_LC_10_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_LC_10_20_2 .LUT_INIT=16'b0001000101010000;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_LC_10_20_2  (
            .in0(N__8224),
            .in1(N__7433),
            .in2(N__7423),
            .in3(N__18335),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g3_0_2_LC_10_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g3_0_2_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g3_0_2_LC_10_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_g3_0_2_LC_10_20_3  (
            .in0(N__9792),
            .in1(N__7466),
            .in2(N__11463),
            .in3(N__8944),
            .lcout(),
            .ltout(\this_vga_signals.g3_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_19_LC_10_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_19_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_19_LC_10_20_4 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \this_vga_signals.un16_address_g0_19_LC_10_20_4  (
            .in0(N__7595),
            .in1(N__8003),
            .in2(N__7457),
            .in3(N__17310),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_3_c_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_18_LC_10_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_18_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_18_LC_10_20_5 .LUT_INIT=16'b0000010000001101;
    LogicCell40 \this_vga_signals.un16_address_g0_18_LC_10_20_5  (
            .in0(N__17311),
            .in1(N__7454),
            .in2(N__7448),
            .in3(N__7964),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABC21_LC_10_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABC21_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABC21_LC_10_20_6 .LUT_INIT=16'b1111100000000111;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABC21_LC_10_20_6  (
            .in0(N__8221),
            .in1(N__8289),
            .in2(N__9391),
            .in3(N__9732),
            .lcout(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABCZ0Z21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_axbxc3_LC_10_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_axbxc3_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_axbxc3_LC_10_20_7 .LUT_INIT=16'b1000101101000111;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_axbxc3_LC_10_20_7  (
            .in0(N__9791),
            .in1(N__7548),
            .in2(N__7519),
            .in3(N__8223),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIG8C01_LC_10_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIG8C01_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIG8C01_LC_10_21_0 .LUT_INIT=16'b0001100001100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIG8C01_LC_10_21_0  (
            .in0(N__8412),
            .in1(N__8326),
            .in2(N__9485),
            .in3(N__8461),
            .lcout(\this_vga_signals.d_N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_10_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_10_21_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_10_21_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_10_21_1  (
            .in0(N__8513),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18213),
            .ce(N__8676),
            .sr(N__8645));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_10_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_10_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_10_21_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__8581),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18213),
            .ce(N__8676),
            .sr(N__8645));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_21_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8534),
            .lcout(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18213),
            .ce(N__8676),
            .sr(N__8645));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_21_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8752),
            .lcout(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18213),
            .ce(N__8676),
            .sr(N__8645));
    defparam \this_vga_signals.un16_address_if_m13_ns_1_LC_10_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m13_ns_1_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m13_ns_1_LC_10_21_5 .LUT_INIT=16'b0000111101110111;
    LogicCell40 \this_vga_signals.un16_address_if_m13_ns_1_LC_10_21_5  (
            .in0(N__8462),
            .in1(N__7654),
            .in2(N__7574),
            .in3(N__8288),
            .lcout(),
            .ltout(\this_vga_signals.if_m13_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m13_ns_LC_10_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m13_ns_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m13_ns_LC_10_21_6 .LUT_INIT=16'b0000111101000100;
    LogicCell40 \this_vga_signals.un16_address_if_m13_ns_LC_10_21_6  (
            .in0(N__9390),
            .in1(N__7535),
            .in2(N__7562),
            .in3(N__18296),
            .lcout(\this_vga_signals.if_m13_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m6_LC_10_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m6_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m6_LC_10_21_7 .LUT_INIT=16'b0100100110010011;
    LogicCell40 \this_vga_signals.un16_address_if_m6_LC_10_21_7  (
            .in0(N__8327),
            .in1(N__9469),
            .in2(N__8291),
            .in3(N__8413),
            .lcout(\this_vga_signals.if_N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_ns_LC_10_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_ns_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_ns_LC_10_22_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_ns_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__14337),
            .in2(N__7475),
            .in3(N__7798),
            .lcout(\this_vga_signals.rgb_1_4 ),
            .ltout(\this_vga_signals.rgb_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIET844_LC_10_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIET844_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIET844_LC_10_22_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIET844_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__7529),
            .in2(N__7523),
            .in3(N__7496),
            .lcout(\this_vga_signals.M_vcounter_q_9_rep1_esr_RNIETZ0Z844 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_LC_10_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_LC_10_22_2 .LUT_INIT=16'b1001111011111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_LC_10_22_2  (
            .in0(N__8321),
            .in1(N__8411),
            .in2(N__8380),
            .in3(N__8453),
            .lcout(\this_vga_signals.d_N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_10_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_10_22_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_10_22_3  (
            .in0(N__8064),
            .in1(N__7604),
            .in2(N__8047),
            .in3(N__8020),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1 ),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_x1_LC_10_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_x1_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_x1_LC_10_22_4 .LUT_INIT=16'b1111001011100100;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_x1_LC_10_22_4  (
            .in0(N__9211),
            .in1(N__8362),
            .in2(N__7478),
            .in3(N__9697),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_i_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_N_2L1_LC_10_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_N_2L1_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_N_2L1_LC_10_22_5 .LUT_INIT=16'b0101111101001100;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_N_2L1_LC_10_22_5  (
            .in0(N__8063),
            .in1(N__7603),
            .in2(N__8046),
            .in3(N__8019),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_2_N_2L1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_LC_10_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_LC_10_22_6 .LUT_INIT=16'b1111011110001111;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_LC_10_22_6  (
            .in0(N__8320),
            .in1(N__8410),
            .in2(N__7607),
            .in3(N__8452),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_22_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_22_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_22_7  (
            .in0(N__8512),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18215),
            .ce(N__8677),
            .sr(N__8643));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_23_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8574),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18221),
            .ce(N__8679),
            .sr(N__8641));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_23_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_23_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_23_1  (
            .in0(N__8530),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18221),
            .ce(N__8679),
            .sr(N__8641));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_23_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8505),
            .lcout(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18221),
            .ce(N__8679),
            .sr(N__8641));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8550),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18221),
            .ce(N__8679),
            .sr(N__8641));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_10_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_10_23_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_10_23_4  (
            .in0(N__8551),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18221),
            .ce(N__8679),
            .sr(N__8641));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_10_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_10_23_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_10_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_10_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8529),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18221),
            .ce(N__8679),
            .sr(N__8641));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_24_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(N__11270),
            .in2(_gnd_net_),
            .in3(N__9874),
            .lcout(\this_vga_signals.un11_address_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA9V41_9_LC_10_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA9V41_9_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA9V41_9_LC_10_24_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIA9V41_9_LC_10_24_6  (
            .in0(N__9261),
            .in1(N__12258),
            .in2(_gnd_net_),
            .in3(N__9875),
            .lcout(\this_vga_signals.vsync_1_0_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNII2LG_7_LC_10_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNII2LG_7_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNII2LG_7_LC_10_24_7 .LUT_INIT=16'b0001000110001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNII2LG_7_LC_10_24_7  (
            .in0(N__7684),
            .in1(N__7672),
            .in2(_gnd_net_),
            .in3(N__8363),
            .lcout(\this_vga_signals.d_N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_11_1_LC_11_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_11_1_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_11_1_LC_11_17_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \this_vga_signals.un16_address_g0_11_1_LC_11_17_1  (
            .in0(N__9860),
            .in1(N__9406),
            .in2(N__11460),
            .in3(N__9143),
            .lcout(\this_vga_signals.g0_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_11_LC_11_17_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_11_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_11_LC_11_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vram.mem_radreg_11_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__20323),
            .in2(_gnd_net_),
            .in3(N__17168),
            .lcout(this_vram_mem_radreg_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18196),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_11_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_11_17_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__11428),
            .in2(_gnd_net_),
            .in3(N__9859),
            .lcout(),
            .ltout(\this_vga_signals.un11_address_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_6_0_LC_11_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_6_0_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_6_0_LC_11_17_7 .LUT_INIT=16'b1001000001010000;
    LogicCell40 \this_vga_signals.un16_address_g0_6_0_LC_11_17_7  (
            .in0(N__9019),
            .in1(N__7907),
            .in2(N__7637),
            .in3(N__7843),
            .lcout(\this_vga_signals.g0_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_11_LC_11_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_11_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_11_LC_11_18_0 .LUT_INIT=16'b1111110111011100;
    LogicCell40 \this_vga_signals.un16_address_g0_11_LC_11_18_0  (
            .in0(N__7634),
            .in1(N__9092),
            .in2(N__7628),
            .in3(N__18358),
            .lcout(),
            .ltout(\this_vga_signals.g2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g3_LC_11_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g3_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g3_LC_11_18_1 .LUT_INIT=16'b1001011000110011;
    LogicCell40 \this_vga_signals.un16_address_g3_LC_11_18_1  (
            .in0(N__7613),
            .in1(N__11169),
            .in2(N__7619),
            .in3(N__17102),
            .lcout(),
            .ltout(\this_vga_signals.g3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_0_i_a4_0_LC_11_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_0_i_a4_0_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_0_i_a4_0_LC_11_18_2 .LUT_INIT=16'b0000001000000001;
    LogicCell40 \this_vga_signals.un16_address_g0_0_i_a4_0_LC_11_18_2  (
            .in0(N__8804),
            .in1(N__12336),
            .in2(N__7616),
            .in3(N__11462),
            .lcout(\this_vga_signals.N_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g2_4_0_LC_11_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g2_4_0_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g2_4_0_LC_11_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un16_address_g2_4_0_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__11331),
            .in2(_gnd_net_),
            .in3(N__11504),
            .lcout(\this_vga_signals.g2_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_11_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_11_18_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_11_18_4  (
            .in0(N__7769),
            .in1(N__7703),
            .in2(_gnd_net_),
            .in3(N__17320),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g1_8_LC_11_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g1_8_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g1_8_LC_11_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un16_address_g1_8_LC_11_18_5  (
            .in0(N__12459),
            .in1(N__12140),
            .in2(_gnd_net_),
            .in3(N__11028),
            .lcout(\this_vga_signals.g1_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6 .LUT_INIT=16'b0110100101011010;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6  (
            .in0(N__11503),
            .in1(N__12508),
            .in2(N__11408),
            .in3(N__12548),
            .lcout(\this_vga_signals.mult1_un54_sum_i_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_x2_LC_11_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_x2_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_x2_LC_11_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un16_address_g0_i_x2_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__12139),
            .in2(N__7697),
            .in3(N__17101),
            .lcout(\this_vga_signals.g0_i_x2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_1_N_3L3_LC_11_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_1_N_3L3_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_1_N_3L3_LC_11_19_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un16_address_g0_1_N_3L3_LC_11_19_0  (
            .in0(N__11505),
            .in1(N__17118),
            .in2(_gnd_net_),
            .in3(N__10899),
            .lcout(\this_vga_signals.g0_1_N_3L3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_11_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_11_19_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_11_19_1  (
            .in0(N__9835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8237),
            .lcout(),
            .ltout(\this_vga_signals.un11_address_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_5_1_LC_11_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_5_1_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_5_1_LC_11_19_2 .LUT_INIT=16'b1001000001010000;
    LogicCell40 \this_vga_signals.un16_address_g0_5_1_LC_11_19_2  (
            .in0(N__9013),
            .in1(N__7906),
            .in2(N__7694),
            .in3(N__7844),
            .lcout(\this_vga_signals.g0_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_x0_3_LC_11_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_x0_3_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_x0_3_LC_11_19_3 .LUT_INIT=16'b0110001100111001;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_x0_3_LC_11_19_3  (
            .in0(N__7963),
            .in1(N__7750),
            .in2(N__7985),
            .in3(N__17299),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_i_x0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_ns_3_LC_11_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_ns_3_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_ns_3_LC_11_19_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_ns_3_LC_11_19_4  (
            .in0(N__17300),
            .in1(N__7751),
            .in2(N__7691),
            .in3(N__7942),
            .lcout(this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_c_LC_11_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_c_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_c_LC_11_19_5 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_c_LC_11_19_5  (
            .in0(N__8102),
            .in1(N__7765),
            .in2(N__17319),
            .in3(N__8002),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_3_c ),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_3_c_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_19_6 .LUT_INIT=16'b0000010000001101;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_19_6  (
            .in0(N__17298),
            .in1(N__7984),
            .in2(N__7967),
            .in3(N__7962),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_1_N_5L8_LC_11_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_1_N_5L8_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_1_N_5L8_LC_11_19_7 .LUT_INIT=16'b0001000001010001;
    LogicCell40 \this_vga_signals.un16_address_g0_1_N_5L8_LC_11_19_7  (
            .in0(N__7943),
            .in1(N__7934),
            .in2(N__7922),
            .in3(N__17301),
            .lcout(\this_vga_signals.g0_1_N_5L8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb2_0_LC_11_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb2_0_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb2_0_LC_11_20_0 .LUT_INIT=16'b0110100111000011;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb2_0_LC_11_20_0  (
            .in0(N__7898),
            .in1(N__8090),
            .in2(N__9020),
            .in3(N__7834),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_axb1_LC_11_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_axb1_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_axb1_LC_11_20_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_axb1_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__8119),
            .in2(_gnd_net_),
            .in3(N__8894),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un40_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_11_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_11_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_11_20_3  (
            .in0(N__9011),
            .in1(N__7730),
            .in2(N__7754),
            .in3(N__18337),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_5_LC_11_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_5_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_5_LC_11_20_4 .LUT_INIT=16'b1100001101101001;
    LogicCell40 \this_vga_signals.un16_address_g0_5_LC_11_20_4  (
            .in0(N__7739),
            .in1(N__11496),
            .in2(N__11457),
            .in3(N__12509),
            .lcout(\this_vga_signals.if_N_13_i_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_11_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_11_20_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_11_20_5  (
            .in0(N__9010),
            .in1(N__7729),
            .in2(N__17318),
            .in3(N__18338),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_1_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_11_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_11_20_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_11_20_6  (
            .in0(N__7712),
            .in1(_gnd_net_),
            .in2(N__7706),
            .in3(N__9135),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_35_LC_11_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_35_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_35_LC_11_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un16_address_g0_35_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(N__11413),
            .in2(N__8147),
            .in3(N__12297),
            .lcout(\this_vga_signals.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIL7SG_4_LC_11_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIL7SG_4_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIL7SG_4_LC_11_21_0 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIL7SG_4_LC_11_21_0  (
            .in0(N__8066),
            .in1(N__8325),
            .in2(N__8290),
            .in3(N__8460),
            .lcout(\this_vga_signals.un11_address_c4_i ),
            .ltout(\this_vga_signals.un11_address_c4_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_1_LC_11_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_1_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_1_LC_11_21_1 .LUT_INIT=16'b0110010101101001;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_1_LC_11_21_1  (
            .in0(N__8091),
            .in1(N__9475),
            .in2(N__8132),
            .in3(N__8474),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_5_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_LC_11_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_LC_11_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_LC_11_21_2  (
            .in0(N__8125),
            .in1(N__8891),
            .in2(N__8129),
            .in3(N__18303),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_5_4 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_5_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_LC_11_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_LC_11_21_3 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_LC_11_21_3  (
            .in0(N__8892),
            .in1(N__8126),
            .in2(N__8108),
            .in3(N__8986),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_21_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_21_4  (
            .in0(N__8280),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8218),
            .lcout(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_21_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8701),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18208),
            .ce(N__8678),
            .sr(N__8644));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_21_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_21_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_21_6  (
            .in0(N__8700),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18208),
            .ce(N__8678),
            .sr(N__8644));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_5_LC_11_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_5_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_5_LC_11_21_7 .LUT_INIT=16'b0000000000111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_5_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__8065),
            .in2(N__8048),
            .in3(N__8021),
            .lcout(\this_vga_signals.SUM_2_i_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_0_LC_11_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_0_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_0_LC_11_22_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_0_LC_11_22_0  (
            .in0(N__8323),
            .in1(N__8367),
            .in2(N__8414),
            .in3(N__8446),
            .lcout(\this_vga_signals.SUM_2_i_a4_a0_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJK9S_8_LC_11_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJK9S_8_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJK9S_8_LC_11_22_1 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIJK9S_8_LC_11_22_1  (
            .in0(N__9465),
            .in1(N__8486),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\this_vga_signals.SUM_2_i_a4_1_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIJ3MB6_LC_11_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIJ3MB6_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIJ3MB6_LC_11_22_2 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIJ3MB6_LC_11_22_2  (
            .in0(N__8473),
            .in1(N__8165),
            .in2(N__8480),
            .in3(N__8153),
            .lcout(\this_vga_signals.SUM_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIHIQV_LC_11_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIHIQV_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIHIQV_LC_11_22_3 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIHIQV_LC_11_22_3  (
            .in0(N__8447),
            .in1(_gnd_net_),
            .in2(N__8379),
            .in3(N__8324),
            .lcout(),
            .ltout(\this_vga_signals.un11_address_c5_a0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPM1_LC_11_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPM1_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPM1_LC_11_22_4 .LUT_INIT=16'b1000111101110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPM1_LC_11_22_4  (
            .in0(N__8281),
            .in1(N__8220),
            .in2(N__8477),
            .in3(N__9257),
            .lcout(\this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPMZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_1_LC_11_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_1_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_1_LC_11_22_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_1_LC_11_22_5  (
            .in0(N__8448),
            .in1(N__8409),
            .in2(N__8378),
            .in3(N__8322),
            .lcout(\this_vga_signals.SUM_2_i_a4_0_a0_2_3 ),
            .ltout(\this_vga_signals.SUM_2_i_a4_0_a0_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUK2_LC_11_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUK2_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUK2_LC_11_22_6 .LUT_INIT=16'b0111011101110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUK2_LC_11_22_6  (
            .in0(N__8282),
            .in1(N__8219),
            .in2(N__8174),
            .in3(N__8171),
            .lcout(\this_vga_signals.SUM_2_i_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_9_LC_11_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_9_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_9_LC_11_22_7 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_9_LC_11_22_7  (
            .in0(N__9258),
            .in1(N__9709),
            .in2(N__9484),
            .in3(N__8159),
            .lcout(\this_vga_signals.SUM_2_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_11_23_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_11_23_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_11_23_0  (
            .in0(N__11686),
            .in1(N__9901),
            .in2(N__9575),
            .in3(N__9574),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__18216),
            .ce(),
            .sr(N__8640));
    defparam \this_vga_signals.M_vcounter_q_1_LC_11_23_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_11_23_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_11_23_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_11_23_1  (
            .in0(N__11688),
            .in1(N__12441),
            .in2(_gnd_net_),
            .in3(N__8597),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__18216),
            .ce(),
            .sr(N__8640));
    defparam \this_vga_signals.M_vcounter_q_2_LC_11_23_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_11_23_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_11_23_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_11_23_2  (
            .in0(N__11687),
            .in1(N__12108),
            .in2(_gnd_net_),
            .in3(N__8594),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__18216),
            .ce(),
            .sr(N__8640));
    defparam \this_vga_signals.M_vcounter_q_3_LC_11_23_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_11_23_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_11_23_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_11_23_3  (
            .in0(N__11689),
            .in1(N__12257),
            .in2(_gnd_net_),
            .in3(N__8591),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__18216),
            .ce(),
            .sr(N__8640));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_11_23_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_11_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(N__11289),
            .in2(_gnd_net_),
            .in3(N__8588),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_11_23_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_11_23_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9873),
            .in3(N__8561),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_11_23_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_11_23_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9410),
            .in3(N__8537),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_11_23_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_11_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_11_23_7  (
            .in0(_gnd_net_),
            .in1(N__9721),
            .in2(_gnd_net_),
            .in3(N__8516),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_11_24_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_11_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_11_24_0  (
            .in0(_gnd_net_),
            .in1(N__9497),
            .in2(_gnd_net_),
            .in3(N__8489),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_11_24_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_11_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_11_24_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_11_24_1  (
            .in0(_gnd_net_),
            .in1(N__9259),
            .in2(_gnd_net_),
            .in3(N__8756),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIAA7K1_9_LC_11_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIAA7K1_9_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIAA7K1_9_LC_11_24_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIAA7K1_9_LC_11_24_6  (
            .in0(N__8708),
            .in1(N__10702),
            .in2(N__10778),
            .in3(N__10741),
            .lcout(N_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIC1AR_4_LC_11_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIC1AR_4_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIC1AR_4_LC_11_24_7 .LUT_INIT=16'b0111011111101110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIC1AR_4_LC_11_24_7  (
            .in0(N__10511),
            .in1(N__10639),
            .in2(_gnd_net_),
            .in3(N__10595),
            .lcout(\this_vga_signals.hsync_1_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_11_25_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_11_25_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_11_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_11_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8702),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18223),
            .ce(N__8681),
            .sr(N__8639));
    defparam \this_vga_signals.rgb_cnst_i_o2_0_4_LC_12_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.rgb_cnst_i_o2_0_4_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.rgb_cnst_i_o2_0_4_LC_12_16_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.rgb_cnst_i_o2_0_4_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__13750),
            .in2(N__10410),
            .in3(N__12959),
            .lcout(\this_vga_signals.N_381_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.rgb_cnst_i_a5_0_4_LC_12_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.rgb_cnst_i_a5_0_4_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.rgb_cnst_i_a5_0_4_LC_12_16_1 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \this_vga_signals.rgb_cnst_i_a5_0_4_LC_12_16_1  (
            .in0(N__15881),
            .in1(N__10392),
            .in2(N__13769),
            .in3(N__12958),
            .lcout(),
            .ltout(\this_vga_signals.N_390_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIS1MK91_9_LC_12_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIS1MK91_9_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIS1MK91_9_LC_12_16_2 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIS1MK91_9_LC_12_16_2  (
            .in0(N__20324),
            .in1(N__8609),
            .in2(N__8603),
            .in3(N__15880),
            .lcout(\this_vga_signals.N_371_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_0_9_LC_12_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_0_9_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_0_9_LC_12_17_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_0_9_LC_12_17_0  (
            .in0(N__10376),
            .in1(N__12987),
            .in2(N__13770),
            .in3(N__20289),
            .lcout(),
            .ltout(\this_vga_signals.rgb_cnst_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIO6OD01_9_LC_12_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIO6OD01_9_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIO6OD01_9_LC_12_17_1 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIO6OD01_9_LC_12_17_1  (
            .in0(N__12986),
            .in1(N__13751),
            .in2(N__8600),
            .in3(N__15902),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_esr_RNIO6OD01Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR0T9KU3_9_LC_12_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR0T9KU3_9_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR0T9KU3_9_LC_12_17_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIR0T9KU3_9_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__14077),
            .in2(N__8831),
            .in3(N__12908),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_x2_5_LC_12_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_x2_5_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_x2_5_LC_12_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un16_address_g0_i_x2_5_LC_12_18_0  (
            .in0(N__16083),
            .in1(N__16121),
            .in2(N__8816),
            .in3(N__8795),
            .lcout(\this_vga_signals.g0_i_x2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_o2_1_x2_LC_12_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_o2_1_x2_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_o2_1_x2_LC_12_18_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un16_address_g0_i_o2_1_x2_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10914),
            .in3(N__10964),
            .lcout(\this_vga_signals.N_10_i ),
            .ltout(\this_vga_signals.N_10_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_x2_5_1_LC_12_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_x2_5_1_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_x2_5_1_LC_12_18_2 .LUT_INIT=16'b0110010110100110;
    LogicCell40 \this_vga_signals.un16_address_g0_i_x2_5_1_LC_12_18_2  (
            .in0(N__17116),
            .in1(N__12335),
            .in2(N__8798),
            .in3(N__11451),
            .lcout(\this_vga_signals.g0_i_x2_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g4_0_0_LC_12_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g4_0_0_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g4_0_0_LC_12_18_3 .LUT_INIT=16'b1110110111011110;
    LogicCell40 \this_vga_signals.un16_address_g4_0_0_LC_12_18_3  (
            .in0(N__10906),
            .in1(N__12332),
            .in2(N__11465),
            .in3(N__10966),
            .lcout(),
            .ltout(\this_vga_signals.g4_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g4_1_LC_12_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g4_1_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g4_1_LC_12_18_4 .LUT_INIT=16'b1111001011111101;
    LogicCell40 \this_vga_signals.un16_address_g4_1_LC_12_18_4  (
            .in0(N__17117),
            .in1(N__8789),
            .in2(N__8780),
            .in3(N__11144),
            .lcout(\this_vga_signals.g4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_0_N_5L7_LC_12_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_0_N_5L7_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_0_N_5L7_LC_12_18_5 .LUT_INIT=16'b0100000000100000;
    LogicCell40 \this_vga_signals.un16_address_g0_i_0_N_5L7_LC_12_18_5  (
            .in0(N__8777),
            .in1(N__8768),
            .in2(N__12170),
            .in3(N__16082),
            .lcout(\this_vga_signals.g0_i_0_N_5L7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_x2_0_LC_12_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_x2_0_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_x2_0_LC_12_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un16_address_g0_i_x2_0_LC_12_18_6  (
            .in0(N__12331),
            .in1(N__11450),
            .in2(_gnd_net_),
            .in3(N__10902),
            .lcout(\this_vga_signals.g0_i_x2_1_1 ),
            .ltout(\this_vga_signals.g0_i_x2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_x1_LC_12_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_x1_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_x1_LC_12_18_7 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \this_vga_signals.un16_address_g0_i_x1_LC_12_18_7  (
            .in0(N__11143),
            .in1(N__10965),
            .in2(N__8759),
            .in3(N__17115),
            .lcout(\this_vga_signals.g0_i_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_12_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_12_19_0 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17158),
            .in3(N__11147),
            .lcout(this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1),
            .ltout(this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_0_i_a4_LC_12_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_0_i_a4_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_0_i_a4_LC_12_19_1 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \this_vga_signals.un16_address_g0_0_i_a4_LC_12_19_1  (
            .in0(N__12333),
            .in1(N__9149),
            .in2(N__8861),
            .in3(N__16057),
            .lcout(\this_vga_signals.N_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_x0_LC_12_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_x0_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_x0_LC_12_19_2 .LUT_INIT=16'b0010100000010100;
    LogicCell40 \this_vga_signals.un16_address_g0_i_x0_LC_12_19_2  (
            .in0(N__10967),
            .in1(N__11148),
            .in2(N__17159),
            .in3(N__8858),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_ns_LC_12_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_ns_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_ns_LC_12_19_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.un16_address_g0_i_ns_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__8852),
            .in2(N__8846),
            .in3(N__16056),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g1_1_1_a3_LC_12_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g1_1_1_a3_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g1_1_1_a3_LC_12_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un16_address_g1_1_1_a3_LC_12_19_4  (
            .in0(N__10968),
            .in1(N__11455),
            .in2(_gnd_net_),
            .in3(N__10900),
            .lcout(\this_vga_signals.g1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m3_4_LC_12_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m3_4_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m3_4_LC_12_19_5 .LUT_INIT=16'b1111001100110000;
    LogicCell40 \this_vga_signals.un16_address_if_m3_4_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__17103),
            .in2(N__11005),
            .in3(N__11027),
            .lcout(this_vga_signals_un16_address_if_i1_mux_0),
            .ltout(this_vga_signals_un16_address_if_i1_mux_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_x2_0_i_o3_LC_12_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_x2_0_i_o3_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_x2_0_i_o3_LC_12_19_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un16_address_g0_i_x2_0_i_o3_LC_12_19_6  (
            .in0(N__17110),
            .in1(_gnd_net_),
            .in2(N__8843),
            .in3(N__11149),
            .lcout(\this_vga_signals.N_6_i ),
            .ltout(\this_vga_signals.N_6_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g1_0_a3_LC_12_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g1_0_a3_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g1_0_a3_LC_12_19_7 .LUT_INIT=16'b1011001001001101;
    LogicCell40 \this_vga_signals.un16_address_g1_0_a3_LC_12_19_7  (
            .in0(N__12334),
            .in1(N__12168),
            .in2(N__8840),
            .in3(N__8837),
            .lcout(\this_vga_signals.g1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_20_0 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_20_0  (
            .in0(N__10883),
            .in1(_gnd_net_),
            .in2(N__10971),
            .in3(N__11437),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m5_0_LC_12_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m5_0_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m5_0_LC_12_20_1 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un16_address_if_m5_0_LC_12_20_1  (
            .in0(N__12304),
            .in1(N__10880),
            .in2(N__11461),
            .in3(N__10949),
            .lcout(\this_vga_signals.if_N_1_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_0_i_x2_1_LC_12_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_0_i_x2_1_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_0_i_x2_1_LC_12_20_2 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un16_address_g0_0_i_x2_1_LC_12_20_2  (
            .in0(N__10882),
            .in1(_gnd_net_),
            .in2(N__10970),
            .in3(N__11436),
            .lcout(\this_vga_signals.N_11_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_25_1_LC_12_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_25_1_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_25_1_LC_12_20_3 .LUT_INIT=16'b0000100110011111;
    LogicCell40 \this_vga_signals.un16_address_g0_25_1_LC_12_20_3  (
            .in0(N__9012),
            .in1(N__9142),
            .in2(N__9110),
            .in3(N__18359),
            .lcout(),
            .ltout(\this_vga_signals.g0_25_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_25_LC_12_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_25_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_25_LC_12_20_4 .LUT_INIT=16'b1001100101101001;
    LogicCell40 \this_vga_signals.un16_address_g0_25_LC_12_20_4  (
            .in0(N__9101),
            .in1(N__8870),
            .in2(N__9095),
            .in3(N__9091),
            .lcout(),
            .ltout(\this_vga_signals.if_N_13_i_i_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_9_LC_12_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_9_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_9_LC_12_20_5 .LUT_INIT=16'b1000001010001000;
    LogicCell40 \this_vga_signals.un16_address_g0_9_LC_12_20_5  (
            .in0(N__9050),
            .in1(N__11190),
            .in2(N__9053),
            .in3(N__17132),
            .lcout(\this_vga_signals.g2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g2_0_LC_12_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g2_0_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g2_0_LC_12_20_6 .LUT_INIT=16'b0001001000100001;
    LogicCell40 \this_vga_signals.un16_address_g2_0_LC_12_20_6  (
            .in0(N__10881),
            .in1(N__12305),
            .in2(N__10969),
            .in3(N__11435),
            .lcout(\this_vga_signals.g2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVRQGTU3_9_LC_12_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVRQGTU3_9_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVRQGTU3_9_LC_12_21_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIVRQGTU3_9_LC_12_21_1  (
            .in0(N__14090),
            .in1(N__13082),
            .in2(_gnd_net_),
            .in3(N__9044),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_12_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_12_21_5 .LUT_INIT=16'b1110110000010011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_12_21_5  (
            .in0(N__9861),
            .in1(N__9405),
            .in2(N__11418),
            .in3(N__9742),
            .lcout(),
            .ltout(\this_vga_signals.un11_address_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_3_0_LC_12_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_3_0_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_3_0_LC_12_21_6 .LUT_INIT=16'b0110010110100110;
    LogicCell40 \this_vga_signals.un16_address_g0_3_0_LC_12_21_6  (
            .in0(N__11348),
            .in1(N__9014),
            .in2(N__8897),
            .in3(N__8893),
            .lcout(\this_vga_signals.g0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_12_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_12_22_0 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_12_22_0  (
            .in0(N__12440),
            .in1(N__9897),
            .in2(N__12138),
            .in3(N__12247),
            .lcout(),
            .ltout(\this_vga_signals.N_28_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_8_LC_12_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_8_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_8_LC_12_22_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_8_LC_12_22_1  (
            .in0(N__9650),
            .in1(N__9404),
            .in2(N__9521),
            .in3(N__9496),
            .lcout(),
            .ltout(\this_vga_signals.N_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVV6F6_9_LC_12_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVV6F6_9_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVV6F6_9_LC_12_22_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIVV6F6_9_LC_12_22_2  (
            .in0(N__11660),
            .in1(N__9570),
            .in2(N__9518),
            .in3(N__9263),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNIVV6F6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clock.M_counter_q_1_LC_12_22_3 .C_ON=1'b0;
    defparam \this_pixel_clock.M_counter_q_1_LC_12_22_3 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clock.M_counter_q_1_LC_12_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_pixel_clock.M_counter_q_1_LC_12_22_3  (
            .in0(N__15257),
            .in1(N__13040),
            .in2(_gnd_net_),
            .in3(N__9550),
            .lcout(\this_pixel_clock.M_counter_q_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18209),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_22_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(N__9495),
            .in2(_gnd_net_),
            .in3(N__9743),
            .lcout(),
            .ltout(\this_vga_signals.rgb297_i_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_22_5 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_22_5  (
            .in0(N__11406),
            .in1(N__9862),
            .in2(N__9413),
            .in3(N__9403),
            .lcout(\this_vga_signals.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI38HR1_5_LC_12_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI38HR1_5_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI38HR1_5_LC_12_22_6 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI38HR1_5_LC_12_22_6  (
            .in0(N__9863),
            .in1(N__9287),
            .in2(_gnd_net_),
            .in3(N__11407),
            .lcout(\this_vga_signals.CO0_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clock.M_counter_q_RNIJR071_1_LC_12_22_7 .C_ON=1'b0;
    defparam \this_pixel_clock.M_counter_q_RNIJR071_1_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \this_pixel_clock.M_counter_q_RNIJR071_1_LC_12_22_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_pixel_clock.M_counter_q_RNIJR071_1_LC_12_22_7  (
            .in0(N__15256),
            .in1(N__13039),
            .in2(_gnd_net_),
            .in3(N__9549),
            .lcout(M_counter_q_RNIJR071_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_12_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_12_23_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_12_23_1  (
            .in0(N__10772),
            .in1(N__10705),
            .in2(_gnd_net_),
            .in3(N__10739),
            .lcout(\this_vga_signals.N_33_0 ),
            .ltout(\this_vga_signals.N_33_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICLUO4_9_LC_12_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICLUO4_9_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICLUO4_9_LC_12_23_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICLUO4_9_LC_12_23_2  (
            .in0(N__9262),
            .in1(N__9163),
            .in2(N__9152),
            .in3(N__9589),
            .lcout(\this_vga_signals.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_23_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_23_5  (
            .in0(N__10637),
            .in1(N__10738),
            .in2(_gnd_net_),
            .in3(N__10593),
            .lcout(),
            .ltout(\this_vga_signals.N_45_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_23_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_23_6  (
            .in0(N__10706),
            .in1(_gnd_net_),
            .in2(N__9578),
            .in3(N__10773),
            .lcout(N_23_0),
            .ltout(N_23_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clock.M_counter_q_RNIQR4I2_1_LC_12_23_7 .C_ON=1'b0;
    defparam \this_pixel_clock.M_counter_q_RNIQR4I2_1_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \this_pixel_clock.M_counter_q_RNIQR4I2_1_LC_12_23_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_pixel_clock.M_counter_q_RNIQR4I2_1_LC_12_23_7  (
            .in0(N__15306),
            .in1(N__13038),
            .in2(N__9554),
            .in3(N__9551),
            .lcout(M_counter_q_RNIQR4I2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_24_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__11747),
            .in2(N__11618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_24_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_24_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_24_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_12_24_1  (
            .in0(N__11702),
            .in1(N__10325),
            .in2(_gnd_net_),
            .in3(N__9536),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__18217),
            .ce(),
            .sr(N__11582));
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_24_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_24_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_24_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_12_24_2  (
            .in0(N__11699),
            .in1(N__10548),
            .in2(_gnd_net_),
            .in3(N__9533),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__18217),
            .ce(),
            .sr(N__11582));
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_24_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_24_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_24_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_12_24_3  (
            .in0(N__11703),
            .in1(N__10510),
            .in2(_gnd_net_),
            .in3(N__9530),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__18217),
            .ce(),
            .sr(N__11582));
    defparam \this_vga_signals.M_hcounter_q_5_LC_12_24_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_12_24_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_12_24_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_12_24_4  (
            .in0(N__11700),
            .in1(N__10638),
            .in2(_gnd_net_),
            .in3(N__9527),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__18217),
            .ce(),
            .sr(N__11582));
    defparam \this_vga_signals.M_hcounter_q_6_LC_12_24_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_12_24_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_12_24_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_12_24_5  (
            .in0(N__11704),
            .in1(N__10594),
            .in2(_gnd_net_),
            .in3(N__9524),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__18217),
            .ce(),
            .sr(N__11582));
    defparam \this_vga_signals.M_hcounter_q_7_LC_12_24_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_12_24_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_12_24_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_12_24_6  (
            .in0(N__11701),
            .in1(N__10740),
            .in2(_gnd_net_),
            .in3(N__9638),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__18217),
            .ce(),
            .sr(N__11582));
    defparam \this_vga_signals.M_hcounter_q_8_LC_12_24_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_12_24_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_12_24_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_12_24_7  (
            .in0(N__11705),
            .in1(N__10774),
            .in2(_gnd_net_),
            .in3(N__9635),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__18217),
            .ce(),
            .sr(N__11582));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_12_25_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_12_25_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_12_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(N__10701),
            .in2(_gnd_net_),
            .in3(N__9632),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18222),
            .ce(N__10466),
            .sr(N__11577));
    defparam \this_vga_signals.un16_address_g0_10_LC_13_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_10_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_10_LC_13_18_0 .LUT_INIT=16'b0001010010000010;
    LogicCell40 \this_vga_signals.un16_address_g0_10_LC_13_18_0  (
            .in0(N__16060),
            .in1(N__16136),
            .in2(N__12365),
            .in3(N__12055),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_30_LC_13_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_30_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_30_LC_13_18_1 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \this_vga_signals.un16_address_g0_30_LC_13_18_1  (
            .in0(N__12178),
            .in1(N__9629),
            .in2(N__9620),
            .in3(N__9617),
            .lcout(\this_vga_signals.N_9_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m2_0_LC_13_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m2_0_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m2_0_LC_13_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_if_m2_0_LC_13_18_2  (
            .in0(N__16058),
            .in1(N__11183),
            .in2(N__12364),
            .in3(N__17181),
            .lcout(\this_vga_signals.if_N_3_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_x2_1_LC_13_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_x2_1_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_x2_1_LC_13_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_g0_i_x2_1_LC_13_18_3  (
            .in0(N__9611),
            .in1(N__16059),
            .in2(N__16146),
            .in3(N__10802),
            .lcout(\this_vga_signals.g0_i_x2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_1_0_LC_13_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_1_0_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_1_0_LC_13_18_5 .LUT_INIT=16'b0100000100101000;
    LogicCell40 \this_vga_signals.un16_address_g0_1_0_LC_13_18_5  (
            .in0(N__12056),
            .in1(N__12356),
            .in2(N__16147),
            .in3(N__16061),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_LC_13_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_LC_13_18_6 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \this_vga_signals.un16_address_g0_LC_13_18_6  (
            .in0(N__12180),
            .in1(N__9602),
            .in2(N__9596),
            .in3(N__11077),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_i_LC_13_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_i_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_i_LC_13_18_7 .LUT_INIT=16'b1000001000010100;
    LogicCell40 \this_vga_signals.un16_address_g0_i_i_LC_13_18_7  (
            .in0(N__12179),
            .in1(N__10112),
            .in2(N__10106),
            .in3(N__12475),
            .lcout(\this_vga_signals.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_7_LC_13_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_7_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_7_LC_13_19_0 .LUT_INIT=16'b1111000010011001;
    LogicCell40 \this_vga_signals.un16_address_g0_7_LC_13_19_0  (
            .in0(N__10103),
            .in1(N__9911),
            .in2(N__10097),
            .in3(N__9938),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3CNE3O2_9_LC_13_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3CNE3O2_9_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3CNE3O2_9_LC_13_19_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI3CNE3O2_9_LC_13_19_1  (
            .in0(N__20291),
            .in1(N__10085),
            .in2(N__10079),
            .in3(N__10808),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_0_N_4L5_LC_13_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_0_N_4L5_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_0_N_4L5_LC_13_19_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.un16_address_g0_i_0_N_4L5_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__9959),
            .in2(_gnd_net_),
            .in3(N__11076),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_0_N_4L5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_0_LC_13_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_0_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_0_LC_13_19_3 .LUT_INIT=16'b0010001010000010;
    LogicCell40 \this_vga_signals.un16_address_g0_i_0_LC_13_19_3  (
            .in0(N__9881),
            .in1(N__9953),
            .in2(N__9947),
            .in3(N__9944),
            .lcout(\this_vga_signals.if_i4_mux_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g1_7_LC_13_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g1_7_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g1_7_LC_13_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_g1_7_LC_13_19_4  (
            .in0(N__10838),
            .in1(N__9932),
            .in2(N__9926),
            .in3(N__17164),
            .lcout(\this_vga_signals.g1_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_0_N_2L1_LC_13_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_0_N_2L1_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_0_N_2L1_LC_13_20_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un16_address_g0_i_0_N_2L1_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__12460),
            .in2(_gnd_net_),
            .in3(N__9905),
            .lcout(\this_vga_signals.g0_i_0_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIU721_7_LC_13_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIU721_7_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIU721_7_LC_13_20_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIU721_7_LC_13_20_2  (
            .in0(N__11438),
            .in1(N__9867),
            .in2(_gnd_net_),
            .in3(N__9741),
            .lcout(\this_vga_signals.M_vcounter_d_1_sqmuxa_i_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI39EPS4_9_LC_13_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI39EPS4_9_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI39EPS4_9_LC_13_22_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI39EPS4_9_LC_13_22_0  (
            .in0(N__10124),
            .in1(N__10142),
            .in2(N__20290),
            .in3(N__10130),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_m1_LC_13_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_m1_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_m1_LC_13_22_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un4_address_if_m1_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__10330),
            .in2(_gnd_net_),
            .in3(N__20148),
            .lcout(\this_vga_signals.mult1_un82_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_m7_0_x4_LC_13_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_m7_0_x4_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_m7_0_x4_LC_13_22_2 .LUT_INIT=16'b0110101001010110;
    LogicCell40 \this_vga_signals.un4_address_if_m7_0_x4_LC_13_22_2  (
            .in0(N__10277),
            .in1(N__10331),
            .in2(N__17779),
            .in3(N__10551),
            .lcout(),
            .ltout(\this_vga_signals.if_N_8_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_m7_0_m2_LC_13_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_m7_0_m2_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_m7_0_m2_LC_13_22_3 .LUT_INIT=16'b0011001110001110;
    LogicCell40 \this_vga_signals.un4_address_if_m7_0_m2_LC_13_22_3  (
            .in0(N__11610),
            .in1(N__11746),
            .in2(N__10151),
            .in3(N__10148),
            .lcout(\this_vga_signals.mult1_un89_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_m7_0_m2_0_LC_13_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_m7_0_m2_0_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_m7_0_m2_0_LC_13_22_4 .LUT_INIT=16'b0000100101101111;
    LogicCell40 \this_vga_signals.un4_address_if_m7_0_m2_0_LC_13_22_4  (
            .in0(N__17769),
            .in1(N__10549),
            .in2(N__10334),
            .in3(N__10283),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_13_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_13_22_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_13_22_5  (
            .in0(N__10550),
            .in1(N__17770),
            .in2(N__10136),
            .in3(N__10276),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0 ),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_13_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_13_22_6 .LUT_INIT=16'b1110000101111000;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_13_22_6  (
            .in0(N__17774),
            .in1(N__10333),
            .in2(N__10133),
            .in3(N__10552),
            .lcout(\this_vga_signals.mult1_un89_sum_axbxc3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_c2_LC_13_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_c2_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_c2_LC_13_22_7 .LUT_INIT=16'b0010001010111011;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_c2_LC_13_22_7  (
            .in0(N__10332),
            .in1(N__11745),
            .in2(_gnd_net_),
            .in3(N__20149),
            .lcout(\this_vga_signals.mult1_un82_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_13_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_13_23_0 .LUT_INIT=16'b0010101111010100;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_13_23_0  (
            .in0(N__10553),
            .in1(N__17775),
            .in2(N__10326),
            .in3(N__10118),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un54_sum_c3_LC_13_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un54_sum_c3_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un54_sum_c3_LC_13_23_1 .LUT_INIT=16'b0101110101000101;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un54_sum_c3_LC_13_23_1  (
            .in0(N__10664),
            .in1(N__10655),
            .in2(N__10640),
            .in3(N__10592),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_23_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__10636),
            .in2(N__10349),
            .in3(N__10508),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axbxc3_LC_13_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axbxc3_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axbxc3_LC_13_23_3 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axbxc3_LC_13_23_3  (
            .in0(N__11901),
            .in1(N__11871),
            .in2(N__10346),
            .in3(N__10475),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_c3_LC_13_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_c3_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_c3_LC_13_23_4 .LUT_INIT=16'b1100110001110001;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_c3_LC_13_23_4  (
            .in0(N__10309),
            .in1(N__10535),
            .in2(N__10343),
            .in3(N__10275),
            .lcout(\this_vga_signals.mult1_un75_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_13_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_13_23_5 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_13_23_5  (
            .in0(N__11872),
            .in1(N__10340),
            .in2(N__11903),
            .in3(N__10474),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_m7_0_o4_1_LC_13_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_m7_0_o4_1_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_m7_0_o4_1_LC_13_23_6 .LUT_INIT=16'b0001011101110001;
    LogicCell40 \this_vga_signals.un4_address_if_m7_0_o4_1_LC_13_23_6  (
            .in0(N__10308),
            .in1(N__11736),
            .in2(N__10286),
            .in3(N__10274),
            .lcout(\this_vga_signals.if_N_9_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axb1_LC_13_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axb1_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axb1_LC_13_23_7 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axb1_LC_13_23_7  (
            .in0(N__10509),
            .in1(N__11897),
            .in2(_gnd_net_),
            .in3(N__11870),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_13_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_13_24_0 .LUT_INIT=16'b1101010111010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_13_24_0  (
            .in0(N__10771),
            .in1(N__10737),
            .in2(N__10704),
            .in3(N__10591),
            .lcout(\this_vga_signals.SUM_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_13_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_13_24_1 .LUT_INIT=16'b1100000101111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_13_24_1  (
            .in0(N__10588),
            .in1(N__10689),
            .in2(N__10742),
            .in3(N__10769),
            .lcout(\this_vga_signals.SUM_3 ),
            .ltout(\this_vga_signals.SUM_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_13_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_13_24_2 .LUT_INIT=16'b1100011111111111;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_13_24_2  (
            .in0(N__10506),
            .in1(N__10631),
            .in2(N__10781),
            .in3(N__10589),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_13_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_13_24_4 .LUT_INIT=16'b1011110101000010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_13_24_4  (
            .in0(N__10770),
            .in1(N__10733),
            .in2(N__10703),
            .in3(N__10587),
            .lcout(\this_vga_signals.N_34 ),
            .ltout(\this_vga_signals.N_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_24_5 .LUT_INIT=16'b0001011100011111;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_24_5  (
            .in0(N__10630),
            .in1(N__10505),
            .in2(N__10658),
            .in3(N__10653),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_24_6 .LUT_INIT=16'b1111100011100000;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_24_6  (
            .in0(N__10654),
            .in1(N__10632),
            .in2(N__10598),
            .in3(N__10590),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_c2_0_LC_13_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_c2_0_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_c2_0_LC_13_24_7 .LUT_INIT=16'b0100110111011101;
    LogicCell40 \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_c2_0_LC_13_24_7  (
            .in0(N__10534),
            .in1(N__10507),
            .in2(N__10478),
            .in3(N__11896),
            .lcout(\this_vga_signals.mult1_un68_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_25_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_25_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(N__11567),
            .in2(_gnd_net_),
            .in3(N__11693),
            .lcout(\this_vga_signals.N_469_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_RNI18AF_4_LC_14_16_3 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_RNI18AF_4_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \this_delay_clk.M_pipe_q_RNI18AF_4_LC_14_16_3 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \this_delay_clk.M_pipe_q_RNI18AF_4_LC_14_16_3  (
            .in0(N__12824),
            .in1(N__12841),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(debug_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.rgb_cnst_i_a5_0_0_3_LC_14_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.rgb_cnst_i_a5_0_0_3_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.rgb_cnst_i_a5_0_0_3_LC_14_16_7 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \this_vga_signals.rgb_cnst_i_a5_0_0_3_LC_14_16_7  (
            .in0(N__15816),
            .in1(N__18943),
            .in2(N__15879),
            .in3(N__18404),
            .lcout(\this_vga_signals.rgb_cnst_i_a5_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIETEJ4_2_11_LC_14_17_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIETEJ4_2_11_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIETEJ4_2_11_LC_14_17_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_radreg_RNIETEJ4_2_11_LC_14_17_7  (
            .in0(N__18944),
            .in1(N__18397),
            .in2(_gnd_net_),
            .in3(N__15800),
            .lcout(M_this_vram_read_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m3_5_LC_14_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m3_5_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m3_5_LC_14_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un16_address_if_m3_5_LC_14_18_0  (
            .in0(N__17180),
            .in1(N__10832),
            .in2(N__12398),
            .in3(N__11043),
            .lcout(),
            .ltout(\this_vga_signals.if_m3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m5_4_LC_14_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m5_4_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m5_4_LC_14_18_1 .LUT_INIT=16'b1010101000010111;
    LogicCell40 \this_vga_signals.un16_address_if_m5_4_LC_14_18_1  (
            .in0(N__12181),
            .in1(N__12473),
            .in2(N__10820),
            .in3(N__10817),
            .lcout(),
            .ltout(\this_vga_signals.if_m5_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIC40KO51_3_LC_14_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIC40KO51_3_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIC40KO51_3_LC_14_18_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIC40KO51_3_LC_14_18_2  (
            .in0(N__10793),
            .in1(N__11057),
            .in2(N__10811),
            .in3(N__12057),
            .lcout(\this_vga_signals.g1_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_o2_1_LC_14_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_o2_1_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_o2_1_LC_14_18_3 .LUT_INIT=16'b0001011100101011;
    LogicCell40 \this_vga_signals.un16_address_g0_i_o2_1_LC_14_18_3  (
            .in0(N__10980),
            .in1(N__12348),
            .in2(N__11458),
            .in3(N__10915),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_1_LC_14_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_1_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_1_LC_14_18_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_1_LC_14_18_5  (
            .in0(N__11422),
            .in1(N__10916),
            .in2(_gnd_net_),
            .in3(N__17178),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_axb2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_LC_14_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_LC_14_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_LC_14_18_6  (
            .in0(N__12347),
            .in1(N__11173),
            .in2(N__10796),
            .in3(N__10981),
            .lcout(\this_vga_signals.mult1_un68_sum_axb2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIRV8NA3_3_LC_14_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIRV8NA3_3_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIRV8NA3_3_LC_14_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIRV8NA3_3_LC_14_18_7  (
            .in0(N__11174),
            .in1(N__12349),
            .in2(_gnd_net_),
            .in3(N__17179),
            .lcout(\this_vga_signals.g1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_m2_5_0_LC_14_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_m2_5_0_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_m2_5_0_LC_14_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un16_address_if_m2_5_0_LC_14_19_0  (
            .in0(N__16086),
            .in1(N__10787),
            .in2(_gnd_net_),
            .in3(N__16140),
            .lcout(\this_vga_signals.if_m2_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_14_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_14_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_14_19_2  (
            .in0(N__12394),
            .in1(N__11044),
            .in2(_gnd_net_),
            .in3(N__17162),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_1_1_LC_14_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_1_1_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_1_1_LC_14_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un16_address_g0_1_1_LC_14_19_3  (
            .in0(N__17163),
            .in1(N__12351),
            .in2(_gnd_net_),
            .in3(N__11192),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_21_LC_14_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_21_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_21_LC_14_19_4 .LUT_INIT=16'b0100000000001000;
    LogicCell40 \this_vga_signals.un16_address_g0_21_LC_14_19_4  (
            .in0(N__16085),
            .in1(N__12172),
            .in2(N__11096),
            .in3(N__12058),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_ac0_3_d_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_17_LC_14_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_17_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_17_LC_14_19_5 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \this_vga_signals.un16_address_g0_17_LC_14_19_5  (
            .in0(N__11093),
            .in1(N__12578),
            .in2(N__11084),
            .in3(N__11081),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_o2_0_0_x2_0_LC_14_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_o2_0_0_x2_0_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_o2_0_0_x2_0_LC_14_19_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un16_address_g0_i_o2_0_0_x2_0_LC_14_19_6  (
            .in0(N__11191),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17161),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_o2_0_0_x2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_o2_0_0_o4_LC_14_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_o2_0_0_o4_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_o2_0_0_o4_LC_14_19_7 .LUT_INIT=16'b0100110111010100;
    LogicCell40 \this_vga_signals.un16_address_g0_i_o2_0_0_o4_LC_14_19_7  (
            .in0(N__12171),
            .in1(N__12352),
            .in2(N__11060),
            .in3(N__16084),
            .lcout(\this_vga_signals.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_i_3_LC_14_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_i_3_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_i_3_LC_14_20_2 .LUT_INIT=16'b1001001100110110;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_i_3_LC_14_20_2  (
            .in0(N__17187),
            .in1(N__11193),
            .in2(N__11051),
            .in3(N__11006),
            .lcout(rgb_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_c2_LC_14_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_c2_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_c2_LC_14_20_3 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_c2_LC_14_20_3  (
            .in0(N__11442),
            .in1(N__10987),
            .in2(N__12354),
            .in3(N__10912),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_o2_LC_14_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_o2_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_o2_LC_14_20_7 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un16_address_g0_i_o2_LC_14_20_7  (
            .in0(N__11443),
            .in1(N__10988),
            .in2(N__12355),
            .in3(N__10913),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_0_LC_14_21_7.C_ON=1'b0;
    defparam M_current_address_q_0_LC_14_21_7.SEQ_MODE=4'b1000;
    defparam M_current_address_q_0_LC_14_21_7.LUT_INIT=16'b1011100011100010;
    LogicCell40 M_current_address_q_0_LC_14_21_7 (
            .in0(N__12593),
            .in1(N__15576),
            .in2(N__11912),
            .in3(N__16327),
            .lcout(M_current_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18201),
            .ce(),
            .sr(N__15321));
    defparam M_current_address_q_RNO_0_0_LC_14_22_3.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_0_LC_14_22_3.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_0_LC_14_22_3.LUT_INIT=16'b1100110011100100;
    LogicCell40 M_current_address_q_RNO_0_0_LC_14_22_3 (
            .in0(N__16460),
            .in1(N__12627),
            .in2(N__17622),
            .in3(N__16326),
            .lcout(N_401),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKNO0B_9_LC_14_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKNO0B_9_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKNO0B_9_LC_14_23_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIKNO0B_9_LC_14_23_0  (
            .in0(N__20266),
            .in1(N__11902),
            .in2(_gnd_net_),
            .in3(N__11873),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_14_25_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_14_25_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_14_25_0 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(N__11707),
            .in2(N__11614),
            .in3(N__11735),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18214),
            .ce(),
            .sr(N__11578));
    defparam \this_vga_signals.M_hcounter_q_0_LC_14_25_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_14_25_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_14_25_1 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_14_25_1  (
            .in0(N__11708),
            .in1(N__11606),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18214),
            .ce(),
            .sr(N__11578));
    defparam \this_vga_signals.un16_address_g0_1_N_7L13_LC_15_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_1_N_7L13_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_1_N_7L13_LC_15_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un16_address_g0_1_N_7L13_LC_15_18_2  (
            .in0(N__12350),
            .in1(N__11194),
            .in2(_gnd_net_),
            .in3(N__17197),
            .lcout(\this_vga_signals.g0_1_N_7L13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.rgb_bm_1_LC_15_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.rgb_bm_1_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.rgb_bm_1_LC_15_18_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vga_signals.rgb_bm_1_LC_15_18_4  (
            .in0(N__14889),
            .in1(N__14006),
            .in2(_gnd_net_),
            .in3(N__13066),
            .lcout(\this_vga_signals.rgb_bmZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_15_18_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_15_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11531),
            .lcout(\this_delay_clk.M_this_delay_clk_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18189),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_23_LC_15_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_23_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_23_LC_15_18_6 .LUT_INIT=16'b1100001101101001;
    LogicCell40 \this_vga_signals.un16_address_g0_23_LC_15_18_6  (
            .in0(N__12563),
            .in1(N__11513),
            .in2(N__11459),
            .in3(N__12527),
            .lcout(),
            .ltout(\this_vga_signals.if_N_13_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_20_LC_15_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_20_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_20_LC_15_18_7 .LUT_INIT=16'b0000101011110101;
    LogicCell40 \this_vga_signals.un16_address_g0_20_LC_15_18_7  (
            .in0(N__17198),
            .in1(_gnd_net_),
            .in2(N__11198),
            .in3(N__11195),
            .lcout(\this_vga_signals.if_N_16_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_1_N_6L11_LC_15_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_1_N_6L11_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_1_N_6L11_LC_15_19_0 .LUT_INIT=16'b1010011001011001;
    LogicCell40 \this_vga_signals.un16_address_g0_1_N_6L11_LC_15_19_0  (
            .in0(N__12572),
            .in1(N__12562),
            .in2(N__12523),
            .in3(N__12485),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_N_6L11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_1_N_8L15_LC_15_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_1_N_8L15_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_1_N_8L15_LC_15_19_1 .LUT_INIT=16'b0010010001000010;
    LogicCell40 \this_vga_signals.un16_address_g0_1_N_8L15_LC_15_19_1  (
            .in0(N__12173),
            .in1(N__12474),
            .in2(N__12401),
            .in3(N__12390),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_N_8L15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_1_LC_15_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_1_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_1_LC_15_19_2 .LUT_INIT=16'b1010011010101001;
    LogicCell40 \this_vga_signals.un16_address_g0_1_LC_15_19_2  (
            .in0(N__12174),
            .in1(N__12374),
            .in2(N__12368),
            .in3(N__16087),
            .lcout(\this_vga_signals.if_N_6_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_vga_signals_address_a0_b_0_LC_15_19_3.C_ON=1'b0;
    defparam un1_M_this_vga_signals_address_a0_b_0_LC_15_19_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_vga_signals_address_a0_b_0_LC_15_19_3.LUT_INIT=16'b0110011000000000;
    LogicCell40 un1_M_this_vga_signals_address_a0_b_0_LC_15_19_3 (
            .in0(N__16142),
            .in1(N__16093),
            .in2(_gnd_net_),
            .in3(N__17879),
            .lcout(a0_b_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_i_o2_0_LC_15_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_i_o2_0_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_i_o2_0_LC_15_19_4 .LUT_INIT=16'b0010101110001110;
    LogicCell40 \this_vga_signals.un16_address_g0_i_o2_0_LC_15_19_4  (
            .in0(N__12353),
            .in1(N__16141),
            .in2(N__12182),
            .in3(N__16088),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un16_address_g0_0_LC_15_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un16_address_g0_0_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un16_address_g0_0_LC_15_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un16_address_g0_0_LC_15_19_5  (
            .in0(N__16089),
            .in1(N__12059),
            .in2(N__12032),
            .in3(N__12029),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI10UUE23_9_LC_15_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI10UUE23_9_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI10UUE23_9_LC_15_19_6 .LUT_INIT=16'b0100100010000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI10UUE23_9_LC_15_19_6  (
            .in0(N__20473),
            .in1(N__20298),
            .in2(N__12023),
            .in3(N__20449),
            .lcout(M_this_vga_signals_address_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_15_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_15_20_1 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_15_20_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_15_20_1  (
            .in0(N__12823),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12857),
            .lcout(this_start_data_delay_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18193),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIMM211_LC_15_20_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIMM211_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIMM211_LC_15_20_2 .LUT_INIT=16'b0110011001101110;
    LogicCell40 \this_start_data_delay.M_last_q_RNIMM211_LC_15_20_2  (
            .in0(N__15558),
            .in1(N__16301),
            .in2(N__12746),
            .in3(N__12800),
            .lcout(N_312_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_RNIBJQQ_4_LC_15_20_4 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_RNIBJQQ_4_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \this_delay_clk.M_pipe_q_RNIBJQQ_4_LC_15_20_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \this_delay_clk.M_pipe_q_RNIBJQQ_4_LC_15_20_4  (
            .in0(N__12744),
            .in1(N__12856),
            .in2(_gnd_net_),
            .in3(N__12822),
            .lcout(N_349_0),
            .ltout(N_349_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_8_LC_15_20_5.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_8_LC_15_20_5.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_8_LC_15_20_5.LUT_INIT=16'b1101111110000000;
    LogicCell40 M_current_address_q_RNO_0_8_LC_15_20_5 (
            .in0(N__16302),
            .in1(N__16636),
            .in2(N__12860),
            .in3(N__13870),
            .lcout(N_409),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_RNI18AF_0_4_LC_15_20_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_RNI18AF_0_4_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \this_delay_clk.M_pipe_q_RNI18AF_0_4_LC_15_20_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_delay_clk.M_pipe_q_RNI18AF_0_4_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__12855),
            .in2(_gnd_net_),
            .in3(N__12821),
            .lcout(debug_0),
            .ltout(debug_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_address_ibuf_RNIR5I81_7_LC_15_20_7.C_ON=1'b0;
    defparam port_address_ibuf_RNIR5I81_7_LC_15_20_7.SEQ_MODE=4'b0000;
    defparam port_address_ibuf_RNIR5I81_7_LC_15_20_7.LUT_INIT=16'b0001000000000000;
    LogicCell40 port_address_ibuf_RNIR5I81_7_LC_15_20_7 (
            .in0(N__12794),
            .in1(N__12770),
            .in2(N__12749),
            .in3(N__12745),
            .lcout(M_state_q_ns_0_a3_0_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_0_LC_15_21_0.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_0_LC_15_21_0.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_0_LC_15_21_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_0_LC_15_21_0 (
            .in0(_gnd_net_),
            .in1(N__12628),
            .in2(N__12608),
            .in3(N__12607),
            .lcout(M_current_address_q_RNO_1Z0Z_0),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(un1_M_current_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_1_LC_15_21_1.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_1_LC_15_21_1.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_1_LC_15_21_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_1_LC_15_21_1 (
            .in0(_gnd_net_),
            .in1(N__13135),
            .in2(_gnd_net_),
            .in3(N__12587),
            .lcout(M_current_address_q_RNO_1Z0Z_1),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_0),
            .carryout(un1_M_current_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_2_LC_15_21_2.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_2_LC_15_21_2.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_2_LC_15_21_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_2_LC_15_21_2 (
            .in0(_gnd_net_),
            .in1(N__15619),
            .in2(_gnd_net_),
            .in3(N__12584),
            .lcout(M_current_address_q_RNO_1Z0Z_2),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_1),
            .carryout(un1_M_current_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_3_LC_15_21_3.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_3_LC_15_21_3.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_3_LC_15_21_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_3_LC_15_21_3 (
            .in0(_gnd_net_),
            .in1(N__13407),
            .in2(_gnd_net_),
            .in3(N__12581),
            .lcout(M_current_address_q_RNO_1Z0Z_3),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_2),
            .carryout(un1_M_current_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_4_LC_15_21_4.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_4_LC_15_21_4.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_4_LC_15_21_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_4_LC_15_21_4 (
            .in0(_gnd_net_),
            .in1(N__14575),
            .in2(_gnd_net_),
            .in3(N__12887),
            .lcout(M_current_address_q_RNO_1Z0Z_4),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_3),
            .carryout(un1_M_current_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_5_LC_15_21_5.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_5_LC_15_21_5.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_5_LC_15_21_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_5_LC_15_21_5 (
            .in0(_gnd_net_),
            .in1(N__13270),
            .in2(_gnd_net_),
            .in3(N__12884),
            .lcout(M_current_address_q_RNO_1Z0Z_5),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_4),
            .carryout(un1_M_current_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_6_LC_15_21_6.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_6_LC_15_21_6.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_6_LC_15_21_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_6_LC_15_21_6 (
            .in0(_gnd_net_),
            .in1(N__15358),
            .in2(_gnd_net_),
            .in3(N__12881),
            .lcout(M_current_address_q_RNO_1Z0Z_6),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_5),
            .carryout(un1_M_current_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_7_LC_15_21_7.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_7_LC_15_21_7.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_7_LC_15_21_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_7_LC_15_21_7 (
            .in0(_gnd_net_),
            .in1(N__14716),
            .in2(_gnd_net_),
            .in3(N__12878),
            .lcout(M_current_address_q_RNO_1Z0Z_7),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_6),
            .carryout(un1_M_current_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_8_LC_15_22_0.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_8_LC_15_22_0.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_8_LC_15_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_8_LC_15_22_0 (
            .in0(_gnd_net_),
            .in1(N__13866),
            .in2(_gnd_net_),
            .in3(N__12875),
            .lcout(M_current_address_q_RNO_1Z0Z_8),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(un1_M_current_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_9_LC_15_22_1.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_9_LC_15_22_1.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_9_LC_15_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_9_LC_15_22_1 (
            .in0(_gnd_net_),
            .in1(N__15127),
            .in2(_gnd_net_),
            .in3(N__12872),
            .lcout(M_current_address_q_RNO_1Z0Z_9),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_8),
            .carryout(un1_M_current_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_10_LC_15_22_2.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_10_LC_15_22_2.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_10_LC_15_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_10_LC_15_22_2 (
            .in0(_gnd_net_),
            .in1(N__13543),
            .in2(_gnd_net_),
            .in3(N__12869),
            .lcout(M_current_address_q_RNO_1Z0Z_10),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_9),
            .carryout(un1_M_current_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_11_LC_15_22_3.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_11_LC_15_22_3.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_11_LC_15_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_11_LC_15_22_3 (
            .in0(_gnd_net_),
            .in1(N__19390),
            .in2(_gnd_net_),
            .in3(N__12866),
            .lcout(M_current_address_q_RNO_1Z0Z_11),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_10),
            .carryout(un1_M_current_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_12_LC_15_22_4.C_ON=1'b1;
    defparam M_current_address_q_RNO_1_12_LC_15_22_4.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_12_LC_15_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNO_1_12_LC_15_22_4 (
            .in0(_gnd_net_),
            .in1(N__19544),
            .in2(_gnd_net_),
            .in3(N__12863),
            .lcout(M_current_address_q_RNO_1Z0Z_12),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_11),
            .carryout(un1_M_current_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_1_13_LC_15_22_5.C_ON=1'b0;
    defparam M_current_address_q_RNO_1_13_LC_15_22_5.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_1_13_LC_15_22_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 M_current_address_q_RNO_1_13_LC_15_22_5 (
            .in0(_gnd_net_),
            .in1(N__19462),
            .in2(_gnd_net_),
            .in3(N__13043),
            .lcout(M_current_address_q_RNO_1Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clock.M_counter_q_0_LC_15_23_5 .C_ON=1'b0;
    defparam \this_pixel_clock.M_counter_q_0_LC_15_23_5 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clock.M_counter_q_0_LC_15_23_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_pixel_clock.M_counter_q_0_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__15308),
            .in2(_gnd_net_),
            .in3(N__13032),
            .lcout(\this_pixel_clock.M_counter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18204),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIMTEJ4_1_11_LC_16_16_3 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIMTEJ4_1_11_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIMTEJ4_1_11_LC_16_16_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_radreg_RNIMTEJ4_1_11_LC_16_16_3  (
            .in0(N__18974),
            .in1(N__18485),
            .in2(_gnd_net_),
            .in3(N__15836),
            .lcout(M_this_vram_read_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.rgb_bm_0_LC_16_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.rgb_bm_0_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.rgb_bm_0_LC_16_17_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vga_signals.rgb_bm_0_LC_16_17_0  (
            .in0(N__12896),
            .in1(N__14479),
            .in2(_gnd_net_),
            .in3(N__14904),
            .lcout(\this_vga_signals.rgb_bmZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.rgb_bm_2_LC_16_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.rgb_bm_2_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.rgb_bm_2_LC_16_17_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vga_signals.rgb_bm_2_LC_16_17_2  (
            .in0(N__14905),
            .in1(N__14480),
            .in2(_gnd_net_),
            .in3(N__13100),
            .lcout(\this_vga_signals.rgb_bmZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m7_am_LC_16_18_2.C_ON=1'b0;
    defparam rgb_2_5_0__m7_am_LC_16_18_2.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m7_am_LC_16_18_2.LUT_INIT=16'b0000010110101110;
    LogicCell40 rgb_2_5_0__m7_am_LC_16_18_2 (
            .in0(N__16768),
            .in1(N__16931),
            .in2(N__17006),
            .in3(N__16847),
            .lcout(),
            .ltout(m7_am_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m7_ns_LC_16_18_3.C_ON=1'b0;
    defparam rgb_2_5_0__m7_ns_LC_16_18_3.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m7_ns_LC_16_18_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 rgb_2_5_0__m7_ns_LC_16_18_3 (
            .in0(_gnd_net_),
            .in1(N__14948),
            .in2(N__12899),
            .in3(N__13112),
            .lcout(m7_ns),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m28_LC_16_18_5.C_ON=1'b0;
    defparam rgb_2_5_0__m28_LC_16_18_5.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m28_LC_16_18_5.LUT_INIT=16'b0001000100101000;
    LogicCell40 rgb_2_5_0__m28_LC_16_18_5 (
            .in0(N__16846),
            .in1(N__17002),
            .in2(N__16934),
            .in3(N__16767),
            .lcout(),
            .ltout(m28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m29_LC_16_18_6.C_ON=1'b0;
    defparam rgb_2_5_0__m29_LC_16_18_6.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m29_LC_16_18_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 rgb_2_5_0__m29_LC_16_18_6 (
            .in0(N__14947),
            .in1(_gnd_net_),
            .in2(N__12890),
            .in3(N__14513),
            .lcout(m29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m32_am_LC_16_19_3.C_ON=1'b0;
    defparam rgb_2_5_0__m32_am_LC_16_19_3.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m32_am_LC_16_19_3.LUT_INIT=16'b0010000101001000;
    LogicCell40 rgb_2_5_0__m32_am_LC_16_19_3 (
            .in0(N__16999),
            .in1(N__16843),
            .in2(N__16932),
            .in3(N__16762),
            .lcout(),
            .ltout(m32_am_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m32_ns_LC_16_19_4.C_ON=1'b0;
    defparam rgb_2_5_0__m32_ns_LC_16_19_4.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m32_ns_LC_16_19_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 rgb_2_5_0__m32_ns_LC_16_19_4 (
            .in0(N__14938),
            .in1(_gnd_net_),
            .in2(N__13115),
            .in3(N__13106),
            .lcout(m32_ns),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m7_bm_LC_16_19_5.C_ON=1'b0;
    defparam rgb_2_5_0__m7_bm_LC_16_19_5.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m7_bm_LC_16_19_5.LUT_INIT=16'b0000001011000000;
    LogicCell40 rgb_2_5_0__m7_bm_LC_16_19_5 (
            .in0(N__17001),
            .in1(N__16845),
            .in2(N__16933),
            .in3(N__16766),
            .lcout(m7_bm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m32_bm_LC_16_19_6.C_ON=1'b0;
    defparam rgb_2_5_0__m32_bm_LC_16_19_6.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m32_bm_LC_16_19_6.LUT_INIT=16'b0101001101010010;
    LogicCell40 rgb_2_5_0__m32_bm_LC_16_19_6 (
            .in0(N__16844),
            .in1(N__17000),
            .in2(N__16769),
            .in3(N__16924),
            .lcout(m32_bm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_11_LC_16_20_0.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_11_LC_16_20_0.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_11_LC_16_20_0.LUT_INIT=16'b1110101000101010;
    LogicCell40 M_current_address_q_RNO_0_11_LC_16_20_0 (
            .in0(N__19382),
            .in1(N__16436),
            .in2(N__16310),
            .in3(N__13828),
            .lcout(N_412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m42_LC_16_20_1.C_ON=1'b0;
    defparam rgb_2_5_0__m42_LC_16_20_1.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m42_LC_16_20_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 rgb_2_5_0__m42_LC_16_20_1 (
            .in0(N__14890),
            .in1(N__13099),
            .in2(_gnd_net_),
            .in3(N__14498),
            .lcout(rgb_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_5_LC_16_20_3.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_5_LC_16_20_3.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_5_LC_16_20_3.LUT_INIT=16'b1101100011001100;
    LogicCell40 M_current_address_q_RNO_0_5_LC_16_20_3 (
            .in0(N__16285),
            .in1(N__13269),
            .in2(N__13696),
            .in3(N__16450),
            .lcout(N_406),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_RNO_1_1_LC_16_20_4.C_ON=1'b0;
    defparam M_state_q_RNO_1_1_LC_16_20_4.SEQ_MODE=4'b0000;
    defparam M_state_q_RNO_1_1_LC_16_20_4.LUT_INIT=16'b0011001100000000;
    LogicCell40 M_state_q_RNO_1_1_LC_16_20_4 (
            .in0(_gnd_net_),
            .in1(N__16437),
            .in2(_gnd_net_),
            .in3(N__15529),
            .lcout(N_352),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.rgb_bm_3_LC_16_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.rgb_bm_3_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.rgb_bm_3_LC_16_20_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.rgb_bm_3_LC_16_20_5  (
            .in0(N__14447),
            .in1(N__14891),
            .in2(_gnd_net_),
            .in3(N__13070),
            .lcout(\this_vga_signals.rgb_bmZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_10_LC_16_20_6.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_10_LC_16_20_6.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_10_LC_16_20_6.LUT_INIT=16'b1110001010101010;
    LogicCell40 M_current_address_q_RNO_0_10_LC_16_20_6 (
            .in0(N__13542),
            .in1(N__16438),
            .in2(N__18050),
            .in3(N__16286),
            .lcout(N_411),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_3_LC_16_20_7.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_3_LC_16_20_7.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_3_LC_16_20_7.LUT_INIT=16'b1110010011110000;
    LogicCell40 M_current_address_q_RNO_0_3_LC_16_20_7 (
            .in0(N__16284),
            .in1(N__18049),
            .in2(N__13408),
            .in3(N__16449),
            .lcout(N_404),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_12_LC_16_21_1.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_12_LC_16_21_1.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_12_LC_16_21_1.LUT_INIT=16'b1110001010101010;
    LogicCell40 M_current_address_q_RNO_0_12_LC_16_21_1 (
            .in0(N__19545),
            .in1(N__16451),
            .in2(N__13697),
            .in3(N__16294),
            .lcout(),
            .ltout(N_413_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_12_LC_16_21_2.C_ON=1'b0;
    defparam M_current_address_q_12_LC_16_21_2.SEQ_MODE=4'b1000;
    defparam M_current_address_q_12_LC_16_21_2.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_12_LC_16_21_2 (
            .in0(N__16295),
            .in1(N__15575),
            .in2(N__13664),
            .in3(N__13661),
            .lcout(M_current_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18192),
            .ce(),
            .sr(N__15323));
    defparam M_current_address_q_10_LC_16_21_3.C_ON=1'b0;
    defparam M_current_address_q_10_LC_16_21_3.SEQ_MODE=4'b1000;
    defparam M_current_address_q_10_LC_16_21_3.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_10_LC_16_21_3 (
            .in0(N__15573),
            .in1(N__16296),
            .in2(N__13655),
            .in3(N__13646),
            .lcout(M_current_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18192),
            .ce(),
            .sr(N__15323));
    defparam M_current_address_q_3_LC_16_21_5.C_ON=1'b0;
    defparam M_current_address_q_3_LC_16_21_5.SEQ_MODE=4'b1000;
    defparam M_current_address_q_3_LC_16_21_5.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_3_LC_16_21_5 (
            .in0(N__15574),
            .in1(N__16297),
            .in2(N__13523),
            .in3(N__13514),
            .lcout(M_current_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18192),
            .ce(),
            .sr(N__15323));
    defparam M_current_address_q_5_LC_16_21_7.C_ON=1'b0;
    defparam M_current_address_q_5_LC_16_21_7.SEQ_MODE=4'b1000;
    defparam M_current_address_q_5_LC_16_21_7.LUT_INIT=16'b1011100011100010;
    LogicCell40 M_current_address_q_5_LC_16_21_7 (
            .in0(N__13382),
            .in1(N__15555),
            .in2(N__13376),
            .in3(N__16298),
            .lcout(M_current_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18192),
            .ce(),
            .sr(N__15323));
    defparam M_current_address_q_RNO_0_1_LC_16_22_0.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_1_LC_16_22_0.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_1_LC_16_22_0.LUT_INIT=16'b1100110011100100;
    LogicCell40 M_current_address_q_RNO_0_1_LC_16_22_0 (
            .in0(N__16462),
            .in1(N__13134),
            .in2(N__16635),
            .in3(N__16312),
            .lcout(),
            .ltout(N_402_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_1_LC_16_22_1.C_ON=1'b0;
    defparam M_current_address_q_1_LC_16_22_1.SEQ_MODE=4'b1000;
    defparam M_current_address_q_1_LC_16_22_1.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_1_LC_16_22_1 (
            .in0(N__15569),
            .in1(N__16328),
            .in2(N__13250),
            .in3(N__13247),
            .lcout(M_current_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18195),
            .ce(),
            .sr(N__15307));
    defparam M_current_address_q_8_LC_16_22_3.C_ON=1'b0;
    defparam M_current_address_q_8_LC_16_22_3.SEQ_MODE=4'b1000;
    defparam M_current_address_q_8_LC_16_22_3.LUT_INIT=16'b1101111010000100;
    LogicCell40 M_current_address_q_8_LC_16_22_3 (
            .in0(N__16314),
            .in1(N__13991),
            .in2(N__15578),
            .in3(N__13985),
            .lcout(M_current_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18195),
            .ce(),
            .sr(N__15307));
    defparam M_current_address_q_11_LC_16_22_5.C_ON=1'b0;
    defparam M_current_address_q_11_LC_16_22_5.SEQ_MODE=4'b1000;
    defparam M_current_address_q_11_LC_16_22_5.LUT_INIT=16'b1110110101001000;
    LogicCell40 M_current_address_q_11_LC_16_22_5 (
            .in0(N__16313),
            .in1(N__13844),
            .in2(N__15577),
            .in3(N__13835),
            .lcout(M_current_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18195),
            .ce(),
            .sr(N__15307));
    defparam M_current_address_q_RNO_0_4_LC_16_22_7.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_4_LC_16_22_7.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_4_LC_16_22_7.LUT_INIT=16'b1101100011001100;
    LogicCell40 M_current_address_q_RNO_0_4_LC_16_22_7 (
            .in0(N__16311),
            .in1(N__14568),
            .in2(N__13829),
            .in3(N__16461),
            .lcout(N_405),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_9_LC_16_23_7.C_ON=1'b0;
    defparam M_current_address_q_9_LC_16_23_7.SEQ_MODE=4'b1000;
    defparam M_current_address_q_9_LC_16_23_7.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_9_LC_16_23_7 (
            .in0(N__16321),
            .in1(N__15565),
            .in2(N__15107),
            .in3(N__13799),
            .lcout(M_current_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18200),
            .ce(),
            .sr(N__15312));
    defparam \this_vram.mem_radreg_RNIETEJ4_1_11_LC_17_14_3 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIETEJ4_1_11_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIETEJ4_1_11_LC_17_14_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \this_vram.mem_radreg_RNIETEJ4_1_11_LC_17_14_3  (
            .in0(N__15841),
            .in1(N__18737),
            .in2(N__18518),
            .in3(_gnd_net_),
            .lcout(M_this_vram_read_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_17_14_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_17_14_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_17_14_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_17_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb291_cry_0_c_LC_17_16_0.C_ON=1'b1;
    defparam rgb291_cry_0_c_LC_17_16_0.SEQ_MODE=4'b0000;
    defparam rgb291_cry_0_c_LC_17_16_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 rgb291_cry_0_c_LC_17_16_0 (
            .in0(_gnd_net_),
            .in1(N__14018),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(rgb291_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb291_cry_1_c_LC_17_16_1.C_ON=1'b1;
    defparam rgb291_cry_1_c_LC_17_16_1.SEQ_MODE=4'b0000;
    defparam rgb291_cry_1_c_LC_17_16_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 rgb291_cry_1_c_LC_17_16_1 (
            .in0(_gnd_net_),
            .in1(N__14150),
            .in2(N__14978),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(rgb291_cry_0),
            .carryout(rgb291_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb291_cry_2_c_LC_17_16_2.C_ON=1'b1;
    defparam rgb291_cry_2_c_LC_17_16_2.SEQ_MODE=4'b0000;
    defparam rgb291_cry_2_c_LC_17_16_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 rgb291_cry_2_c_LC_17_16_2 (
            .in0(_gnd_net_),
            .in1(N__15773),
            .in2(N__14182),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(rgb291_cry_1),
            .carryout(rgb291_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb291_cry_3_c_LC_17_16_3.C_ON=1'b1;
    defparam rgb291_cry_3_c_LC_17_16_3.SEQ_MODE=4'b0000;
    defparam rgb291_cry_3_c_LC_17_16_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 rgb291_cry_3_c_LC_17_16_3 (
            .in0(_gnd_net_),
            .in1(N__14024),
            .in2(N__14183),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(rgb291_cry_2),
            .carryout(rgb291),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI4ODS4_9_LC_17_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI4ODS4_9_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI4ODS4_9_LC_17_16_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI4ODS4_9_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__20329),
            .in2(_gnd_net_),
            .in3(N__14096),
            .lcout(\this_vga_signals.rgb_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_17_16_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_17_16_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_17_16_5  (
            .in0(N__15838),
            .in1(N__18973),
            .in2(_gnd_net_),
            .in3(N__18484),
            .lcout(mem_radreg_RNIMTEJ4_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIETEJ4_0_11_LC_17_16_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIETEJ4_0_11_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIETEJ4_0_11_LC_17_16_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_radreg_RNIETEJ4_0_11_LC_17_16_6  (
            .in0(N__18396),
            .in1(N__18936),
            .in2(_gnd_net_),
            .in3(N__15837),
            .lcout(mem_radreg_RNIETEJ4_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m44_LC_17_18_0.C_ON=1'b0;
    defparam rgb_2_5_0__m44_LC_17_18_0.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m44_LC_17_18_0.LUT_INIT=16'b0000110011010000;
    LogicCell40 rgb_2_5_0__m44_LC_17_18_0 (
            .in0(N__16908),
            .in1(N__16986),
            .in2(N__16842),
            .in3(N__16747),
            .lcout(),
            .ltout(m44_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m46_bm_LC_17_18_1.C_ON=1'b0;
    defparam rgb_2_5_0__m46_bm_LC_17_18_1.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m46_bm_LC_17_18_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 rgb_2_5_0__m46_bm_LC_17_18_1 (
            .in0(N__14512),
            .in1(_gnd_net_),
            .in2(N__14012),
            .in3(N__14951),
            .lcout(m46_bm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m22_am_LC_17_18_3.C_ON=1'b0;
    defparam rgb_2_5_0__m22_am_LC_17_18_3.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m22_am_LC_17_18_3.LUT_INIT=16'b0000101010110000;
    LogicCell40 rgb_2_5_0__m22_am_LC_17_18_3 (
            .in0(N__16984),
            .in1(N__16906),
            .in2(N__16760),
            .in3(N__16825),
            .lcout(),
            .ltout(m22_am_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m22_ns_LC_17_18_4.C_ON=1'b0;
    defparam rgb_2_5_0__m22_ns_LC_17_18_4.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m22_ns_LC_17_18_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 rgb_2_5_0__m22_ns_LC_17_18_4 (
            .in0(N__13997),
            .in1(_gnd_net_),
            .in2(N__14009),
            .in3(N__14937),
            .lcout(m22_ns),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m22_bm_LC_17_18_5.C_ON=1'b0;
    defparam rgb_2_5_0__m22_bm_LC_17_18_5.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m22_bm_LC_17_18_5.LUT_INIT=16'b0000111110101100;
    LogicCell40 rgb_2_5_0__m22_bm_LC_17_18_5 (
            .in0(N__16985),
            .in1(N__16907),
            .in2(N__16761),
            .in3(N__16826),
            .lcout(m22_bm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m24_LC_17_19_0.C_ON=1'b0;
    defparam rgb_2_5_0__m24_LC_17_19_0.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m24_LC_17_19_0.LUT_INIT=16'b0101100001001000;
    LogicCell40 rgb_2_5_0__m24_LC_17_19_0 (
            .in0(N__16809),
            .in1(N__16970),
            .in2(N__16740),
            .in3(N__16887),
            .lcout(m24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m40_LC_17_19_1.C_ON=1'b0;
    defparam rgb_2_5_0__m40_LC_17_19_1.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m40_LC_17_19_1.LUT_INIT=16'b0011000010101001;
    LogicCell40 rgb_2_5_0__m40_LC_17_19_1 (
            .in0(N__16971),
            .in1(N__16810),
            .in2(N__16905),
            .in3(N__16727),
            .lcout(),
            .ltout(m40_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m41_LC_17_19_2.C_ON=1'b0;
    defparam rgb_2_5_0__m41_LC_17_19_2.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m41_LC_17_19_2.LUT_INIT=16'b1010101011110000;
    LogicCell40 rgb_2_5_0__m41_LC_17_19_2 (
            .in0(N__14492),
            .in1(_gnd_net_),
            .in2(N__14501),
            .in3(N__14936),
            .lcout(m41),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m10_LC_17_19_3.C_ON=1'b0;
    defparam rgb_2_5_0__m10_LC_17_19_3.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m10_LC_17_19_3.LUT_INIT=16'b0000000010111100;
    LogicCell40 rgb_2_5_0__m10_LC_17_19_3 (
            .in0(N__16968),
            .in1(N__16807),
            .in2(N__16903),
            .in3(N__16722),
            .lcout(m10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1UGICK_9_LC_17_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1UGICK_9_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1UGICK_9_LC_17_19_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI1UGICK_9_LC_17_19_4  (
            .in0(N__14465),
            .in1(N__17873),
            .in2(_gnd_net_),
            .in3(N__17169),
            .lcout(rgb_1_axb_0),
            .ltout(rgb_1_axb_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m15_LC_17_19_5.C_ON=1'b0;
    defparam rgb_2_5_0__m15_LC_17_19_5.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m15_LC_17_19_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 rgb_2_5_0__m15_LC_17_19_5 (
            .in0(_gnd_net_),
            .in1(N__14491),
            .in2(N__14483),
            .in3(N__15767),
            .lcout(m15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m19_LC_17_19_7.C_ON=1'b0;
    defparam rgb_2_5_0__m19_LC_17_19_7.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m19_LC_17_19_7.LUT_INIT=16'b0010001110001000;
    LogicCell40 rgb_2_5_0__m19_LC_17_19_7 (
            .in0(N__16969),
            .in1(N__16808),
            .in2(N__16904),
            .in3(N__16723),
            .lcout(m19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_1_cry_0_0_c_RNO_LC_17_20_1.C_ON=1'b0;
    defparam rgb_1_cry_0_0_c_RNO_LC_17_20_1.SEQ_MODE=4'b0000;
    defparam rgb_1_cry_0_0_c_RNO_LC_17_20_1.LUT_INIT=16'b1001101011000000;
    LogicCell40 rgb_1_cry_0_0_c_RNO_LC_17_20_1 (
            .in0(N__17869),
            .in1(N__14461),
            .in2(N__17878),
            .in3(N__17199),
            .lcout(rgb_1_cry_0_0_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m37_LC_17_20_2.C_ON=1'b0;
    defparam rgb_2_5_0__m37_LC_17_20_2.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m37_LC_17_20_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 rgb_2_5_0__m37_LC_17_20_2 (
            .in0(N__14949),
            .in1(N__14962),
            .in2(_gnd_net_),
            .in3(N__16687),
            .lcout(m37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m46_am_LC_17_20_3.C_ON=1'b0;
    defparam rgb_2_5_0__m46_am_LC_17_20_3.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m46_am_LC_17_20_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 rgb_2_5_0__m46_am_LC_17_20_3 (
            .in0(N__16688),
            .in1(N__14963),
            .in2(_gnd_net_),
            .in3(N__14950),
            .lcout(),
            .ltout(m46_am_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m46_ns_LC_17_20_4.C_ON=1'b0;
    defparam rgb_2_5_0__m46_ns_LC_17_20_4.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m46_ns_LC_17_20_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 rgb_2_5_0__m46_ns_LC_17_20_4 (
            .in0(_gnd_net_),
            .in1(N__14906),
            .in2(N__14861),
            .in3(N__14858),
            .lcout(rgb_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_1_LC_17_20_5.C_ON=1'b0;
    defparam M_state_q_1_LC_17_20_5.SEQ_MODE=4'b1000;
    defparam M_state_q_1_LC_17_20_5.LUT_INIT=16'b0101010001000100;
    LogicCell40 M_state_q_1_LC_17_20_5 (
            .in0(N__15325),
            .in1(N__14834),
            .in2(N__14549),
            .in3(N__16643),
            .lcout(M_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18194),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_0_LC_17_20_6.C_ON=1'b0;
    defparam M_state_q_0_LC_17_20_6.SEQ_MODE=4'b1000;
    defparam M_state_q_0_LC_17_20_6.LUT_INIT=16'b0011000000110010;
    LogicCell40 M_state_q_0_LC_17_20_6 (
            .in0(N__16241),
            .in1(N__15326),
            .in2(N__14522),
            .in3(N__16453),
            .lcout(M_state_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18194),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_RNIMM211_1_LC_17_20_7.C_ON=1'b0;
    defparam M_state_q_RNIMM211_1_LC_17_20_7.SEQ_MODE=4'b0000;
    defparam M_state_q_RNIMM211_1_LC_17_20_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 M_state_q_RNIMM211_1_LC_17_20_7 (
            .in0(N__16452),
            .in1(N__15522),
            .in2(_gnd_net_),
            .in3(N__16240),
            .lcout(M_this_vram_write_en_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_7_LC_17_21_0.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_7_LC_17_21_0.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_7_LC_17_21_0.LUT_INIT=16'b1110101000101010;
    LogicCell40 M_current_address_q_RNO_0_7_LC_17_21_0 (
            .in0(N__14712),
            .in1(N__16473),
            .in2(N__16325),
            .in3(N__17623),
            .lcout(),
            .ltout(N_408_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_7_LC_17_21_1.C_ON=1'b0;
    defparam M_current_address_q_7_LC_17_21_1.SEQ_MODE=4'b1000;
    defparam M_current_address_q_7_LC_17_21_1.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_7_LC_17_21_1 (
            .in0(N__16299),
            .in1(N__15557),
            .in2(N__14828),
            .in3(N__14825),
            .lcout(M_current_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18197),
            .ce(),
            .sr(N__15324));
    defparam M_current_address_q_4_LC_17_21_2.C_ON=1'b0;
    defparam M_current_address_q_4_LC_17_21_2.SEQ_MODE=4'b1000;
    defparam M_current_address_q_4_LC_17_21_2.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_4_LC_17_21_2 (
            .in0(N__15556),
            .in1(N__16300),
            .in2(N__14693),
            .in3(N__14684),
            .lcout(M_current_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18197),
            .ce(),
            .sr(N__15324));
    defparam M_state_q_RNO_0_0_LC_17_21_6.C_ON=1'b0;
    defparam M_state_q_RNO_0_0_LC_17_21_6.SEQ_MODE=4'b0000;
    defparam M_state_q_RNO_0_0_LC_17_21_6.LUT_INIT=16'b0000000001000000;
    LogicCell40 M_state_q_RNO_0_0_LC_17_21_6 (
            .in0(N__16678),
            .in1(N__14545),
            .in2(N__19964),
            .in3(N__15530),
            .lcout(N_351),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_2_LC_17_22_1.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_2_LC_17_22_1.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_2_LC_17_22_1.LUT_INIT=16'b1011101010001010;
    LogicCell40 M_current_address_q_RNO_0_2_LC_17_22_1 (
            .in0(N__15606),
            .in1(N__16317),
            .in2(N__16478),
            .in3(N__19771),
            .lcout(),
            .ltout(N_403_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_2_LC_17_22_2.C_ON=1'b0;
    defparam M_current_address_q_2_LC_17_22_2.SEQ_MODE=4'b1000;
    defparam M_current_address_q_2_LC_17_22_2.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_2_LC_17_22_2 (
            .in0(N__16318),
            .in1(N__15564),
            .in2(N__15725),
            .in3(N__15722),
            .lcout(M_current_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18202),
            .ce(),
            .sr(N__15322));
    defparam M_current_address_q_13_LC_17_22_3.C_ON=1'b0;
    defparam M_current_address_q_13_LC_17_22_3.SEQ_MODE=4'b1000;
    defparam M_current_address_q_13_LC_17_22_3.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_13_LC_17_22_3 (
            .in0(N__15562),
            .in1(N__16319),
            .in2(N__16160),
            .in3(N__15587),
            .lcout(M_current_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18202),
            .ce(),
            .sr(N__15322));
    defparam M_current_address_q_RNO_0_6_LC_17_22_4.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_6_LC_17_22_4.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_6_LC_17_22_4.LUT_INIT=16'b1101100011001100;
    LogicCell40 M_current_address_q_RNO_0_6_LC_17_22_4 (
            .in0(N__16316),
            .in1(N__15345),
            .in2(N__16376),
            .in3(N__16477),
            .lcout(),
            .ltout(N_407_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_6_LC_17_22_5.C_ON=1'b0;
    defparam M_current_address_q_6_LC_17_22_5.SEQ_MODE=4'b1000;
    defparam M_current_address_q_6_LC_17_22_5.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_6_LC_17_22_5 (
            .in0(N__15563),
            .in1(N__16320),
            .in2(N__15473),
            .in3(N__15470),
            .lcout(M_current_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18202),
            .ce(),
            .sr(N__15322));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICJRF0D_9_LC_17_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICJRF0D_9_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICJRF0D_9_LC_17_23_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICJRF0D_9_LC_17_23_1  (
            .in0(N__17874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17201),
            .lcout(M_vcounter_q_esr_RNICJRF0D_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_9_LC_17_23_3.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_9_LC_17_23_3.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_9_LC_17_23_3.LUT_INIT=16'b1110001010101010;
    LogicCell40 M_current_address_q_RNO_0_9_LC_17_23_3 (
            .in0(N__15126),
            .in1(N__16472),
            .in2(N__19772),
            .in3(N__16315),
            .lcout(N_410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRM6F7_9_LC_17_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRM6F7_9_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRM6F7_9_LC_17_23_6 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIRM6F7_9_LC_17_23_6  (
            .in0(N__20262),
            .in1(N__15098),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIETEJ4_11_LC_18_14_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIETEJ4_11_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIETEJ4_11_LC_18_14_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_radreg_RNIETEJ4_11_LC_18_14_7  (
            .in0(N__18514),
            .in1(N__18736),
            .in2(_gnd_net_),
            .in3(N__15842),
            .lcout(mem_radreg_RNIETEJ4_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIMTEJ4_2_11_LC_18_16_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIMTEJ4_2_11_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIMTEJ4_2_11_LC_18_16_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_radreg_RNIMTEJ4_2_11_LC_18_16_0  (
            .in0(N__15840),
            .in1(N__19067),
            .in2(_gnd_net_),
            .in3(N__18821),
            .lcout(M_this_vram_read_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIMTEJ4_11_LC_18_16_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIMTEJ4_11_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIMTEJ4_11_LC_18_16_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_radreg_RNIMTEJ4_11_LC_18_16_5  (
            .in0(N__18820),
            .in1(N__19066),
            .in2(_gnd_net_),
            .in3(N__15839),
            .lcout(mem_radreg_RNIMTEJ4_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIB9J4TN_9_LC_18_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIB9J4TN_9_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIB9J4TN_9_LC_18_19_0 .LUT_INIT=16'b1011100001001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIB9J4TN_9_LC_18_19_0  (
            .in0(N__17846),
            .in1(N__17170),
            .in2(N__17865),
            .in3(N__17351),
            .lcout(M_vcounter_q_esr_RNIB9J4TN_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m14_LC_18_19_6.C_ON=1'b0;
    defparam rgb_2_5_0__m14_LC_18_19_6.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m14_LC_18_19_6.LUT_INIT=16'b0000100100110100;
    LogicCell40 rgb_2_5_0__m14_LC_18_19_6 (
            .in0(N__16880),
            .in1(N__16967),
            .in2(N__16824),
            .in3(N__16721),
            .lcout(m14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_1_cry_0_0_c_LC_18_20_0.C_ON=1'b1;
    defparam rgb_1_cry_0_0_c_LC_18_20_0.SEQ_MODE=4'b0000;
    defparam rgb_1_cry_0_0_c_LC_18_20_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 rgb_1_cry_0_0_c_LC_18_20_0 (
            .in0(_gnd_net_),
            .in1(N__15761),
            .in2(N__17021),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(rgb_1_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_1_cry_0_0_c_RNIFFTTT41_LC_18_20_1.C_ON=1'b1;
    defparam rgb_1_cry_0_0_c_RNIFFTTT41_LC_18_20_1.SEQ_MODE=4'b0000;
    defparam rgb_1_cry_0_0_c_RNIFFTTT41_LC_18_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rgb_1_cry_0_0_c_RNIFFTTT41_LC_18_20_1 (
            .in0(_gnd_net_),
            .in1(N__15755),
            .in2(N__15749),
            .in3(N__15737),
            .lcout(rgb_1_3),
            .ltout(),
            .carryin(rgb_1_cry_0),
            .carryout(rgb_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_1_cry_1_0_c_RNIPTLTE01_LC_18_20_2.C_ON=1'b1;
    defparam rgb_1_cry_1_0_c_RNIPTLTE01_LC_18_20_2.SEQ_MODE=4'b0000;
    defparam rgb_1_cry_1_0_c_RNIPTLTE01_LC_18_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rgb_1_cry_1_0_c_RNIPTLTE01_LC_18_20_2 (
            .in0(_gnd_net_),
            .in1(N__17012),
            .in2(N__17795),
            .in3(N__15734),
            .lcout(rgb_1_4),
            .ltout(),
            .carryin(rgb_1_cry_1),
            .carryout(rgb_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_1_cry_2_0_c_RNISLC8LA_LC_18_20_3.C_ON=1'b1;
    defparam rgb_1_cry_2_0_c_RNISLC8LA_LC_18_20_3.SEQ_MODE=4'b0000;
    defparam rgb_1_cry_2_0_c_RNISLC8LA_LC_18_20_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 rgb_1_cry_2_0_c_RNISLC8LA_LC_18_20_3 (
            .in0(_gnd_net_),
            .in1(N__17885),
            .in2(_gnd_net_),
            .in3(N__15731),
            .lcout(rgb_1_5),
            .ltout(),
            .carryin(rgb_1_cry_2),
            .carryout(rgb_1_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_1_6_THRU_LUT4_0_LC_18_20_4.C_ON=1'b0;
    defparam rgb_1_6_THRU_LUT4_0_LC_18_20_4.SEQ_MODE=4'b0000;
    defparam rgb_1_6_THRU_LUT4_0_LC_18_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 rgb_1_6_THRU_LUT4_0_LC_18_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15728),
            .lcout(rgb_1_6_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_1_cry_0_0_c_RNO_0_LC_18_20_5.C_ON=1'b0;
    defparam rgb_1_cry_0_0_c_RNO_0_LC_18_20_5.SEQ_MODE=4'b0000;
    defparam rgb_1_cry_0_0_c_RNO_0_LC_18_20_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 rgb_1_cry_0_0_c_RNO_0_LC_18_20_5 (
            .in0(_gnd_net_),
            .in1(N__17832),
            .in2(_gnd_net_),
            .in3(N__17200),
            .lcout(rgb_1_cry_0_0_c_RNOZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1H9RHL_9_LC_18_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1H9RHL_9_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1H9RHL_9_LC_18_20_6 .LUT_INIT=16'b1001101011000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI1H9RHL_9_LC_18_20_6  (
            .in0(N__17833),
            .in1(N__18363),
            .in2(N__17853),
            .in3(N__17350),
            .lcout(M_vcounter_q_esr_RNI1H9RHL_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_2_5_0__m36_LC_18_20_7.C_ON=1'b0;
    defparam rgb_2_5_0__m36_LC_18_20_7.SEQ_MODE=4'b0000;
    defparam rgb_2_5_0__m36_LC_18_20_7.LUT_INIT=16'b0000110101111110;
    LogicCell40 rgb_2_5_0__m36_LC_18_20_7 (
            .in0(N__16966),
            .in1(N__16879),
            .in2(N__16823),
            .in3(N__16720),
            .lcout(m36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_RNO_0_1_LC_18_21_0.C_ON=1'b0;
    defparam M_state_q_RNO_0_1_LC_18_21_0.SEQ_MODE=4'b0000;
    defparam M_state_q_RNO_0_1_LC_18_21_0.LUT_INIT=16'b0000000001100000;
    LogicCell40 M_state_q_RNO_0_1_LC_18_21_0 (
            .in0(N__16679),
            .in1(N__16655),
            .in2(N__19963),
            .in3(N__16287),
            .lcout(M_state_q_ns_0_a3_0_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_ibuf_RNI2PEE1_1_LC_18_21_5.C_ON=1'b0;
    defparam port_data_ibuf_RNI2PEE1_1_LC_18_21_5.SEQ_MODE=4'b0000;
    defparam port_data_ibuf_RNI2PEE1_1_LC_18_21_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 port_data_ibuf_RNI2PEE1_1_LC_18_21_5 (
            .in0(_gnd_net_),
            .in1(N__16637),
            .in2(_gnd_net_),
            .in3(N__19251),
            .lcout(M_this_vram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNO_0_13_LC_18_22_0.C_ON=1'b0;
    defparam M_current_address_q_RNO_0_13_LC_18_22_0.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNO_0_13_LC_18_22_0.LUT_INIT=16'b1110001010101010;
    LogicCell40 M_current_address_q_RNO_0_13_LC_18_22_0 (
            .in0(N__19432),
            .in1(N__16471),
            .in2(N__16375),
            .in3(N__16309),
            .lcout(N_414),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRN34U9_9_LC_19_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRN34U9_9_LC_19_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRN34U9_9_LC_19_19_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIRN34U9_9_LC_19_19_7  (
            .in0(N__20325),
            .in1(N__16148),
            .in2(_gnd_net_),
            .in3(N__16094),
            .lcout(M_this_vga_signals_address_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIRB7JA_9_LC_19_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIRB7JA_9_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIRB7JA_9_LC_19_20_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIRB7JA_9_LC_19_20_3  (
            .in0(N__17647),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15919),
            .lcout(rgbZ0Z_1),
            .ltout(rgbZ0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI2RH6LA_9_LC_19_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI2RH6LA_9_LC_19_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI2RH6LA_9_LC_19_20_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI2RH6LA_9_LC_19_20_4  (
            .in0(N__18370),
            .in1(_gnd_net_),
            .in2(N__17888),
            .in3(_gnd_net_),
            .lcout(M_vcounter_q_esr_RNI2RH6LA_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVLNKSA_9_LC_19_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVLNKSA_9_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIVLNKSA_9_LC_19_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIVLNKSA_9_LC_19_20_5  (
            .in0(N__17831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17339),
            .lcout(M_vcounter_q_esr_RNIVLNKSA_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIN383L_9_LC_19_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIN383L_9_LC_19_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIN383L_9_LC_19_23_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIN383L_9_LC_19_23_1  (
            .in0(_gnd_net_),
            .in1(N__20308),
            .in2(_gnd_net_),
            .in3(N__17783),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_ibuf_RNI1OEE1_0_LC_20_22_2.C_ON=1'b0;
    defparam port_data_ibuf_RNI1OEE1_0_LC_20_22_2.SEQ_MODE=4'b0000;
    defparam port_data_ibuf_RNI1OEE1_0_LC_20_22_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 port_data_ibuf_RNI1OEE1_0_LC_20_22_2 (
            .in0(_gnd_net_),
            .in1(N__17627),
            .in2(_gnd_net_),
            .in3(N__19297),
            .lcout(M_this_vram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIFAVQ5_9_LC_20_25_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIFAVQ5_9_LC_20_25_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIFAVQ5_9_LC_20_25_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIFAVQ5_9_LC_20_25_1  (
            .in0(_gnd_net_),
            .in1(N__20310),
            .in2(_gnd_net_),
            .in3(N__17498),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_21_15_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_21_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_21_15_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vram.mem_mem_1_0_wclke_3_LC_21_15_5  (
            .in0(N__19595),
            .in1(N__19391),
            .in2(N__19499),
            .in3(N__19309),
            .lcout(\this_vram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_12_LC_21_18_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_12_LC_21_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_12_LC_21_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vram.mem_radreg_12_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(N__20338),
            .in2(_gnd_net_),
            .in3(N__17349),
            .lcout(\this_vram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18203),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_22_15_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_22_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_22_15_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vram.mem_mem_3_0_wclke_3_LC_22_15_1  (
            .in0(N__19579),
            .in1(N__19394),
            .in2(N__19500),
            .in3(N__19310),
            .lcout(\this_vram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNISOI11_0_LC_23_12_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNISOI11_0_LC_23_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNISOI11_0_LC_23_12_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_0_1_RNISOI11_0_LC_23_12_1  (
            .in0(N__17219),
            .in1(N__19871),
            .in2(_gnd_net_),
            .in3(N__18533),
            .lcout(\this_vram.mem_mem_0_1_RNISOI11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_13_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_13_0  (
            .in0(N__18877),
            .in1(N__18680),
            .in2(_gnd_net_),
            .in3(N__18653),
            .lcout(\this_vram.mem_N_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5GH72_12_LC_23_14_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5GH72_12_LC_23_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5GH72_12_LC_23_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_radreg_RNI5GH72_12_LC_23_14_4  (
            .in0(N__18593),
            .in1(N__18494),
            .in2(_gnd_net_),
            .in3(N__18866),
            .lcout(\this_vram.mem_N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_23_15_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_23_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_23_15_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_vram.mem_mem_2_0_wclke_3_LC_23_15_3  (
            .in0(N__19312),
            .in1(N__19496),
            .in2(N__19601),
            .in3(N__19393),
            .lcout(\this_vram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_23_15_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_23_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_23_15_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vram.mem_mem_0_0_wclke_3_LC_23_15_6  (
            .in0(N__19596),
            .in1(N__19392),
            .in2(N__19502),
            .in3(N__19311),
            .lcout(\this_vram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI1GH72_12_LC_23_17_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI1GH72_12_LC_23_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI1GH72_12_LC_23_17_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_radreg_RNI1GH72_12_LC_23_17_2  (
            .in0(N__18851),
            .in1(N__19799),
            .in2(_gnd_net_),
            .in3(N__19937),
            .lcout(this_vram_mem_N_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_13_LC_23_17_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_13_LC_23_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_13_LC_23_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vram.mem_radreg_13_LC_23_17_7  (
            .in0(_gnd_net_),
            .in1(N__20339),
            .in2(_gnd_net_),
            .in3(N__18371),
            .lcout(\this_vram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18205),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_ibuf_RNI4REE1_3_LC_23_20_2.C_ON=1'b0;
    defparam port_data_ibuf_RNI4REE1_3_LC_23_20_2.SEQ_MODE=4'b0000;
    defparam port_data_ibuf_RNI4REE1_3_LC_23_20_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 port_data_ibuf_RNI4REE1_3_LC_23_20_2 (
            .in0(_gnd_net_),
            .in1(N__18045),
            .in2(_gnd_net_),
            .in3(N__19276),
            .lcout(M_this_vram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_12_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_12_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_12_3  (
            .in0(N__17915),
            .in1(N__17903),
            .in2(_gnd_net_),
            .in3(N__19878),
            .lcout(\this_vram.mem_mem_0_0_RNIQOI11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_12_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_12_6  (
            .in0(N__19879),
            .in1(N__18776),
            .in2(_gnd_net_),
            .in3(N__18764),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_0_RNIU0N11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_12_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_12_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_12_7  (
            .in0(N__18746),
            .in1(_gnd_net_),
            .in2(N__18740),
            .in3(N__18878),
            .lcout(\this_vram.mem_N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_13_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_13_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_13_1  (
            .in0(N__18707),
            .in1(N__19872),
            .in2(_gnd_net_),
            .in3(N__18695),
            .lcout(\this_vram.mem_mem_1_0_RNISSK11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_3  (
            .in0(N__18674),
            .in1(N__19877),
            .in2(_gnd_net_),
            .in3(N__18668),
            .lcout(\this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_13_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_13_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \this_vram.mem_mem_1_0_RNISSK11_LC_24_13_4  (
            .in0(N__18647),
            .in1(_gnd_net_),
            .in2(N__19880),
            .in3(N__18635),
            .lcout(\this_vram.mem_mem_1_0_RNISSKZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_13_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_13_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_13_5  (
            .in0(N__18620),
            .in1(N__19876),
            .in2(_gnd_net_),
            .in3(N__18611),
            .lcout(\this_vram.mem_mem_2_1_RNI01N11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_14_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_14_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_0_1_RNISOI11_LC_24_14_1  (
            .in0(N__18587),
            .in1(N__19868),
            .in2(_gnd_net_),
            .in3(N__18572),
            .lcout(\this_vram.mem_mem_0_1_RNISOIZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_14_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_14_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_1_1_RNIUSK11_LC_24_14_2  (
            .in0(N__19869),
            .in1(N__18560),
            .in2(_gnd_net_),
            .in3(N__18548),
            .lcout(\this_vram.mem_mem_1_1_RNIUSKZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_14_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_2_1_RNI01N11_LC_24_14_5  (
            .in0(N__19103),
            .in1(N__19094),
            .in2(_gnd_net_),
            .in3(N__19870),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_14_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_14_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_14_6  (
            .in0(N__18876),
            .in1(_gnd_net_),
            .in2(N__19076),
            .in3(N__19073),
            .lcout(\this_vram.mem_N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_15_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_15_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_15_0  (
            .in0(N__19046),
            .in1(N__19031),
            .in2(_gnd_net_),
            .in3(N__19841),
            .lcout(\this_vram.mem_mem_1_1_RNIUSK11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_1  (
            .in0(N__19842),
            .in1(_gnd_net_),
            .in2(N__19016),
            .in3(N__19007),
            .lcout(),
            .ltout(\this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI9OL72_12_LC_24_15_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI9OL72_12_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI9OL72_12_LC_24_15_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vram.mem_radreg_RNI9OL72_12_LC_24_15_2  (
            .in0(N__18865),
            .in1(_gnd_net_),
            .in2(N__18986),
            .in3(N__18983),
            .lcout(\this_vram.mem_N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5OL72_12_LC_24_15_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5OL72_12_LC_24_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5OL72_12_LC_24_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_radreg_RNI5OL72_12_LC_24_15_5  (
            .in0(N__18953),
            .in1(N__19907),
            .in2(_gnd_net_),
            .in3(N__18863),
            .lcout(this_vram_mem_N_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6  (
            .in0(N__18911),
            .in1(N__18905),
            .in2(_gnd_net_),
            .in3(N__19843),
            .lcout(),
            .ltout(\this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_15_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_15_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_15_7  (
            .in0(N__18887),
            .in1(_gnd_net_),
            .in2(N__18881),
            .in3(N__18864),
            .lcout(\this_vram.mem_N_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_16_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_16_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_2_0_RNIU0N11_LC_24_16_3  (
            .in0(N__19822),
            .in1(N__18803),
            .in2(_gnd_net_),
            .in3(N__18788),
            .lcout(\this_vram.mem_mem_2_0_RNIU0NZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_16_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_16_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_3_0_RNI05P11_LC_24_16_6  (
            .in0(N__19931),
            .in1(N__19823),
            .in2(_gnd_net_),
            .in3(N__19916),
            .lcout(\this_vram.mem_mem_3_0_RNI05PZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_3  (
            .in0(N__19901),
            .in1(N__19886),
            .in2(_gnd_net_),
            .in3(N__19821),
            .lcout(\this_vram.mem_mem_0_0_RNIQOIZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_24_18_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_24_18_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vram.mem_mem_4_0_wclke_3_LC_24_18_7  (
            .in0(N__19597),
            .in1(N__19402),
            .in2(N__19501),
            .in3(N__19316),
            .lcout(\this_vram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_ibuf_RNI3QEE1_2_LC_24_20_3.C_ON=1'b0;
    defparam port_data_ibuf_RNI3QEE1_2_LC_24_20_3.SEQ_MODE=4'b0000;
    defparam port_data_ibuf_RNI3QEE1_2_LC_24_20_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 port_data_ibuf_RNI3QEE1_2_LC_24_20_3 (
            .in0(_gnd_net_),
            .in1(N__19767),
            .in2(_gnd_net_),
            .in3(N__19277),
            .lcout(M_this_vram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_21_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_21_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vram.mem_mem_5_0_wclke_3_LC_24_21_5  (
            .in0(N__19580),
            .in1(N__19403),
            .in2(N__19498),
            .in3(N__19313),
            .lcout(\this_vram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_22_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_22_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vram.mem_mem_7_0_wclke_3_LC_24_22_4  (
            .in0(N__19315),
            .in1(N__19581),
            .in2(N__19497),
            .in3(N__19386),
            .lcout(\this_vram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_24_22_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_24_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_24_22_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vram.mem_mem_6_0_wclke_3_LC_24_22_7  (
            .in0(N__19582),
            .in1(N__19480),
            .in2(N__19401),
            .in3(N__19314),
            .lcout(\this_vram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI51C6S_9_LC_24_29_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI51C6S_9_LC_24_29_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI51C6S_9_LC_24_29_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI51C6S_9_LC_24_29_4  (
            .in0(_gnd_net_),
            .in1(N__20332),
            .in2(_gnd_net_),
            .in3(N__20167),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNID2F8IP1_9_LC_24_31_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNID2F8IP1_9_LC_24_31_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNID2F8IP1_9_LC_24_31_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNID2F8IP1_9_LC_24_31_4  (
            .in0(N__20333),
            .in1(N__20480),
            .in2(_gnd_net_),
            .in3(N__20459),
            .lcout(M_this_vga_signals_address_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGD3HC3_9_LC_24_31_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGD3HC3_9_LC_24_31_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGD3HC3_9_LC_24_31_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGD3HC3_9_LC_24_31_7  (
            .in0(N__20334),
            .in1(N__20168),
            .in2(_gnd_net_),
            .in3(N__20135),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_address_ibuf_RNIPG5P_5_LC_32_21_6.C_ON=1'b0;
    defparam port_address_ibuf_RNIPG5P_5_LC_32_21_6.SEQ_MODE=4'b0000;
    defparam port_address_ibuf_RNIPG5P_5_LC_32_21_6.LUT_INIT=16'b0000000001010101;
    LogicCell40 port_address_ibuf_RNIPG5P_5_LC_32_21_6 (
            .in0(N__20024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20018),
            .lcout(M_state_q_ns_0_a3_0_0_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_address_ibuf_RNI7ITU1_2_LC_32_23_2.C_ON=1'b0;
    defparam port_address_ibuf_RNI7ITU1_2_LC_32_23_2.SEQ_MODE=4'b0000;
    defparam port_address_ibuf_RNI7ITU1_2_LC_32_23_2.LUT_INIT=16'b0000000100000000;
    LogicCell40 port_address_ibuf_RNI7ITU1_2_LC_32_23_2 (
            .in0(N__20006),
            .in1(N__19994),
            .in2(N__19982),
            .in3(N__19973),
            .lcout(M_state_q_ns_0_a3_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
