-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 28 2022 16:04:31

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    led : out std_logic_vector(7 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__36351\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \this_vga_signals.N_692_0\ : std_logic;
signal port_clk_c : std_logic;
signal port_data_rw_0_i : std_logic;
signal port_nmib_0_i : std_logic;
signal this_vga_signals_vvisibility_i : std_logic;
signal rgb_c_0 : std_logic;
signal rgb_c_1 : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.g0_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_1_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_0\ : std_logic;
signal \this_vga_signals.N_4_0_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_1_cascade_\ : std_logic;
signal \this_vga_signals.g2_1_cascade_\ : std_logic;
signal \this_vga_signals.g2\ : std_logic;
signal \this_vga_signals.vsync_1_3_cascade_\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \this_vga_signals.g0_2_0_cascade_\ : std_logic;
signal \this_vga_signals.N_43_1_cascade_\ : std_logic;
signal \this_vga_signals.un2_vsynclt8\ : std_logic;
signal \this_vga_signals.vsync_1_2\ : std_logic;
signal \this_vga_signals.g1_1\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \this_vga_signals.g0_0_0\ : std_logic;
signal \M_this_map_address_qZ0Z_0\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \M_this_map_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_map_address_q_cry_0\ : std_logic;
signal \M_this_map_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_map_address_q_cry_1\ : std_logic;
signal \M_this_map_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_map_address_q_cry_2\ : std_logic;
signal \M_this_map_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_map_address_q_cry_3\ : std_logic;
signal \M_this_map_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_map_address_q_cry_4\ : std_logic;
signal \M_this_map_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_5\ : std_logic;
signal \M_this_map_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_map_address_q_cry_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_7\ : std_logic;
signal \M_this_map_address_qZ0Z_8\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \un1_M_this_map_address_q_cry_8\ : std_logic;
signal \M_this_map_address_qZ0Z_9\ : std_logic;
signal \N_89_0\ : std_logic;
signal \N_83_0\ : std_logic;
signal \N_85_0\ : std_logic;
signal \this_vga_signals.vaddress_3_0_5_cascade_\ : std_logic;
signal \this_vga_signals.g0_6_0_0_0\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_1_3_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_1_1_3\ : std_logic;
signal \this_vga_signals.N_1_3_1\ : std_logic;
signal \this_vga_signals.N_1_3_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.vaddress_1_0_5_cascade_\ : std_logic;
signal \this_vga_signals.un6_vvisibilitylt8_cascade_\ : std_logic;
signal \this_vga_signals.vvisibility_1\ : std_logic;
signal \this_vga_signals.vaddress_0_5\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_3_cascade_\ : std_logic;
signal \this_vga_signals.g0_6_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d\ : std_logic;
signal \this_vga_signals.i6_mux_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_a2_1\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_2\ : std_logic;
signal \this_vga_signals.SUM_3_1_tz\ : std_logic;
signal this_vga_signals_hvisibility_i : std_logic;
signal \M_stage_q_RNIC68K4_9\ : std_logic;
signal \this_vga_signals.vaddress_3_5\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_5_cascade_\ : std_logic;
signal \this_vga_signals.g0_6_0_0\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_0\ : std_logic;
signal \this_vga_signals.N_5_i_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.M_vcounter_q_8_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_9_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_c2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_0\ : std_logic;
signal \this_vga_signals.vaddress_2_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_x0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_1\ : std_logic;
signal \this_vga_signals.if_N_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_cascade_\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_6\ : std_logic;
signal \this_vga_signals.N_5_i_0\ : std_logic;
signal \this_vga_signals.g1_2_1_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_4_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_2_0\ : std_logic;
signal \this_vga_signals.g1_0_4\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_4\ : std_logic;
signal \this_vga_signals.g1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_1_0_0_0\ : std_logic;
signal \this_vga_signals.g2_1_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g3_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0_0\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lt7_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3_0_1_cascade_\ : std_logic;
signal \this_vga_signals.haddress_1_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lto7_1\ : std_logic;
signal \this_vga_signals.un2_hsynclto3_0\ : std_logic;
signal \this_vga_signals.un2_hsynclto3_0_cascade_\ : std_logic;
signal \this_vga_signals.un2_hsynclto6_0_cascade_\ : std_logic;
signal rgb_c_4 : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal \this_vga_signals.N_692_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_379_0\ : std_logic;
signal \this_vga_signals.g0_3_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_0\ : std_logic;
signal \this_vga_signals.g1_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_0\ : std_logic;
signal \this_vga_signals.g1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1\ : std_logic;
signal \this_vga_signals.g0_1_0_0\ : std_logic;
signal \this_vga_signals.g1_2_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_0_0_0\ : std_logic;
signal \this_vga_signals.g0_2_0_a2_1\ : std_logic;
signal \this_vga_signals.g0_2_0_a2_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_3_x1\ : std_logic;
signal \this_vga_signals.g0_13_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_2_cascade_\ : std_logic;
signal \this_vga_signals.g0_13_x1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_x0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_x1\ : std_logic;
signal \this_vga_signals.g1_2_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNITVMCUZ0Z_3_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNIANU4QZ0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_2\ : std_logic;
signal \this_vga_signals.g2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_0_a3_0\ : std_logic;
signal \this_vga_signals.vaddress_c3_0\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_1_3\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_2_3\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_0\ : std_logic;
signal \this_vga_signals.g0_i_x4_4_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_4\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \this_vga_signals.g2_0\ : std_logic;
signal \this_vga_signals.g0_2_0_a2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_ns\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_571\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3\ : std_logic;
signal \this_vga_signals.N_4_0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_cascade_\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \this_vga_signals.if_m2_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb2_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \this_vga_signals.SUM_3\ : std_logic;
signal \this_vga_signals.SUM_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0\ : std_logic;
signal \this_vga_signals.N_6_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_0_0_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.un4_hsynclt4_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \N_91_0\ : std_logic;
signal \N_93_0\ : std_logic;
signal \M_this_map_ram_read_data_3\ : std_logic;
signal \M_this_ppu_sprites_addr_9\ : std_logic;
signal \M_this_map_ram_read_data_0\ : std_logic;
signal \M_this_ppu_sprites_addr_6\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.N_692_0_g\ : std_logic;
signal \this_vga_signals.N_988_g\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.un4_hsynclt8_0\ : std_logic;
signal \this_vga_signals.un2_hsynclt8_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal this_vga_signals_hsync_1_i : std_logic;
signal rgb_c_3 : std_logic;
signal \N_95_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \M_this_map_ram_read_data_2\ : std_logic;
signal \M_this_ppu_sprites_addr_8\ : std_logic;
signal \this_vga_ramdac.N_24_mux\ : std_logic;
signal \this_vga_ramdac.N_2862_reto\ : std_logic;
signal \this_pixel_clk_M_counter_q_i_1\ : std_logic;
signal rgb_c_2 : std_logic;
signal \this_vga_ramdac.m6\ : std_logic;
signal \this_vga_ramdac.N_2863_reto\ : std_logic;
signal \this_vga_ramdac.i2_mux_0\ : std_logic;
signal \this_vga_ramdac.m19\ : std_logic;
signal \this_vga_ramdac.N_2866_reto\ : std_logic;
signal \this_vga_signals.M_this_vga_signals_pixel_clk_0_0\ : std_logic;
signal \M_this_vga_ramdac_en_0\ : std_logic;
signal \M_pcounter_q_ret_2_RNIH7PG8_cascade_\ : std_logic;
signal \this_vga_ramdac.i2_mux\ : std_logic;
signal \this_vga_ramdac.N_2864_reto\ : std_logic;
signal dma_0_i : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_0\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_1\ : std_logic;
signal \this_vga_signals.N_3_0\ : std_logic;
signal \this_vga_signals.N_3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_3_1\ : std_logic;
signal \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\ : std_logic;
signal \this_vga_ramdac.N_2867_reto\ : std_logic;
signal rgb_c_5 : std_logic;
signal \this_vga_signals.N_2_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_3_0\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \M_this_data_count_q_cry_0\ : std_logic;
signal \M_this_data_count_q_cry_1\ : std_logic;
signal \M_this_data_count_q_cry_2\ : std_logic;
signal \M_this_data_count_q_cry_3\ : std_logic;
signal \M_this_data_count_q_cry_4\ : std_logic;
signal \M_this_data_count_q_cry_5\ : std_logic;
signal \M_this_data_count_q_cry_6\ : std_logic;
signal \M_this_data_count_q_cry_7\ : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal \M_this_data_count_q_cry_8\ : std_logic;
signal \M_this_data_count_q_s_10\ : std_logic;
signal \M_this_data_count_q_cry_9\ : std_logic;
signal \M_this_data_count_q_cry_10\ : std_logic;
signal \M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_data_count_q_cry_12\ : std_logic;
signal \M_this_data_count_q_s_13\ : std_logic;
signal \N_87_0\ : std_logic;
signal \N_81_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt8_0\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lto8_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_d8_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\ : std_logic;
signal \this_pixel_clk_M_counter_q_0\ : std_logic;
signal \M_pcounter_q_ret_2_RNIH7PG8\ : std_logic;
signal \this_vga_ramdac.N_2865_reto\ : std_logic;
signal \dma_ac0_5_0_cascade_\ : std_logic;
signal \M_this_state_q_RNIOE1SZ0Z_11\ : std_logic;
signal un20_i_a2_x_3 : std_logic;
signal \M_this_state_q_RNIG01LZ0Z_12\ : std_logic;
signal \this_vga_signals.N_419_i_i_0Z0Z_1_cascade_\ : std_logic;
signal \M_this_data_count_q_s_6\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \M_this_data_count_q_cry_3_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \M_this_data_count_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \M_this_data_count_q_cry_2_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_10_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_11_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \M_this_data_count_q_cry_7_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \M_this_data_count_q_cry_1_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_8_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \M_this_map_ram_read_data_1\ : std_logic;
signal \M_this_ppu_sprites_addr_7\ : std_logic;
signal \this_ppu.M_count_d_0_sqmuxa_1_7_cascade_\ : std_logic;
signal \this_vga_signals.un4_lvisibility_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_6_s1\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_7\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_5\ : std_logic;
signal \this_ppu.M_count_qZ0Z_4\ : std_logic;
signal \this_ppu.M_count_qZ0Z_6\ : std_logic;
signal \this_ppu.M_count_qZ0Z_2\ : std_logic;
signal \this_ppu.M_count_d_1_sqmuxa_1_i_a2_4\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \this_vga_signals.un20_i_a2_sxZ0Z_3_cascade_\ : std_logic;
signal \this_vga_signals.N_322_cascade_\ : std_logic;
signal \this_vga_signals_M_this_state_q_ns_i_o3_0_10\ : std_logic;
signal \M_this_state_qZ0Z_10\ : std_logic;
signal \N_212\ : std_logic;
signal \N_160_0\ : std_logic;
signal \M_this_state_qc_3_1\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_4_cascade_\ : std_logic;
signal \N_465_0\ : std_logic;
signal \N_610_0_i\ : std_logic;
signal \M_this_data_count_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_data_count_qe_0_i\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_this_state_d55Z0Z_9\ : std_logic;
signal \this_vga_signals.M_this_state_d55Z0Z_8\ : std_logic;
signal \this_vga_signals.M_this_state_d55Z0Z_7_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_d55Z0Z_6\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \this_vga_ramdac.m16\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_5\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_8\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_6\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_7\ : std_logic;
signal \this_ppu.M_count_qZ0Z_7\ : std_logic;
signal \this_ppu.M_count_d_1_sqmuxa_1_i_a2_3\ : std_logic;
signal \this_ppu.N_132_0_cascade_\ : std_logic;
signal \this_ppu.M_count_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_d8\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d7_1_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_d7_0\ : std_logic;
signal \this_vga_signals.GZ0Z_330\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d7_1_0\ : std_logic;
signal \this_vga_signals.CO0_cascade_\ : std_logic;
signal \this_ppu.N_1157_0_1\ : std_logic;
signal \this_ppu.un16_0\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\ : std_logic;
signal \this_ppu.un16_0_cascade_\ : std_logic;
signal \this_ppu.N_1157_0\ : std_logic;
signal \this_ppu.M_count_qZ0Z_3\ : std_logic;
signal \N_459_0_cascade_\ : std_logic;
signal \N_458_0_cascade_\ : std_logic;
signal \this_vga_signals_N_419_i_i_0_a3_1_0\ : std_logic;
signal \N_496_0_cascade_\ : std_logic;
signal \N_278\ : std_logic;
signal \M_this_state_qsr_0_cascade_\ : std_logic;
signal \N_462_0\ : std_logic;
signal \M_this_state_qsr_2_cascade_\ : std_logic;
signal \N_484_0\ : std_logic;
signal \this_vga_signals.N_159_0_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_9\ : std_logic;
signal \N_168_0\ : std_logic;
signal \N_168_0_cascade_\ : std_logic;
signal \this_vga_signals.M_this_external_address_d_0_sqmuxa_1Z0Z_2\ : std_logic;
signal \M_this_state_qZ0Z_11\ : std_logic;
signal \N_456_0_1\ : std_logic;
signal \N_500\ : std_logic;
signal \M_this_sprites_ram_write_data_0\ : std_logic;
signal \M_this_state_d_2_sqmuxa\ : std_logic;
signal \M_this_substate_qZ0\ : std_logic;
signal \this_vga_signals_M_this_state_q_ns_0_a3_0_0_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_0\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_3\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_4\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_2\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\ : std_logic;
signal \M_this_map_ram_read_data_7\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_2\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.line_clk_1\ : std_logic;
signal \M_this_sprites_ram_write_data_3\ : std_logic;
signal \this_vga_signals.N_169_0\ : std_logic;
signal \N_210_cascade_\ : std_logic;
signal \this_vga_signals.N_159_0\ : std_logic;
signal \this_vga_signals.N_167_0_cascade_\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_5_cascade_\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_6\ : std_logic;
signal \M_this_state_d55\ : std_logic;
signal \this_vga_signals_M_this_state_q_ns_i_o3_0_7_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0\ : std_logic;
signal \this_vga_signals.N_279\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \N_210\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \this_vga_signals.N_166\ : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_1\ : std_logic;
signal \M_this_map_ram_read_data_5\ : std_logic;
signal \M_this_ppu_vram_data_3\ : std_logic;
signal \M_this_ppu_vram_data_2\ : std_logic;
signal \M_this_ppu_vram_data_3_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_0\ : std_logic;
signal \this_ppu.N_156_cascade_\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_2\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_3_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_3_c5\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_3\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_3\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_start_data_delay_M_last_q\ : std_logic;
signal port_enb_c : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal \N_156_0_cascade_\ : std_logic;
signal \N_35_0\ : std_logic;
signal port_rw_in : std_logic;
signal led_c_1 : std_logic;
signal \N_459_0\ : std_logic;
signal \un1_M_this_state_q_12_0\ : std_logic;
signal \bfn_19_22_0_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3\ : std_logic;
signal \M_this_sprites_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4\ : std_logic;
signal \M_this_sprites_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7\ : std_logic;
signal \bfn_19_23_0_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12\ : std_logic;
signal \M_this_state_d25\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_9_cascade_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_2_cascade_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3_cascade_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_7\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\ : std_logic;
signal \M_this_ppu_vram_data_1\ : std_logic;
signal \this_sprites_ram.mem_WE_14\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_1\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_3\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\ : std_logic;
signal this_vga_signals_vvisibility : std_logic;
signal dma_0 : std_logic;
signal \this_ppu.N_150_cascade_\ : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal \M_this_ppu_sprites_addr_2\ : std_logic;
signal \M_this_ppu_vram_en_0\ : std_logic;
signal \this_ppu.N_156\ : std_logic;
signal \this_ppu.un2_hscroll_axb_0_cascade_\ : std_logic;
signal \M_this_ppu_sprites_addr_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_3_c2\ : std_logic;
signal \this_ppu.M_state_q_RNIGL6V4Z0Z_0\ : std_logic;
signal \this_sprites_ram.mem_WE_8\ : std_logic;
signal \this_ppu.N_1046_0_cascade_\ : std_logic;
signal \this_ppu.M_state_qZ0Z_5\ : std_logic;
signal \this_ppu.un1_M_oam_idx_q_1_c1_cascade_\ : std_logic;
signal \this_ppu.un1_M_oam_idx_q_1_c3\ : std_logic;
signal \M_this_ppu_oam_addr_2\ : std_logic;
signal \M_this_ppu_oam_addr_0\ : std_logic;
signal \this_ppu.M_oam_idx_qZ0Z_4\ : std_logic;
signal \this_ppu.N_144_4_cascade_\ : std_logic;
signal \this_ppu.M_state_qZ0Z_4\ : std_logic;
signal \this_ppu.N_1046_0\ : std_logic;
signal \this_ppu.un1_M_oam_idx_q_1_c1\ : std_logic;
signal \M_this_ppu_oam_addr_1\ : std_logic;
signal \M_this_ppu_oam_addr_3\ : std_logic;
signal \this_ppu.N_144_4\ : std_logic;
signal \this_ppu.N_144\ : std_logic;
signal \M_this_state_qZ0Z_8\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal \M_this_sprites_ram_write_data_2\ : std_logic;
signal \this_sprites_ram.mem_WE_6\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0\ : std_logic;
signal \M_this_sprites_address_q_RNIQ61C7Z0Z_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_11\ : std_logic;
signal \M_this_substate_q_RNOZ0Z_1\ : std_logic;
signal \M_this_substate_q_s_1\ : std_logic;
signal \this_vga_signals_M_this_state_d_2_sqmuxa_0\ : std_logic;
signal \N_17_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_3\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_12\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_13\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_10_cascade_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_10\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10\ : std_logic;
signal \M_this_substate_q_RNOZ0Z_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_1\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_11\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_1\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\ : std_logic;
signal \bfn_21_16_0_\ : std_logic;
signal \this_ppu.un2_hscroll_cry_0\ : std_logic;
signal \this_ppu.un2_hscroll_cry_1\ : std_logic;
signal \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0\ : std_logic;
signal \this_sprites_ram.mem_WE_12\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_2\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\ : std_logic;
signal \M_this_oam_ram_read_data_i_9\ : std_logic;
signal \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0\ : std_logic;
signal \M_this_ppu_sprites_addr_1\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \bfn_21_18_0_\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_0\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_1\ : std_logic;
signal \M_this_oam_ram_read_data_i_11\ : std_logic;
signal \M_this_ppu_map_addr_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_4\ : std_logic;
signal \M_this_ppu_map_addr_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_3\ : std_logic;
signal \M_this_ppu_map_addr_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_4\ : std_logic;
signal \M_this_ppu_map_addr_3\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_5\ : std_logic;
signal \M_this_ppu_map_addr_4\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_6\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_7\ : std_logic;
signal \bfn_21_19_0_\ : std_logic;
signal \this_ppu.vscroll8\ : std_logic;
signal \this_ppu.M_state_qZ0Z_2\ : std_logic;
signal \N_48_0\ : std_logic;
signal \M_this_oam_ram_write_data_28\ : std_logic;
signal \this_ppu.M_state_qZ0Z_3\ : std_logic;
signal \this_ppu.M_state_qZ0Z_1\ : std_logic;
signal \this_ppu.M_count_d_0_sqmuxa_1_7\ : std_logic;
signal \this_ppu.N_148\ : std_logic;
signal \M_this_data_tmp_qZ0Z_20\ : std_logic;
signal \this_sprites_ram.mem_WE_4\ : std_logic;
signal \M_this_state_d22\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11\ : std_logic;
signal port_address_in_0 : std_logic;
signal \this_vga_signals.M_this_state_d21Z0Z_6\ : std_logic;
signal \this_vga_signals.M_this_state_dZ0Z24\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_8\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_8\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_1_cascade_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4\ : std_logic;
signal \this_vga_signals.un1_M_this_state_q_14_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_mZ0Z_4\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_8\ : std_logic;
signal \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\ : std_logic;
signal \M_this_sprites_ram_write_data_1\ : std_logic;
signal \M_this_map_ram_read_data_4\ : std_logic;
signal \M_this_ppu_sprites_addr_10\ : std_logic;
signal \M_this_ppu_sprites_addr_4\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_2_c5\ : std_logic;
signal \bfn_22_17_0_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_0\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_1\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_2\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_3\ : std_logic;
signal \M_this_ppu_map_addr_7\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_4\ : std_logic;
signal \M_this_ppu_map_addr_8\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_5\ : std_logic;
signal \M_this_ppu_map_addr_9\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_7\ : std_logic;
signal \bfn_22_18_0_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_5\ : std_logic;
signal \un1_M_this_oam_address_q_c3_cascade_\ : std_logic;
signal \M_this_data_tmp_qZ0Z_7\ : std_logic;
signal \N_65_0\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_0\ : std_logic;
signal \M_this_oam_ram_read_data_8\ : std_logic;
signal \bfn_22_19_0_\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_1\ : std_logic;
signal \M_this_oam_ram_read_data_9\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_0\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_2\ : std_logic;
signal \M_this_oam_ram_read_data_10\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_1\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_2\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_3\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_4\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_3\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_5\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_4\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_6\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_7\ : std_logic;
signal \bfn_22_20_0_\ : std_logic;
signal \this_ppu.vscroll8_1\ : std_logic;
signal port_address_in_5 : std_logic;
signal port_address_in_6 : std_logic;
signal port_address_in_7 : std_logic;
signal \M_this_state_qZ0Z_12\ : std_logic;
signal \N_56_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_13\ : std_logic;
signal \M_this_state_d21_1\ : std_logic;
signal port_address_in_4 : std_logic;
signal port_address_in_2 : std_logic;
signal \M_this_state_d21_6_x\ : std_logic;
signal \M_this_substate_q_RNOZ0Z_2\ : std_logic;
signal port_address_in_3 : std_logic;
signal port_address_in_1 : std_logic;
signal \this_vga_signals.M_this_state_d24Z0Z_1\ : std_logic;
signal \this_sprites_ram.mem_WE_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_15\ : std_logic;
signal \M_this_oam_ram_write_data_15\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_16\ : std_logic;
signal \bfn_23_16_0_\ : std_logic;
signal \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0\ : std_logic;
signal \this_ppu.un2_vscroll_cry_0\ : std_logic;
signal \this_ppu.un2_vscroll_cry_1\ : std_logic;
signal \M_this_map_ram_read_data_6\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_12\ : std_logic;
signal \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0\ : std_logic;
signal \M_this_ppu_sprites_addr_5\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_1\ : std_logic;
signal \this_ppu.N_132_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_6\ : std_logic;
signal \this_ppu.un2_vscroll_axb_0_cascade_\ : std_logic;
signal \this_ppu.M_state_qZ0Z_7\ : std_logic;
signal \M_this_ppu_sprites_addr_3\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_2\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_2_c2\ : std_logic;
signal \M_this_ppu_map_addr_5\ : std_logic;
signal \M_this_ppu_map_addr_6\ : std_logic;
signal \this_ppu.M_state_qZ0Z_0\ : std_logic;
signal \this_ppu.M_last_q\ : std_logic;
signal \M_this_vga_signals_line_clk_0\ : std_logic;
signal \M_this_ppu_vram_addr_7\ : std_logic;
signal \this_ppu.M_state_q_RNI42KTAZ0Z_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_4\ : std_logic;
signal \N_71_0\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_7\ : std_logic;
signal \M_this_oam_ram_read_data_16\ : std_logic;
signal \bfn_23_19_0_\ : std_logic;
signal \this_ppu.M_vaddress_q_i_1\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_0\ : std_logic;
signal \this_ppu.M_vaddress_q_i_2\ : std_logic;
signal \M_this_oam_ram_read_data_18\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_1\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_5\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_2\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_3\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_7\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_4\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_8\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_5\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_9\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_7\ : std_logic;
signal \bfn_23_20_0_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_7_THRU_CO\ : std_logic;
signal \N_61_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_3\ : std_logic;
signal \N_73_0\ : std_logic;
signal \M_this_oam_address_qZ0Z_4\ : std_logic;
signal \M_this_oam_address_qZ0Z_5\ : std_logic;
signal \N_1152_0\ : std_logic;
signal \M_this_oam_address_qZ0Z_3\ : std_logic;
signal \M_this_oam_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_oam_address_q_c2\ : std_logic;
signal \un1_M_this_oam_address_q_c4\ : std_logic;
signal \N_50_0\ : std_logic;
signal \N_46_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_21\ : std_logic;
signal \M_this_data_tmp_qZ0Z_10\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_3\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_WE_10\ : std_logic;
signal \M_this_oam_ram_read_data_17\ : std_logic;
signal \M_this_oam_ram_read_data_i_17\ : std_logic;
signal \M_this_oam_ram_read_data_2\ : std_logic;
signal \M_this_oam_ram_read_data_1\ : std_logic;
signal \M_this_oam_ram_read_data_0\ : std_logic;
signal \M_this_oam_ram_read_data_3\ : std_logic;
signal \this_ppu.un9lto7Z0Z_5\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_6\ : std_logic;
signal \M_this_oam_ram_read_data_4\ : std_logic;
signal \M_this_oam_ram_read_data_6\ : std_logic;
signal \M_this_oam_ram_read_data_7\ : std_logic;
signal \M_this_oam_ram_read_data_5\ : std_logic;
signal \this_ppu.un9lto7Z0Z_4\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_4\ : std_logic;
signal \M_this_oam_ram_read_data_11\ : std_logic;
signal \M_this_oam_ram_read_data_12\ : std_logic;
signal \M_this_oam_ram_read_data_15\ : std_logic;
signal \M_this_oam_ram_read_data_14\ : std_logic;
signal \this_ppu.un1_oam_data_1_c2_cascade_\ : std_logic;
signal \M_this_oam_ram_read_data_13\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_7\ : std_logic;
signal \M_this_data_tmp_qZ0Z_6\ : std_logic;
signal \N_67_0\ : std_logic;
signal \M_this_oam_ram_read_data_23\ : std_logic;
signal \this_ppu.un1_oam_data_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_7\ : std_logic;
signal \M_this_oam_ram_write_data_22\ : std_logic;
signal \M_this_oam_ram_read_data_22\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_6\ : std_logic;
signal \M_this_oam_ram_write_data_31\ : std_logic;
signal \N_52_0\ : std_logic;
signal \M_this_oam_ram_write_data_16\ : std_logic;
signal \N_158_0\ : std_logic;
signal \M_this_oam_ram_read_data_21\ : std_logic;
signal \M_this_oam_ram_read_data_20\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_5\ : std_logic;
signal \M_this_oam_ram_read_data_19\ : std_logic;
signal \M_this_oam_ram_read_data_i_19\ : std_logic;
signal \M_this_data_tmp_qZ0Z_16\ : std_logic;
signal \M_this_data_tmp_qZ0Z_19\ : std_logic;
signal \M_this_data_tmp_qZ0Z_18\ : std_logic;
signal \M_this_data_tmp_qZ0Z_22\ : std_logic;
signal \M_this_data_tmp_qZ0Z_17\ : std_logic;
signal \N_54_0\ : std_logic;
signal \N_1126_0\ : std_logic;
signal \M_this_oam_ram_write_data_30\ : std_logic;
signal \bfn_24_22_0_\ : std_logic;
signal \un1_M_this_external_address_q_cry_0\ : std_logic;
signal \un1_M_this_external_address_q_cry_1\ : std_logic;
signal \un1_M_this_external_address_q_cry_2\ : std_logic;
signal \un1_M_this_external_address_q_cry_3\ : std_logic;
signal \un1_M_this_external_address_q_cry_4\ : std_logic;
signal \un1_M_this_external_address_q_cry_5\ : std_logic;
signal \un1_M_this_external_address_q_cry_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_7\ : std_logic;
signal \bfn_24_23_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_external_address_q_cry_8_c_RNI09PBZ0\ : std_logic;
signal \un1_M_this_external_address_q_cry_8\ : std_logic;
signal \un1_M_this_external_address_q_cry_9\ : std_logic;
signal \un1_M_this_external_address_q_cry_10\ : std_logic;
signal \un1_M_this_external_address_q_cry_11\ : std_logic;
signal \un1_M_this_external_address_q_cry_12\ : std_logic;
signal \un1_M_this_external_address_q_cry_13\ : std_logic;
signal \un1_M_this_external_address_q_cry_14\ : std_logic;
signal \M_this_sprites_address_qZ0Z_12\ : std_logic;
signal \M_this_sprites_address_qZ0Z_11\ : std_logic;
signal \M_this_sprites_address_qZ0Z_13\ : std_logic;
signal \M_this_sprites_ram_write_en_0_0\ : std_logic;
signal \this_sprites_ram.mem_WE_2\ : std_logic;
signal \M_this_oam_ram_write_data_8\ : std_logic;
signal \M_this_data_tmp_qZ0Z_8\ : std_logic;
signal \N_79_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_0\ : std_logic;
signal \N_43_0\ : std_logic;
signal \N_77_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_1\ : std_logic;
signal \N_58_0\ : std_logic;
signal \M_this_oam_ram_write_data_14\ : std_logic;
signal \N_63_0\ : std_logic;
signal \N_75_0\ : std_logic;
signal \M_this_oam_ram_write_data_11\ : std_logic;
signal \M_this_data_tmp_qZ0Z_11\ : std_logic;
signal \M_this_data_tmp_qZ0Z_12\ : std_logic;
signal \M_this_data_tmp_qZ0Z_9\ : std_logic;
signal \M_this_data_tmp_qZ0Z_14\ : std_logic;
signal \N_1134_0\ : std_logic;
signal \N_39_0\ : std_logic;
signal \M_this_oam_ram_write_data_27\ : std_logic;
signal \M_this_data_tmp_qZ0Z_23\ : std_logic;
signal \M_this_oam_ram_write_data_23\ : std_logic;
signal port_data_c_1 : std_logic;
signal \N_41_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_2\ : std_logic;
signal \un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0\ : std_logic;
signal port_data_c_3 : std_logic;
signal \M_this_external_address_qZ0Z_11\ : std_logic;
signal \un1_M_this_external_address_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_external_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0\ : std_logic;
signal port_data_c_4 : std_logic;
signal \M_this_external_address_qZ0Z_12\ : std_logic;
signal \un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_13\ : std_logic;
signal \un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0\ : std_logic;
signal port_data_c_6 : std_logic;
signal \M_this_external_address_qZ0Z_14\ : std_logic;
signal \un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0\ : std_logic;
signal port_data_c_0 : std_logic;
signal \M_this_external_address_qZ0Z_8\ : std_logic;
signal port_data_c_7 : std_logic;
signal \un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0\ : std_logic;
signal \M_this_external_address_qZ0Z_15\ : std_logic;
signal \un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0\ : std_logic;
signal port_data_c_2 : std_logic;
signal \M_this_external_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_state_q_11_0_i\ : std_logic;
signal \M_this_external_address_qZ0Z_0\ : std_logic;
signal \un1_M_this_external_address_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_external_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_external_address_q_cry_1_THRU_CO\ : std_logic;
signal \M_this_external_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_external_address_q_cry_2_THRU_CO\ : std_logic;
signal \M_this_external_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_external_address_q_cry_3_THRU_CO\ : std_logic;
signal \M_this_external_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_external_address_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_external_address_qZ0Z_5\ : std_logic;
signal \N_458_0\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \un1_M_this_external_address_q_cry_5_THRU_CO\ : std_logic;
signal \M_this_external_address_qZ0Z_6\ : std_logic;
signal \M_this_oam_address_qZ0Z_1\ : std_logic;
signal \N_156_0\ : std_logic;
signal \M_this_oam_address_qZ0Z_0\ : std_logic;
signal \N_69_0\ : std_logic;
signal port_data_c_5 : std_logic;
signal \M_this_data_tmp_qZ0Z_5\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_0_c_g : std_logic;
signal \N_1142_0\ : std_logic;
signal \M_this_reset_cond_out_g_0\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_map_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    led <= led_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \M_this_map_ram_read_data_3\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_2\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_1\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_0\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&\N__27777\&\N__27825\&\N__27870\&\N__29529\&\N__29577\&\N__25155\&\N__25212\&\N__25272\&\N__25335\&\N__25416\;
    \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&\N__11496\&\N__11529\&\N__11559\&\N__11589\&\N__11268\&\N__11298\&\N__11328\&\N__11358\&\N__11388\&\N__11415\;
    \this_map_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&\N__11469\&'0'&'0'&'0'&\N__13761\&'0'&'0'&'0'&\N__13752\&'0'&'0'&'0'&\N__15501\&'0';
    \M_this_map_ram_read_data_7\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_6\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_5\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_4\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&\N__27771\&\N__27819\&\N__27864\&\N__29523\&\N__29571\&\N__25149\&\N__25206\&\N__25265\&\N__25325\&\N__25409\;
    \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&\N__11490\&\N__11523\&\N__11553\&\N__11583\&\N__11262\&\N__11292\&\N__11322\&\N__11352\&\N__11382\&\N__11409\;
    \this_map_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&\N__16158\&'0'&'0'&'0'&\N__11463\&'0'&'0'&'0'&\N__11457\&'0'&'0'&'0'&\N__16170\&'0';
    \M_this_oam_ram_read_data_15\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(15);
    \M_this_oam_ram_read_data_14\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(14);
    \M_this_oam_ram_read_data_13\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_oam_ram_read_data_12\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(12);
    \M_this_oam_ram_read_data_11\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \M_this_oam_ram_read_data_10\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(10);
    \M_this_oam_ram_read_data_9\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_8\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(8);
    \M_this_oam_ram_read_data_7\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_6\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_5\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_4\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_3\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_2\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_1\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_0\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23838\&\N__23469\&\N__23874\&\N__23427\;
    \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__30717\&\N__30198\&\N__30639\&\N__30597\;
    \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ <= \N__29064\&\N__32052\&\N__28605\&\N__32058\&\N__32235\&\N__30234\&\N__32247\&\N__32115\&\N__28056\&\N__30723\&\N__34782\&\N__29226\&\N__30210\&\N__32241\&\N__32073\&\N__32100\;
    \M_this_oam_ram_read_data_23\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_22\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_21\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_20\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_19\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_18\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_17\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_16\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23832\&\N__23463\&\N__23868\&\N__23421\;
    \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__30711\&\N__30192\&\N__30631\&\N__30591\;
    \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ <= \N__31332\&\N__31578\&\N__20772\&\N__25965\&\N__32121\&\N__32127\&\N__32865\&\N__32085\&\N__32994\&\N__31380\&\N__30522\&\N__25980\&\N__30531\&\N__31326\&\N__31455\&\N__31320\;
    \this_sprites_ram.mem_out_bus0_1\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_0\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__27154\&\N__13724\&\N__15127\&\N__17412\&\N__14489\&\N__28948\&\N__26996\&\N__29869\&\N__22800\&\N__25812\&\N__23346\;
    \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__24879\&\N__22558\&\N__26613\&\N__21982\&\N__21360\&\N__21565\&\N__27633\&\N__24163\&\N__22265\&\N__26223\&\N__24468\;
    \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27321\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19652\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus0_3\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_2\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__27204\&\N__13717\&\N__15088\&\N__17407\&\N__14502\&\N__28878\&\N__26986\&\N__29862\&\N__22740\&\N__25808\&\N__23339\;
    \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__24875\&\N__22559\&\N__26609\&\N__22008\&\N__21359\&\N__21564\&\N__27629\&\N__24164\&\N__22293\&\N__26222\&\N__24467\;
    \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19980\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23643\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_1\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_0\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__27196\&\N__13704\&\N__15132\&\N__17347\&\N__14496\&\N__28937\&\N__26985\&\N__29847\&\N__22794\&\N__25800\&\N__23338\;
    \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__24874\&\N__22560\&\N__26608\&\N__22007\&\N__21352\&\N__21563\&\N__27622\&\N__24165\&\N__22289\&\N__26215\&\N__24460\;
    \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27317\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19653\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_3\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_2\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__27175\&\N__13695\&\N__15128\&\N__17392\&\N__14470\&\N__28920\&\N__26960\&\N__29814\&\N__22793\&\N__25784\&\N__23314\;
    \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__24864\&\N__22561\&\N__26598\&\N__22024\&\N__21351\&\N__21566\&\N__27612\&\N__24166\&\N__22282\&\N__26214\&\N__24427\;
    \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19976\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23637\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_1\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_0\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__27144\&\N__13678\&\N__15118\&\N__17391\&\N__14495\&\N__28896\&\N__26946\&\N__29815\&\N__22775\&\N__25715\&\N__23313\;
    \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__24825\&\N__22568\&\N__26584\&\N__22023\&\N__21338\&\N__21538\&\N__27599\&\N__24182\&\N__22253\&\N__26201\&\N__24450\;
    \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27309\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19651\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_3\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_2\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__27131\&\N__13601\&\N__15117\&\N__17358\&\N__14494\&\N__28850\&\N__26907\&\N__29798\&\N__22774\&\N__25757\&\N__23272\;
    \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__24851\&\N__22571\&\N__26563\&\N__22032\&\N__21337\&\N__21537\&\N__27584\&\N__24178\&\N__22271\&\N__26200\&\N__24449\;
    \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19938\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23636\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_1\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_0\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__27080\&\N__13688\&\N__15093\&\N__17277\&\N__14460\&\N__28841\&\N__26859\&\N__29777\&\N__22741\&\N__25722\&\N__23271\;
    \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__24850\&\N__22572\&\N__26535\&\N__22031\&\N__21318\&\N__21578\&\N__27568\&\N__24183\&\N__22228\&\N__26178\&\N__24433\;
    \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27295\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19643\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_3\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_2\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__27119\&\N__13631\&\N__15056\&\N__17348\&\N__14487\&\N__28930\&\N__26897\&\N__29870\&\N__22770\&\N__25794\&\N__23332\;
    \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__24830\&\N__22569\&\N__26597\&\N__21972\&\N__21317\&\N__21572\&\N__27611\&\N__24176\&\N__22237\&\N__26199\&\N__24430\;
    \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19974\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23642\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_1\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_0\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__27182\&\N__13671\&\N__15057\&\N__17384\&\N__14488\&\N__28944\&\N__26970\&\N__29883\&\N__22771\&\N__25807\&\N__23333\;
    \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__24849\&\N__22552\&\N__26580\&\N__22000\&\N__21292\&\N__21576\&\N__27580\&\N__24159\&\N__22281\&\N__26198\&\N__24429\;
    \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27316\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19647\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_3\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_2\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__27200\&\N__13700\&\N__15075\&\N__17405\&\N__14483\&\N__28949\&\N__26990\&\N__29875\&\N__22772\&\N__25780\&\N__23334\;
    \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__24826\&\N__22553\&\N__26579\&\N__22022\&\N__21260\&\N__21577\&\N__27561\&\N__24177\&\N__22267\&\N__26197\&\N__24390\;
    \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19967\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23641\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_1\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_0\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__27201\&\N__13716\&\N__15092\&\N__17406\&\N__14500\&\N__28950\&\N__26991\&\N__29882\&\N__22773\&\N__25799\&\N__23345\;
    \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__24793\&\N__22478\&\N__26578\&\N__22021\&\N__21291\&\N__21579\&\N__27538\&\N__24130\&\N__22227\&\N__26196\&\N__24428\;
    \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27305\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19641\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_3\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_2\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__27165\&\N__13711\&\N__15038\&\N__17399\&\N__14469\&\N__28851\&\N__26947\&\N__29808\&\N__22757\&\N__25740\&\N__23288\;
    \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__24811\&\N__22570\&\N__26527\&\N__21955\&\N__21214\&\N__21550\&\N__27529\&\N__24133\&\N__22246\&\N__26147\&\N__24333\;
    \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19948\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23618\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_1\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_0\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__27189\&\N__13696\&\N__15106\&\N__17400\&\N__14501\&\N__28888\&\N__26977\&\N__29822\&\N__22785\&\N__25741\&\N__23324\;
    \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__24740\&\N__22442\&\N__26491\&\N__21931\&\N__21270\&\N__21570\&\N__27493\&\N__24098\&\N__22185\&\N__26139\&\N__24403\;
    \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27263\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19640\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_3\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_2\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__27202\&\N__13670\&\N__15107\&\N__17401\&\N__14464\&\N__28889\&\N__26978\&\N__29858\&\N__22786\&\N__25775\&\N__23325\;
    \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__24806\&\N__22554\&\N__26528\&\N__21927\&\N__21271\&\N__21571\&\N__27522\&\N__24132\&\N__22241\&\N__26140\&\N__24404\;
    \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19944\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23619\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_1\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_0\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__27164\&\N__13715\&\N__15125\&\N__17380\&\N__14465\&\N__28918\&\N__26992\&\N__29851\&\N__22798\&\N__25776\&\N__23343\;
    \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__24807\&\N__22520\&\N__26561\&\N__21932\&\N__21296\&\N__21548\&\N__27548\&\N__24131\&\N__22242\&\N__26176\&\N__24431\;
    \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27264\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19642\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_3\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_2\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__27203\&\N__13725\&\N__15126\&\N__17411\&\N__14490\&\N__28919\&\N__26997\&\N__29874\&\N__22799\&\N__25798\&\N__23344\;
    \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__24831\&\N__22548\&\N__26562\&\N__21954\&\N__21297\&\N__21549\&\N__27549\&\N__24155\&\N__22266\&\N__26177\&\N__24432\;
    \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19975\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23629\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__11079\&\N__11106\&\N__13428\&\N__11094\&\N__13194\&\N__11115\&\N__13104\&\N__12225\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__29337\&\N__25202\&\N__25268\&\N__25334\&\N__25412\&\N__25476\&\N__25533\&\N__25590\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20739\&\N__20721\&\N__21786\&\N__20694\;

    \this_map_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34586\,
            RE => \N__17947\,
            WCLKE => \N__18250\,
            WCLK => \N__34587\,
            WE => \N__17943\
        );

    \this_map_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34590\,
            RE => \N__17948\,
            WCLKE => \N__18261\,
            WCLK => \N__34591\,
            WE => \N__17989\
        );

    \this_oam_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34546\,
            RE => \N__17738\,
            WCLKE => \N__31314\,
            WCLK => \N__34547\,
            WE => \N__17923\
        );

    \this_oam_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34564\,
            RE => \N__17898\,
            WCLKE => \N__31310\,
            WCLK => \N__34565\,
            WE => \N__17905\
        );

    \this_sprites_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34467\,
            RE => \N__17992\,
            WCLKE => \N__23085\,
            WCLK => \N__34468\,
            WE => \N__17922\
        );

    \this_sprites_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34469\,
            RE => \N__17849\,
            WCLKE => \N__23084\,
            WCLK => \N__34470\,
            WE => \N__17964\
        );

    \this_sprites_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34471\,
            RE => \N__17959\,
            WCLKE => \N__25092\,
            WCLK => \N__34472\,
            WE => \N__17963\
        );

    \this_sprites_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34481\,
            RE => \N__17752\,
            WCLKE => \N__25088\,
            WCLK => \N__34480\,
            WE => \N__17906\
        );

    \this_sprites_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34495\,
            RE => \N__18019\,
            WCLKE => \N__30357\,
            WCLK => \N__34496\,
            WE => \N__18010\
        );

    \this_sprites_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34511\,
            RE => \N__17739\,
            WCLKE => \N__30356\,
            WCLK => \N__34512\,
            WE => \N__18006\
        );

    \this_sprites_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34531\,
            RE => \N__17957\,
            WCLKE => \N__23114\,
            WCLK => \N__34532\,
            WE => \N__17934\
        );

    \this_sprites_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34522\,
            RE => \N__17991\,
            WCLKE => \N__23118\,
            WCLK => \N__34523\,
            WE => \N__17956\
        );

    \this_sprites_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34553\,
            RE => \N__17768\,
            WCLKE => \N__23571\,
            WCLK => \N__34554\,
            WE => \N__17884\
        );

    \this_sprites_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34571\,
            RE => \N__17864\,
            WCLKE => \N__23570\,
            WCLK => \N__34572\,
            WE => \N__17894\
        );

    \this_sprites_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34578\,
            RE => \N__17865\,
            WCLKE => \N__26793\,
            WCLK => \N__34579\,
            WE => \N__17942\
        );

    \this_sprites_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34573\,
            RE => \N__17765\,
            WCLKE => \N__26786\,
            WCLK => \N__34574\,
            WE => \N__17968\
        );

    \this_sprites_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34582\,
            RE => \N__17958\,
            WCLKE => \N__31592\,
            WCLK => \N__34583\,
            WE => \N__17996\
        );

    \this_sprites_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34588\,
            RE => \N__17766\,
            WCLKE => \N__31593\,
            WCLK => \N__34589\,
            WE => \N__17997\
        );

    \this_sprites_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34593\,
            RE => \N__18012\,
            WCLKE => \N__28313\,
            WCLK => \N__34594\,
            WE => \N__18020\
        );

    \this_sprites_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34595\,
            RE => \N__17767\,
            WCLKE => \N__28314\,
            WCLK => \N__34596\,
            WE => \N__18021\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34539\,
            RE => \N__17803\,
            WCLKE => \N__22614\,
            WCLK => \N__34540\,
            WE => \N__17952\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__36349\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36351\,
            DIN => \N__36350\,
            DOUT => \N__36349\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36351\,
            PADOUT => \N__36350\,
            PADIN => \N__36349\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36340\,
            DIN => \N__36339\,
            DOUT => \N__36338\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36340\,
            PADOUT => \N__36339\,
            PADIN => \N__36338\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36331\,
            DIN => \N__36330\,
            DOUT => \N__36329\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36331\,
            PADOUT => \N__36330\,
            PADIN => \N__36329\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36322\,
            DIN => \N__36321\,
            DOUT => \N__36320\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36322\,
            PADOUT => \N__36321\,
            PADIN => \N__36320\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11760\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36313\,
            DIN => \N__36312\,
            DOUT => \N__36311\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36313\,
            PADOUT => \N__36312\,
            PADIN => \N__36311\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14541\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36304\,
            DIN => \N__36303\,
            DOUT => \N__36302\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36304\,
            PADOUT => \N__36303\,
            PADIN => \N__36302\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__18011\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36295\,
            DIN => \N__36294\,
            DOUT => \N__36293\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36295\,
            PADOUT => \N__36294\,
            PADIN => \N__36293\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21699\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36286\,
            DIN => \N__36285\,
            DOUT => \N__36284\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36286\,
            PADOUT => \N__36285\,
            PADIN => \N__36284\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36277\,
            DIN => \N__36276\,
            DOUT => \N__36275\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36277\,
            PADOUT => \N__36276\,
            PADIN => \N__36275\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36268\,
            DIN => \N__36267\,
            DOUT => \N__36266\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36268\,
            PADOUT => \N__36267\,
            PADIN => \N__36266\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36259\,
            DIN => \N__36258\,
            DOUT => \N__36257\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36259\,
            PADOUT => \N__36258\,
            PADIN => \N__36257\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36250\,
            DIN => \N__36249\,
            DOUT => \N__36248\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36250\,
            PADOUT => \N__36249\,
            PADIN => \N__36248\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36241\,
            DIN => \N__36240\,
            DOUT => \N__36239\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36241\,
            PADOUT => \N__36240\,
            PADIN => \N__36239\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36232\,
            DIN => \N__36231\,
            DOUT => \N__36230\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36232\,
            PADOUT => \N__36231\,
            PADIN => \N__36230\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__33279\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16000\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36223\,
            DIN => \N__36222\,
            DOUT => \N__36221\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36223\,
            PADOUT => \N__36222\,
            PADIN => \N__36221\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__33221\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15989\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36214\,
            DIN => \N__36213\,
            DOUT => \N__36212\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36214\,
            PADOUT => \N__36213\,
            PADIN => \N__36212\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__33180\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16056\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36205\,
            DIN => \N__36204\,
            DOUT => \N__36203\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36205\,
            PADOUT => \N__36204\,
            PADIN => \N__36203\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__33132\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16096\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36196\,
            DIN => \N__36195\,
            DOUT => \N__36194\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36196\,
            PADOUT => \N__36195\,
            PADIN => \N__36194\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__33083\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16083\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36187\,
            DIN => \N__36186\,
            DOUT => \N__36185\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36187\,
            PADOUT => \N__36186\,
            PADIN => \N__36185\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__33042\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16061\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36178\,
            DIN => \N__36177\,
            DOUT => \N__36176\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36178\,
            PADOUT => \N__36177\,
            PADIN => \N__36176\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__35526\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16097\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36169\,
            DIN => \N__36168\,
            DOUT => \N__36167\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36169\,
            PADOUT => \N__36168\,
            PADIN => \N__36167\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__32652\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16094\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36160\,
            DIN => \N__36159\,
            DOUT => \N__36158\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36160\,
            PADOUT => \N__36159\,
            PADIN => \N__36158\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__33330\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16027\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36151\,
            DIN => \N__36150\,
            DOUT => \N__36149\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36151\,
            PADOUT => \N__36150\,
            PADIN => \N__36149\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__32691\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16095\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36142\,
            DIN => \N__36141\,
            DOUT => \N__36140\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36142\,
            PADOUT => \N__36141\,
            PADIN => \N__36140\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__32481\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16084\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36133\,
            DIN => \N__36132\,
            DOUT => \N__36131\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36133\,
            PADOUT => \N__36132\,
            PADIN => \N__36131\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__32445\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16062\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36124\,
            DIN => \N__36123\,
            DOUT => \N__36122\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36124\,
            PADOUT => \N__36123\,
            PADIN => \N__36122\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__32277\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16098\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36115\,
            DIN => \N__36114\,
            DOUT => \N__36113\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36115\,
            PADOUT => \N__36114\,
            PADIN => \N__36113\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__33534\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16022\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36106\,
            DIN => \N__36105\,
            DOUT => \N__36104\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36106\,
            PADOUT => \N__36105\,
            PADIN => \N__36104\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__33696\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15999\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36097\,
            DIN => \N__36096\,
            DOUT => \N__36095\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__36097\,
            PADOUT => \N__36096\,
            PADIN => \N__36095\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__32043\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16057\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36088\,
            DIN => \N__36087\,
            DOUT => \N__36086\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36088\,
            PADOUT => \N__36087\,
            PADIN => \N__36086\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36079\,
            DIN => \N__36078\,
            DOUT => \N__36077\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36079\,
            PADOUT => \N__36078\,
            PADIN => \N__36077\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36070\,
            DIN => \N__36069\,
            DOUT => \N__36068\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36070\,
            PADOUT => \N__36069\,
            PADIN => \N__36068\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36061\,
            DIN => \N__36060\,
            DOUT => \N__36059\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36061\,
            PADOUT => \N__36060\,
            PADIN => \N__36059\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36052\,
            DIN => \N__36051\,
            DOUT => \N__36050\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36052\,
            PADOUT => \N__36051\,
            PADIN => \N__36050\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36043\,
            DIN => \N__36042\,
            DOUT => \N__36041\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36043\,
            PADOUT => \N__36042\,
            PADIN => \N__36041\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36034\,
            DIN => \N__36033\,
            DOUT => \N__36032\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36034\,
            PADOUT => \N__36033\,
            PADIN => \N__36032\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36025\,
            DIN => \N__36024\,
            DOUT => \N__36023\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36025\,
            PADOUT => \N__36024\,
            PADIN => \N__36023\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36016\,
            DIN => \N__36015\,
            DOUT => \N__36014\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36016\,
            PADOUT => \N__36015\,
            PADIN => \N__36014\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36007\,
            DIN => \N__36006\,
            DOUT => \N__36005\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36007\,
            PADOUT => \N__36006\,
            PADIN => \N__36005\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11058\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35998\,
            DIN => \N__35997\,
            DOUT => \N__35996\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35998\,
            PADOUT => \N__35997\,
            PADIN => \N__35996\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__22941\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35989\,
            DIN => \N__35988\,
            DOUT => \N__35987\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35989\,
            PADOUT => \N__35988\,
            PADIN => \N__35987\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35980\,
            DIN => \N__35979\,
            DOUT => \N__35978\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35980\,
            PADOUT => \N__35979\,
            PADIN => \N__35978\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11052\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35971\,
            DIN => \N__35970\,
            DOUT => \N__35969\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35971\,
            PADOUT => \N__35970\,
            PADIN => \N__35969\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__17990\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16026\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35962\,
            DIN => \N__35961\,
            DOUT => \N__35960\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35962\,
            PADOUT => \N__35961\,
            PADIN => \N__35960\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11139\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35953\,
            DIN => \N__35952\,
            DOUT => \N__35951\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35953\,
            PADOUT => \N__35952\,
            PADIN => \N__35951\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11124\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35944\,
            DIN => \N__35943\,
            DOUT => \N__35942\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35944\,
            PADOUT => \N__35943\,
            PADIN => \N__35942\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15693\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35935\,
            DIN => \N__35934\,
            DOUT => \N__35933\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35935\,
            PADOUT => \N__35934\,
            PADIN => \N__35933\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15522\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35926\,
            DIN => \N__35925\,
            DOUT => \N__35924\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35926\,
            PADOUT => \N__35925\,
            PADIN => \N__35924\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12309\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35917\,
            DIN => \N__35916\,
            DOUT => \N__35915\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35917\,
            PADOUT => \N__35916\,
            PADIN => \N__35915\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15750\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35908\,
            DIN => \N__35907\,
            DOUT => \N__35906\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35908\,
            PADOUT => \N__35907\,
            PADIN => \N__35906\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35899\,
            DIN => \N__35898\,
            DOUT => \N__35897\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35899\,
            PADOUT => \N__35898\,
            PADIN => \N__35897\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11037\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35890\,
            DIN => \N__35889\,
            DOUT => \N__35888\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35890\,
            PADOUT => \N__35889\,
            PADIN => \N__35888\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11235\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__9096\ : CascadeMux
    port map (
            O => \N__35871\,
            I => \N__35868\
        );

    \I__9095\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35847\
        );

    \I__9094\ : InMux
    port map (
            O => \N__35867\,
            I => \N__35829\
        );

    \I__9093\ : InMux
    port map (
            O => \N__35866\,
            I => \N__35829\
        );

    \I__9092\ : InMux
    port map (
            O => \N__35865\,
            I => \N__35829\
        );

    \I__9091\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35829\
        );

    \I__9090\ : InMux
    port map (
            O => \N__35863\,
            I => \N__35829\
        );

    \I__9089\ : InMux
    port map (
            O => \N__35862\,
            I => \N__35829\
        );

    \I__9088\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35829\
        );

    \I__9087\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35829\
        );

    \I__9086\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35814\
        );

    \I__9085\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35814\
        );

    \I__9084\ : InMux
    port map (
            O => \N__35857\,
            I => \N__35814\
        );

    \I__9083\ : InMux
    port map (
            O => \N__35856\,
            I => \N__35814\
        );

    \I__9082\ : InMux
    port map (
            O => \N__35855\,
            I => \N__35814\
        );

    \I__9081\ : InMux
    port map (
            O => \N__35854\,
            I => \N__35814\
        );

    \I__9080\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35814\
        );

    \I__9079\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35806\
        );

    \I__9078\ : InMux
    port map (
            O => \N__35851\,
            I => \N__35803\
        );

    \I__9077\ : InMux
    port map (
            O => \N__35850\,
            I => \N__35800\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__35847\,
            I => \N__35797\
        );

    \I__9075\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35794\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__35829\,
            I => \N__35788\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35788\
        );

    \I__9072\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35775\
        );

    \I__9071\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35766\
        );

    \I__9070\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35766\
        );

    \I__9069\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35766\
        );

    \I__9068\ : InMux
    port map (
            O => \N__35809\,
            I => \N__35766\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__35806\,
            I => \N__35756\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__35803\,
            I => \N__35756\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__35800\,
            I => \N__35756\
        );

    \I__9064\ : Span4Mux_v
    port map (
            O => \N__35797\,
            I => \N__35750\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__35794\,
            I => \N__35750\
        );

    \I__9062\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35747\
        );

    \I__9061\ : Span4Mux_v
    port map (
            O => \N__35788\,
            I => \N__35744\
        );

    \I__9060\ : InMux
    port map (
            O => \N__35787\,
            I => \N__35741\
        );

    \I__9059\ : InMux
    port map (
            O => \N__35786\,
            I => \N__35738\
        );

    \I__9058\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35731\
        );

    \I__9057\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35731\
        );

    \I__9056\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35731\
        );

    \I__9055\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35728\
        );

    \I__9054\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35725\
        );

    \I__9053\ : InMux
    port map (
            O => \N__35780\,
            I => \N__35718\
        );

    \I__9052\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35718\
        );

    \I__9051\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35718\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__35775\,
            I => \N__35708\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__35766\,
            I => \N__35708\
        );

    \I__9048\ : InMux
    port map (
            O => \N__35765\,
            I => \N__35701\
        );

    \I__9047\ : InMux
    port map (
            O => \N__35764\,
            I => \N__35701\
        );

    \I__9046\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35701\
        );

    \I__9045\ : Span4Mux_v
    port map (
            O => \N__35756\,
            I => \N__35698\
        );

    \I__9044\ : InMux
    port map (
            O => \N__35755\,
            I => \N__35695\
        );

    \I__9043\ : Span4Mux_h
    port map (
            O => \N__35750\,
            I => \N__35692\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__35747\,
            I => \N__35689\
        );

    \I__9041\ : Sp12to4
    port map (
            O => \N__35744\,
            I => \N__35680\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__35741\,
            I => \N__35680\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__35738\,
            I => \N__35680\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__35731\,
            I => \N__35680\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__35728\,
            I => \N__35673\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__35725\,
            I => \N__35673\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__35718\,
            I => \N__35673\
        );

    \I__9034\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35666\
        );

    \I__9033\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35666\
        );

    \I__9032\ : InMux
    port map (
            O => \N__35715\,
            I => \N__35666\
        );

    \I__9031\ : InMux
    port map (
            O => \N__35714\,
            I => \N__35661\
        );

    \I__9030\ : InMux
    port map (
            O => \N__35713\,
            I => \N__35661\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__35708\,
            I => \N_458_0\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__35701\,
            I => \N_458_0\
        );

    \I__9027\ : Odrv4
    port map (
            O => \N__35698\,
            I => \N_458_0\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__35695\,
            I => \N_458_0\
        );

    \I__9025\ : Odrv4
    port map (
            O => \N__35692\,
            I => \N_458_0\
        );

    \I__9024\ : Odrv4
    port map (
            O => \N__35689\,
            I => \N_458_0\
        );

    \I__9023\ : Odrv12
    port map (
            O => \N__35680\,
            I => \N_458_0\
        );

    \I__9022\ : Odrv4
    port map (
            O => \N__35673\,
            I => \N_458_0\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__35666\,
            I => \N_458_0\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__35661\,
            I => \N_458_0\
        );

    \I__9019\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35619\
        );

    \I__9018\ : InMux
    port map (
            O => \N__35639\,
            I => \N__35619\
        );

    \I__9017\ : InMux
    port map (
            O => \N__35638\,
            I => \N__35619\
        );

    \I__9016\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35619\
        );

    \I__9015\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35619\
        );

    \I__9014\ : InMux
    port map (
            O => \N__35635\,
            I => \N__35619\
        );

    \I__9013\ : InMux
    port map (
            O => \N__35634\,
            I => \N__35619\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__35619\,
            I => \N__35606\
        );

    \I__9011\ : InMux
    port map (
            O => \N__35618\,
            I => \N__35589\
        );

    \I__9010\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35589\
        );

    \I__9009\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35589\
        );

    \I__9008\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35589\
        );

    \I__9007\ : InMux
    port map (
            O => \N__35614\,
            I => \N__35589\
        );

    \I__9006\ : InMux
    port map (
            O => \N__35613\,
            I => \N__35589\
        );

    \I__9005\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35589\
        );

    \I__9004\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35589\
        );

    \I__9003\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35586\
        );

    \I__9002\ : CascadeMux
    port map (
            O => \N__35609\,
            I => \N__35583\
        );

    \I__9001\ : Span4Mux_v
    port map (
            O => \N__35606\,
            I => \N__35580\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__35589\,
            I => \N__35573\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__35586\,
            I => \N__35573\
        );

    \I__8998\ : InMux
    port map (
            O => \N__35583\,
            I => \N__35570\
        );

    \I__8997\ : Span4Mux_h
    port map (
            O => \N__35580\,
            I => \N__35567\
        );

    \I__8996\ : InMux
    port map (
            O => \N__35579\,
            I => \N__35564\
        );

    \I__8995\ : InMux
    port map (
            O => \N__35578\,
            I => \N__35561\
        );

    \I__8994\ : Span12Mux_h
    port map (
            O => \N__35573\,
            I => \N__35558\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__35570\,
            I => \N__35555\
        );

    \I__8992\ : Span4Mux_h
    port map (
            O => \N__35567\,
            I => \N__35552\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__35564\,
            I => \N__35549\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__35561\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__8989\ : Odrv12
    port map (
            O => \N__35558\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__35555\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__8987\ : Odrv4
    port map (
            O => \N__35552\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__8986\ : Odrv4
    port map (
            O => \N__35549\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__8985\ : InMux
    port map (
            O => \N__35538\,
            I => \N__35535\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__35535\,
            I => \N__35532\
        );

    \I__8983\ : Span4Mux_h
    port map (
            O => \N__35532\,
            I => \N__35529\
        );

    \I__8982\ : Odrv4
    port map (
            O => \N__35529\,
            I => \un1_M_this_external_address_q_cry_5_THRU_CO\
        );

    \I__8981\ : IoInMux
    port map (
            O => \N__35526\,
            I => \N__35523\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__35523\,
            I => \N__35520\
        );

    \I__8979\ : IoSpan4Mux
    port map (
            O => \N__35520\,
            I => \N__35516\
        );

    \I__8978\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35512\
        );

    \I__8977\ : IoSpan4Mux
    port map (
            O => \N__35516\,
            I => \N__35509\
        );

    \I__8976\ : CascadeMux
    port map (
            O => \N__35515\,
            I => \N__35506\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__35512\,
            I => \N__35503\
        );

    \I__8974\ : Span4Mux_s3_h
    port map (
            O => \N__35509\,
            I => \N__35500\
        );

    \I__8973\ : InMux
    port map (
            O => \N__35506\,
            I => \N__35497\
        );

    \I__8972\ : Span4Mux_h
    port map (
            O => \N__35503\,
            I => \N__35494\
        );

    \I__8971\ : Odrv4
    port map (
            O => \N__35500\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__35497\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__8969\ : Odrv4
    port map (
            O => \N__35494\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__8968\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35470\
        );

    \I__8967\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35470\
        );

    \I__8966\ : InMux
    port map (
            O => \N__35485\,
            I => \N__35470\
        );

    \I__8965\ : InMux
    port map (
            O => \N__35484\,
            I => \N__35470\
        );

    \I__8964\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35463\
        );

    \I__8963\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35460\
        );

    \I__8962\ : InMux
    port map (
            O => \N__35481\,
            I => \N__35453\
        );

    \I__8961\ : InMux
    port map (
            O => \N__35480\,
            I => \N__35453\
        );

    \I__8960\ : InMux
    port map (
            O => \N__35479\,
            I => \N__35453\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__35470\,
            I => \N__35449\
        );

    \I__8958\ : CascadeMux
    port map (
            O => \N__35469\,
            I => \N__35446\
        );

    \I__8957\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35436\
        );

    \I__8956\ : CascadeMux
    port map (
            O => \N__35467\,
            I => \N__35432\
        );

    \I__8955\ : InMux
    port map (
            O => \N__35466\,
            I => \N__35424\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__35463\,
            I => \N__35415\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__35460\,
            I => \N__35410\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__35453\,
            I => \N__35410\
        );

    \I__8951\ : InMux
    port map (
            O => \N__35452\,
            I => \N__35407\
        );

    \I__8950\ : Span4Mux_h
    port map (
            O => \N__35449\,
            I => \N__35404\
        );

    \I__8949\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35401\
        );

    \I__8948\ : InMux
    port map (
            O => \N__35445\,
            I => \N__35392\
        );

    \I__8947\ : InMux
    port map (
            O => \N__35444\,
            I => \N__35392\
        );

    \I__8946\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35383\
        );

    \I__8945\ : InMux
    port map (
            O => \N__35442\,
            I => \N__35383\
        );

    \I__8944\ : InMux
    port map (
            O => \N__35441\,
            I => \N__35383\
        );

    \I__8943\ : InMux
    port map (
            O => \N__35440\,
            I => \N__35383\
        );

    \I__8942\ : InMux
    port map (
            O => \N__35439\,
            I => \N__35380\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__35436\,
            I => \N__35377\
        );

    \I__8940\ : InMux
    port map (
            O => \N__35435\,
            I => \N__35372\
        );

    \I__8939\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35372\
        );

    \I__8938\ : InMux
    port map (
            O => \N__35431\,
            I => \N__35369\
        );

    \I__8937\ : InMux
    port map (
            O => \N__35430\,
            I => \N__35366\
        );

    \I__8936\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35359\
        );

    \I__8935\ : InMux
    port map (
            O => \N__35428\,
            I => \N__35359\
        );

    \I__8934\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35359\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__35424\,
            I => \N__35356\
        );

    \I__8932\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35345\
        );

    \I__8931\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35345\
        );

    \I__8930\ : InMux
    port map (
            O => \N__35421\,
            I => \N__35345\
        );

    \I__8929\ : InMux
    port map (
            O => \N__35420\,
            I => \N__35345\
        );

    \I__8928\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35345\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__35418\,
            I => \N__35342\
        );

    \I__8926\ : Span4Mux_h
    port map (
            O => \N__35415\,
            I => \N__35337\
        );

    \I__8925\ : Span4Mux_h
    port map (
            O => \N__35410\,
            I => \N__35334\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__35407\,
            I => \N__35327\
        );

    \I__8923\ : Span4Mux_v
    port map (
            O => \N__35404\,
            I => \N__35327\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__35401\,
            I => \N__35327\
        );

    \I__8921\ : InMux
    port map (
            O => \N__35400\,
            I => \N__35324\
        );

    \I__8920\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35321\
        );

    \I__8919\ : InMux
    port map (
            O => \N__35398\,
            I => \N__35316\
        );

    \I__8918\ : InMux
    port map (
            O => \N__35397\,
            I => \N__35316\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__35392\,
            I => \N__35313\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__35383\,
            I => \N__35306\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__35380\,
            I => \N__35306\
        );

    \I__8914\ : Span4Mux_v
    port map (
            O => \N__35377\,
            I => \N__35306\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__35372\,
            I => \N__35303\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__35369\,
            I => \N__35292\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__35366\,
            I => \N__35292\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__35359\,
            I => \N__35292\
        );

    \I__8909\ : Span4Mux_v
    port map (
            O => \N__35356\,
            I => \N__35292\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__35345\,
            I => \N__35292\
        );

    \I__8907\ : InMux
    port map (
            O => \N__35342\,
            I => \N__35289\
        );

    \I__8906\ : InMux
    port map (
            O => \N__35341\,
            I => \N__35284\
        );

    \I__8905\ : InMux
    port map (
            O => \N__35340\,
            I => \N__35284\
        );

    \I__8904\ : Span4Mux_h
    port map (
            O => \N__35337\,
            I => \N__35279\
        );

    \I__8903\ : Span4Mux_h
    port map (
            O => \N__35334\,
            I => \N__35279\
        );

    \I__8902\ : Span4Mux_h
    port map (
            O => \N__35327\,
            I => \N__35274\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__35324\,
            I => \N__35274\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__35321\,
            I => \N__35261\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__35316\,
            I => \N__35261\
        );

    \I__8898\ : Span4Mux_v
    port map (
            O => \N__35313\,
            I => \N__35261\
        );

    \I__8897\ : Span4Mux_h
    port map (
            O => \N__35306\,
            I => \N__35261\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__35303\,
            I => \N__35261\
        );

    \I__8895\ : Span4Mux_v
    port map (
            O => \N__35292\,
            I => \N__35261\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__35289\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__35284\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__8892\ : Odrv4
    port map (
            O => \N__35279\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__8891\ : Odrv4
    port map (
            O => \N__35274\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__8890\ : Odrv4
    port map (
            O => \N__35261\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__8889\ : CascadeMux
    port map (
            O => \N__35250\,
            I => \N__35243\
        );

    \I__8888\ : CascadeMux
    port map (
            O => \N__35249\,
            I => \N__35240\
        );

    \I__8887\ : CascadeMux
    port map (
            O => \N__35248\,
            I => \N__35225\
        );

    \I__8886\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35222\
        );

    \I__8885\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35213\
        );

    \I__8884\ : InMux
    port map (
            O => \N__35243\,
            I => \N__35213\
        );

    \I__8883\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35213\
        );

    \I__8882\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35213\
        );

    \I__8881\ : InMux
    port map (
            O => \N__35238\,
            I => \N__35210\
        );

    \I__8880\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35201\
        );

    \I__8879\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35201\
        );

    \I__8878\ : InMux
    port map (
            O => \N__35235\,
            I => \N__35201\
        );

    \I__8877\ : InMux
    port map (
            O => \N__35234\,
            I => \N__35201\
        );

    \I__8876\ : CascadeMux
    port map (
            O => \N__35233\,
            I => \N__35197\
        );

    \I__8875\ : CascadeMux
    port map (
            O => \N__35232\,
            I => \N__35194\
        );

    \I__8874\ : CascadeMux
    port map (
            O => \N__35231\,
            I => \N__35191\
        );

    \I__8873\ : InMux
    port map (
            O => \N__35230\,
            I => \N__35180\
        );

    \I__8872\ : CascadeMux
    port map (
            O => \N__35229\,
            I => \N__35177\
        );

    \I__8871\ : CascadeMux
    port map (
            O => \N__35228\,
            I => \N__35171\
        );

    \I__8870\ : InMux
    port map (
            O => \N__35225\,
            I => \N__35166\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__35222\,
            I => \N__35159\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__35213\,
            I => \N__35159\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__35210\,
            I => \N__35156\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__35201\,
            I => \N__35153\
        );

    \I__8865\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35142\
        );

    \I__8864\ : InMux
    port map (
            O => \N__35197\,
            I => \N__35142\
        );

    \I__8863\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35142\
        );

    \I__8862\ : InMux
    port map (
            O => \N__35191\,
            I => \N__35142\
        );

    \I__8861\ : InMux
    port map (
            O => \N__35190\,
            I => \N__35142\
        );

    \I__8860\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35139\
        );

    \I__8859\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35136\
        );

    \I__8858\ : InMux
    port map (
            O => \N__35187\,
            I => \N__35129\
        );

    \I__8857\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35129\
        );

    \I__8856\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35129\
        );

    \I__8855\ : InMux
    port map (
            O => \N__35184\,
            I => \N__35126\
        );

    \I__8854\ : CascadeMux
    port map (
            O => \N__35183\,
            I => \N__35123\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__35180\,
            I => \N__35116\
        );

    \I__8852\ : InMux
    port map (
            O => \N__35177\,
            I => \N__35111\
        );

    \I__8851\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35111\
        );

    \I__8850\ : InMux
    port map (
            O => \N__35175\,
            I => \N__35106\
        );

    \I__8849\ : InMux
    port map (
            O => \N__35174\,
            I => \N__35106\
        );

    \I__8848\ : InMux
    port map (
            O => \N__35171\,
            I => \N__35099\
        );

    \I__8847\ : InMux
    port map (
            O => \N__35170\,
            I => \N__35099\
        );

    \I__8846\ : InMux
    port map (
            O => \N__35169\,
            I => \N__35099\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__35166\,
            I => \N__35095\
        );

    \I__8844\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35090\
        );

    \I__8843\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35090\
        );

    \I__8842\ : Span4Mux_v
    port map (
            O => \N__35159\,
            I => \N__35081\
        );

    \I__8841\ : Span4Mux_h
    port map (
            O => \N__35156\,
            I => \N__35081\
        );

    \I__8840\ : Span4Mux_v
    port map (
            O => \N__35153\,
            I => \N__35081\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__35142\,
            I => \N__35081\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__35139\,
            I => \N__35071\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__35136\,
            I => \N__35071\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__35129\,
            I => \N__35071\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__35126\,
            I => \N__35071\
        );

    \I__8834\ : InMux
    port map (
            O => \N__35123\,
            I => \N__35064\
        );

    \I__8833\ : InMux
    port map (
            O => \N__35122\,
            I => \N__35064\
        );

    \I__8832\ : InMux
    port map (
            O => \N__35121\,
            I => \N__35064\
        );

    \I__8831\ : InMux
    port map (
            O => \N__35120\,
            I => \N__35061\
        );

    \I__8830\ : InMux
    port map (
            O => \N__35119\,
            I => \N__35058\
        );

    \I__8829\ : Span4Mux_v
    port map (
            O => \N__35116\,
            I => \N__35049\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__35111\,
            I => \N__35049\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__35106\,
            I => \N__35049\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__35099\,
            I => \N__35049\
        );

    \I__8825\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35046\
        );

    \I__8824\ : Span4Mux_h
    port map (
            O => \N__35095\,
            I => \N__35043\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__35090\,
            I => \N__35038\
        );

    \I__8822\ : Span4Mux_h
    port map (
            O => \N__35081\,
            I => \N__35038\
        );

    \I__8821\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35035\
        );

    \I__8820\ : Span12Mux_h
    port map (
            O => \N__35071\,
            I => \N__35032\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__35064\,
            I => \N__35027\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__35061\,
            I => \N__35027\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__35058\,
            I => \N__35020\
        );

    \I__8816\ : Span4Mux_v
    port map (
            O => \N__35049\,
            I => \N__35020\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__35046\,
            I => \N__35020\
        );

    \I__8814\ : Span4Mux_h
    port map (
            O => \N__35043\,
            I => \N__35015\
        );

    \I__8813\ : Span4Mux_h
    port map (
            O => \N__35038\,
            I => \N__35015\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__35035\,
            I => \N_156_0\
        );

    \I__8811\ : Odrv12
    port map (
            O => \N__35032\,
            I => \N_156_0\
        );

    \I__8810\ : Odrv12
    port map (
            O => \N__35027\,
            I => \N_156_0\
        );

    \I__8809\ : Odrv4
    port map (
            O => \N__35020\,
            I => \N_156_0\
        );

    \I__8808\ : Odrv4
    port map (
            O => \N__35015\,
            I => \N_156_0\
        );

    \I__8807\ : CascadeMux
    port map (
            O => \N__35004\,
            I => \N__34991\
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__35003\,
            I => \N__34983\
        );

    \I__8805\ : InMux
    port map (
            O => \N__35002\,
            I => \N__34975\
        );

    \I__8804\ : InMux
    port map (
            O => \N__35001\,
            I => \N__34966\
        );

    \I__8803\ : InMux
    port map (
            O => \N__35000\,
            I => \N__34966\
        );

    \I__8802\ : InMux
    port map (
            O => \N__34999\,
            I => \N__34966\
        );

    \I__8801\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34966\
        );

    \I__8800\ : InMux
    port map (
            O => \N__34997\,
            I => \N__34963\
        );

    \I__8799\ : CascadeMux
    port map (
            O => \N__34996\,
            I => \N__34959\
        );

    \I__8798\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34954\
        );

    \I__8797\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34954\
        );

    \I__8796\ : InMux
    port map (
            O => \N__34991\,
            I => \N__34947\
        );

    \I__8795\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34940\
        );

    \I__8794\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34940\
        );

    \I__8793\ : InMux
    port map (
            O => \N__34988\,
            I => \N__34940\
        );

    \I__8792\ : InMux
    port map (
            O => \N__34987\,
            I => \N__34930\
        );

    \I__8791\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34930\
        );

    \I__8790\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34927\
        );

    \I__8789\ : InMux
    port map (
            O => \N__34982\,
            I => \N__34924\
        );

    \I__8788\ : InMux
    port map (
            O => \N__34981\,
            I => \N__34911\
        );

    \I__8787\ : InMux
    port map (
            O => \N__34980\,
            I => \N__34911\
        );

    \I__8786\ : InMux
    port map (
            O => \N__34979\,
            I => \N__34911\
        );

    \I__8785\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34911\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__34975\,
            I => \N__34908\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__34966\,
            I => \N__34903\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__34963\,
            I => \N__34903\
        );

    \I__8781\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34900\
        );

    \I__8780\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34897\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__34954\,
            I => \N__34894\
        );

    \I__8778\ : InMux
    port map (
            O => \N__34953\,
            I => \N__34882\
        );

    \I__8777\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34882\
        );

    \I__8776\ : InMux
    port map (
            O => \N__34951\,
            I => \N__34882\
        );

    \I__8775\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34879\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__34947\,
            I => \N__34874\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__34940\,
            I => \N__34874\
        );

    \I__8772\ : InMux
    port map (
            O => \N__34939\,
            I => \N__34867\
        );

    \I__8771\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34867\
        );

    \I__8770\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34867\
        );

    \I__8769\ : InMux
    port map (
            O => \N__34936\,
            I => \N__34862\
        );

    \I__8768\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34862\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__34930\,
            I => \N__34857\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__34927\,
            I => \N__34857\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__34924\,
            I => \N__34854\
        );

    \I__8764\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34851\
        );

    \I__8763\ : InMux
    port map (
            O => \N__34922\,
            I => \N__34848\
        );

    \I__8762\ : InMux
    port map (
            O => \N__34921\,
            I => \N__34843\
        );

    \I__8761\ : InMux
    port map (
            O => \N__34920\,
            I => \N__34843\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__34911\,
            I => \N__34836\
        );

    \I__8759\ : Span4Mux_v
    port map (
            O => \N__34908\,
            I => \N__34836\
        );

    \I__8758\ : Span4Mux_v
    port map (
            O => \N__34903\,
            I => \N__34836\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__34900\,
            I => \N__34833\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__34897\,
            I => \N__34828\
        );

    \I__8755\ : Span4Mux_v
    port map (
            O => \N__34894\,
            I => \N__34828\
        );

    \I__8754\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34817\
        );

    \I__8753\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34817\
        );

    \I__8752\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34817\
        );

    \I__8751\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34817\
        );

    \I__8750\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34817\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__34882\,
            I => \N__34814\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__34879\,
            I => \N__34803\
        );

    \I__8747\ : Span4Mux_h
    port map (
            O => \N__34874\,
            I => \N__34803\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__34867\,
            I => \N__34803\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__34862\,
            I => \N__34803\
        );

    \I__8744\ : Span4Mux_h
    port map (
            O => \N__34857\,
            I => \N__34803\
        );

    \I__8743\ : Odrv12
    port map (
            O => \N__34854\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__34851\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__34848\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__34843\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8739\ : Odrv4
    port map (
            O => \N__34836\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8738\ : Odrv4
    port map (
            O => \N__34833\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__34828\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__34817\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8735\ : Odrv4
    port map (
            O => \N__34814\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8734\ : Odrv4
    port map (
            O => \N__34803\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8733\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34779\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__34779\,
            I => \N__34776\
        );

    \I__8731\ : Span4Mux_v
    port map (
            O => \N__34776\,
            I => \N__34773\
        );

    \I__8730\ : Odrv4
    port map (
            O => \N__34773\,
            I => \N_69_0\
        );

    \I__8729\ : CascadeMux
    port map (
            O => \N__34770\,
            I => \N__34767\
        );

    \I__8728\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34763\
        );

    \I__8727\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34758\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__34763\,
            I => \N__34754\
        );

    \I__8725\ : CascadeMux
    port map (
            O => \N__34762\,
            I => \N__34751\
        );

    \I__8724\ : CascadeMux
    port map (
            O => \N__34761\,
            I => \N__34747\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__34758\,
            I => \N__34744\
        );

    \I__8722\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34741\
        );

    \I__8721\ : Span4Mux_v
    port map (
            O => \N__34754\,
            I => \N__34736\
        );

    \I__8720\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34733\
        );

    \I__8719\ : InMux
    port map (
            O => \N__34750\,
            I => \N__34730\
        );

    \I__8718\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34727\
        );

    \I__8717\ : Span4Mux_h
    port map (
            O => \N__34744\,
            I => \N__34722\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__34741\,
            I => \N__34722\
        );

    \I__8715\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34719\
        );

    \I__8714\ : CascadeMux
    port map (
            O => \N__34739\,
            I => \N__34716\
        );

    \I__8713\ : Span4Mux_h
    port map (
            O => \N__34736\,
            I => \N__34707\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__34733\,
            I => \N__34707\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__34730\,
            I => \N__34707\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__34727\,
            I => \N__34707\
        );

    \I__8709\ : Span4Mux_v
    port map (
            O => \N__34722\,
            I => \N__34702\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__34719\,
            I => \N__34699\
        );

    \I__8707\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34696\
        );

    \I__8706\ : Span4Mux_v
    port map (
            O => \N__34707\,
            I => \N__34691\
        );

    \I__8705\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34688\
        );

    \I__8704\ : CascadeMux
    port map (
            O => \N__34705\,
            I => \N__34685\
        );

    \I__8703\ : Span4Mux_h
    port map (
            O => \N__34702\,
            I => \N__34679\
        );

    \I__8702\ : Span4Mux_v
    port map (
            O => \N__34699\,
            I => \N__34679\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__34696\,
            I => \N__34676\
        );

    \I__8700\ : InMux
    port map (
            O => \N__34695\,
            I => \N__34673\
        );

    \I__8699\ : CascadeMux
    port map (
            O => \N__34694\,
            I => \N__34670\
        );

    \I__8698\ : Span4Mux_h
    port map (
            O => \N__34691\,
            I => \N__34665\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__34688\,
            I => \N__34665\
        );

    \I__8696\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34659\
        );

    \I__8695\ : InMux
    port map (
            O => \N__34684\,
            I => \N__34659\
        );

    \I__8694\ : Span4Mux_h
    port map (
            O => \N__34679\,
            I => \N__34652\
        );

    \I__8693\ : Span4Mux_v
    port map (
            O => \N__34676\,
            I => \N__34652\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__34673\,
            I => \N__34652\
        );

    \I__8691\ : InMux
    port map (
            O => \N__34670\,
            I => \N__34649\
        );

    \I__8690\ : Span4Mux_v
    port map (
            O => \N__34665\,
            I => \N__34646\
        );

    \I__8689\ : InMux
    port map (
            O => \N__34664\,
            I => \N__34643\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__34659\,
            I => \N__34640\
        );

    \I__8687\ : Span4Mux_h
    port map (
            O => \N__34652\,
            I => \N__34635\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__34649\,
            I => \N__34635\
        );

    \I__8685\ : Span4Mux_h
    port map (
            O => \N__34646\,
            I => \N__34630\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__34643\,
            I => \N__34630\
        );

    \I__8683\ : Span12Mux_v
    port map (
            O => \N__34640\,
            I => \N__34627\
        );

    \I__8682\ : Span4Mux_h
    port map (
            O => \N__34635\,
            I => \N__34624\
        );

    \I__8681\ : Span4Mux_v
    port map (
            O => \N__34630\,
            I => \N__34621\
        );

    \I__8680\ : Span12Mux_h
    port map (
            O => \N__34627\,
            I => \N__34618\
        );

    \I__8679\ : IoSpan4Mux
    port map (
            O => \N__34624\,
            I => \N__34615\
        );

    \I__8678\ : Span4Mux_h
    port map (
            O => \N__34621\,
            I => \N__34612\
        );

    \I__8677\ : Odrv12
    port map (
            O => \N__34618\,
            I => port_data_c_5
        );

    \I__8676\ : Odrv4
    port map (
            O => \N__34615\,
            I => port_data_c_5
        );

    \I__8675\ : Odrv4
    port map (
            O => \N__34612\,
            I => port_data_c_5
        );

    \I__8674\ : CascadeMux
    port map (
            O => \N__34605\,
            I => \N__34602\
        );

    \I__8673\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34599\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__34599\,
            I => \M_this_data_tmp_qZ0Z_5\
        );

    \I__8671\ : ClkMux
    port map (
            O => \N__34596\,
            I => \N__34206\
        );

    \I__8670\ : ClkMux
    port map (
            O => \N__34595\,
            I => \N__34206\
        );

    \I__8669\ : ClkMux
    port map (
            O => \N__34594\,
            I => \N__34206\
        );

    \I__8668\ : ClkMux
    port map (
            O => \N__34593\,
            I => \N__34206\
        );

    \I__8667\ : ClkMux
    port map (
            O => \N__34592\,
            I => \N__34206\
        );

    \I__8666\ : ClkMux
    port map (
            O => \N__34591\,
            I => \N__34206\
        );

    \I__8665\ : ClkMux
    port map (
            O => \N__34590\,
            I => \N__34206\
        );

    \I__8664\ : ClkMux
    port map (
            O => \N__34589\,
            I => \N__34206\
        );

    \I__8663\ : ClkMux
    port map (
            O => \N__34588\,
            I => \N__34206\
        );

    \I__8662\ : ClkMux
    port map (
            O => \N__34587\,
            I => \N__34206\
        );

    \I__8661\ : ClkMux
    port map (
            O => \N__34586\,
            I => \N__34206\
        );

    \I__8660\ : ClkMux
    port map (
            O => \N__34585\,
            I => \N__34206\
        );

    \I__8659\ : ClkMux
    port map (
            O => \N__34584\,
            I => \N__34206\
        );

    \I__8658\ : ClkMux
    port map (
            O => \N__34583\,
            I => \N__34206\
        );

    \I__8657\ : ClkMux
    port map (
            O => \N__34582\,
            I => \N__34206\
        );

    \I__8656\ : ClkMux
    port map (
            O => \N__34581\,
            I => \N__34206\
        );

    \I__8655\ : ClkMux
    port map (
            O => \N__34580\,
            I => \N__34206\
        );

    \I__8654\ : ClkMux
    port map (
            O => \N__34579\,
            I => \N__34206\
        );

    \I__8653\ : ClkMux
    port map (
            O => \N__34578\,
            I => \N__34206\
        );

    \I__8652\ : ClkMux
    port map (
            O => \N__34577\,
            I => \N__34206\
        );

    \I__8651\ : ClkMux
    port map (
            O => \N__34576\,
            I => \N__34206\
        );

    \I__8650\ : ClkMux
    port map (
            O => \N__34575\,
            I => \N__34206\
        );

    \I__8649\ : ClkMux
    port map (
            O => \N__34574\,
            I => \N__34206\
        );

    \I__8648\ : ClkMux
    port map (
            O => \N__34573\,
            I => \N__34206\
        );

    \I__8647\ : ClkMux
    port map (
            O => \N__34572\,
            I => \N__34206\
        );

    \I__8646\ : ClkMux
    port map (
            O => \N__34571\,
            I => \N__34206\
        );

    \I__8645\ : ClkMux
    port map (
            O => \N__34570\,
            I => \N__34206\
        );

    \I__8644\ : ClkMux
    port map (
            O => \N__34569\,
            I => \N__34206\
        );

    \I__8643\ : ClkMux
    port map (
            O => \N__34568\,
            I => \N__34206\
        );

    \I__8642\ : ClkMux
    port map (
            O => \N__34567\,
            I => \N__34206\
        );

    \I__8641\ : ClkMux
    port map (
            O => \N__34566\,
            I => \N__34206\
        );

    \I__8640\ : ClkMux
    port map (
            O => \N__34565\,
            I => \N__34206\
        );

    \I__8639\ : ClkMux
    port map (
            O => \N__34564\,
            I => \N__34206\
        );

    \I__8638\ : ClkMux
    port map (
            O => \N__34563\,
            I => \N__34206\
        );

    \I__8637\ : ClkMux
    port map (
            O => \N__34562\,
            I => \N__34206\
        );

    \I__8636\ : ClkMux
    port map (
            O => \N__34561\,
            I => \N__34206\
        );

    \I__8635\ : ClkMux
    port map (
            O => \N__34560\,
            I => \N__34206\
        );

    \I__8634\ : ClkMux
    port map (
            O => \N__34559\,
            I => \N__34206\
        );

    \I__8633\ : ClkMux
    port map (
            O => \N__34558\,
            I => \N__34206\
        );

    \I__8632\ : ClkMux
    port map (
            O => \N__34557\,
            I => \N__34206\
        );

    \I__8631\ : ClkMux
    port map (
            O => \N__34556\,
            I => \N__34206\
        );

    \I__8630\ : ClkMux
    port map (
            O => \N__34555\,
            I => \N__34206\
        );

    \I__8629\ : ClkMux
    port map (
            O => \N__34554\,
            I => \N__34206\
        );

    \I__8628\ : ClkMux
    port map (
            O => \N__34553\,
            I => \N__34206\
        );

    \I__8627\ : ClkMux
    port map (
            O => \N__34552\,
            I => \N__34206\
        );

    \I__8626\ : ClkMux
    port map (
            O => \N__34551\,
            I => \N__34206\
        );

    \I__8625\ : ClkMux
    port map (
            O => \N__34550\,
            I => \N__34206\
        );

    \I__8624\ : ClkMux
    port map (
            O => \N__34549\,
            I => \N__34206\
        );

    \I__8623\ : ClkMux
    port map (
            O => \N__34548\,
            I => \N__34206\
        );

    \I__8622\ : ClkMux
    port map (
            O => \N__34547\,
            I => \N__34206\
        );

    \I__8621\ : ClkMux
    port map (
            O => \N__34546\,
            I => \N__34206\
        );

    \I__8620\ : ClkMux
    port map (
            O => \N__34545\,
            I => \N__34206\
        );

    \I__8619\ : ClkMux
    port map (
            O => \N__34544\,
            I => \N__34206\
        );

    \I__8618\ : ClkMux
    port map (
            O => \N__34543\,
            I => \N__34206\
        );

    \I__8617\ : ClkMux
    port map (
            O => \N__34542\,
            I => \N__34206\
        );

    \I__8616\ : ClkMux
    port map (
            O => \N__34541\,
            I => \N__34206\
        );

    \I__8615\ : ClkMux
    port map (
            O => \N__34540\,
            I => \N__34206\
        );

    \I__8614\ : ClkMux
    port map (
            O => \N__34539\,
            I => \N__34206\
        );

    \I__8613\ : ClkMux
    port map (
            O => \N__34538\,
            I => \N__34206\
        );

    \I__8612\ : ClkMux
    port map (
            O => \N__34537\,
            I => \N__34206\
        );

    \I__8611\ : ClkMux
    port map (
            O => \N__34536\,
            I => \N__34206\
        );

    \I__8610\ : ClkMux
    port map (
            O => \N__34535\,
            I => \N__34206\
        );

    \I__8609\ : ClkMux
    port map (
            O => \N__34534\,
            I => \N__34206\
        );

    \I__8608\ : ClkMux
    port map (
            O => \N__34533\,
            I => \N__34206\
        );

    \I__8607\ : ClkMux
    port map (
            O => \N__34532\,
            I => \N__34206\
        );

    \I__8606\ : ClkMux
    port map (
            O => \N__34531\,
            I => \N__34206\
        );

    \I__8605\ : ClkMux
    port map (
            O => \N__34530\,
            I => \N__34206\
        );

    \I__8604\ : ClkMux
    port map (
            O => \N__34529\,
            I => \N__34206\
        );

    \I__8603\ : ClkMux
    port map (
            O => \N__34528\,
            I => \N__34206\
        );

    \I__8602\ : ClkMux
    port map (
            O => \N__34527\,
            I => \N__34206\
        );

    \I__8601\ : ClkMux
    port map (
            O => \N__34526\,
            I => \N__34206\
        );

    \I__8600\ : ClkMux
    port map (
            O => \N__34525\,
            I => \N__34206\
        );

    \I__8599\ : ClkMux
    port map (
            O => \N__34524\,
            I => \N__34206\
        );

    \I__8598\ : ClkMux
    port map (
            O => \N__34523\,
            I => \N__34206\
        );

    \I__8597\ : ClkMux
    port map (
            O => \N__34522\,
            I => \N__34206\
        );

    \I__8596\ : ClkMux
    port map (
            O => \N__34521\,
            I => \N__34206\
        );

    \I__8595\ : ClkMux
    port map (
            O => \N__34520\,
            I => \N__34206\
        );

    \I__8594\ : ClkMux
    port map (
            O => \N__34519\,
            I => \N__34206\
        );

    \I__8593\ : ClkMux
    port map (
            O => \N__34518\,
            I => \N__34206\
        );

    \I__8592\ : ClkMux
    port map (
            O => \N__34517\,
            I => \N__34206\
        );

    \I__8591\ : ClkMux
    port map (
            O => \N__34516\,
            I => \N__34206\
        );

    \I__8590\ : ClkMux
    port map (
            O => \N__34515\,
            I => \N__34206\
        );

    \I__8589\ : ClkMux
    port map (
            O => \N__34514\,
            I => \N__34206\
        );

    \I__8588\ : ClkMux
    port map (
            O => \N__34513\,
            I => \N__34206\
        );

    \I__8587\ : ClkMux
    port map (
            O => \N__34512\,
            I => \N__34206\
        );

    \I__8586\ : ClkMux
    port map (
            O => \N__34511\,
            I => \N__34206\
        );

    \I__8585\ : ClkMux
    port map (
            O => \N__34510\,
            I => \N__34206\
        );

    \I__8584\ : ClkMux
    port map (
            O => \N__34509\,
            I => \N__34206\
        );

    \I__8583\ : ClkMux
    port map (
            O => \N__34508\,
            I => \N__34206\
        );

    \I__8582\ : ClkMux
    port map (
            O => \N__34507\,
            I => \N__34206\
        );

    \I__8581\ : ClkMux
    port map (
            O => \N__34506\,
            I => \N__34206\
        );

    \I__8580\ : ClkMux
    port map (
            O => \N__34505\,
            I => \N__34206\
        );

    \I__8579\ : ClkMux
    port map (
            O => \N__34504\,
            I => \N__34206\
        );

    \I__8578\ : ClkMux
    port map (
            O => \N__34503\,
            I => \N__34206\
        );

    \I__8577\ : ClkMux
    port map (
            O => \N__34502\,
            I => \N__34206\
        );

    \I__8576\ : ClkMux
    port map (
            O => \N__34501\,
            I => \N__34206\
        );

    \I__8575\ : ClkMux
    port map (
            O => \N__34500\,
            I => \N__34206\
        );

    \I__8574\ : ClkMux
    port map (
            O => \N__34499\,
            I => \N__34206\
        );

    \I__8573\ : ClkMux
    port map (
            O => \N__34498\,
            I => \N__34206\
        );

    \I__8572\ : ClkMux
    port map (
            O => \N__34497\,
            I => \N__34206\
        );

    \I__8571\ : ClkMux
    port map (
            O => \N__34496\,
            I => \N__34206\
        );

    \I__8570\ : ClkMux
    port map (
            O => \N__34495\,
            I => \N__34206\
        );

    \I__8569\ : ClkMux
    port map (
            O => \N__34494\,
            I => \N__34206\
        );

    \I__8568\ : ClkMux
    port map (
            O => \N__34493\,
            I => \N__34206\
        );

    \I__8567\ : ClkMux
    port map (
            O => \N__34492\,
            I => \N__34206\
        );

    \I__8566\ : ClkMux
    port map (
            O => \N__34491\,
            I => \N__34206\
        );

    \I__8565\ : ClkMux
    port map (
            O => \N__34490\,
            I => \N__34206\
        );

    \I__8564\ : ClkMux
    port map (
            O => \N__34489\,
            I => \N__34206\
        );

    \I__8563\ : ClkMux
    port map (
            O => \N__34488\,
            I => \N__34206\
        );

    \I__8562\ : ClkMux
    port map (
            O => \N__34487\,
            I => \N__34206\
        );

    \I__8561\ : ClkMux
    port map (
            O => \N__34486\,
            I => \N__34206\
        );

    \I__8560\ : ClkMux
    port map (
            O => \N__34485\,
            I => \N__34206\
        );

    \I__8559\ : ClkMux
    port map (
            O => \N__34484\,
            I => \N__34206\
        );

    \I__8558\ : ClkMux
    port map (
            O => \N__34483\,
            I => \N__34206\
        );

    \I__8557\ : ClkMux
    port map (
            O => \N__34482\,
            I => \N__34206\
        );

    \I__8556\ : ClkMux
    port map (
            O => \N__34481\,
            I => \N__34206\
        );

    \I__8555\ : ClkMux
    port map (
            O => \N__34480\,
            I => \N__34206\
        );

    \I__8554\ : ClkMux
    port map (
            O => \N__34479\,
            I => \N__34206\
        );

    \I__8553\ : ClkMux
    port map (
            O => \N__34478\,
            I => \N__34206\
        );

    \I__8552\ : ClkMux
    port map (
            O => \N__34477\,
            I => \N__34206\
        );

    \I__8551\ : ClkMux
    port map (
            O => \N__34476\,
            I => \N__34206\
        );

    \I__8550\ : ClkMux
    port map (
            O => \N__34475\,
            I => \N__34206\
        );

    \I__8549\ : ClkMux
    port map (
            O => \N__34474\,
            I => \N__34206\
        );

    \I__8548\ : ClkMux
    port map (
            O => \N__34473\,
            I => \N__34206\
        );

    \I__8547\ : ClkMux
    port map (
            O => \N__34472\,
            I => \N__34206\
        );

    \I__8546\ : ClkMux
    port map (
            O => \N__34471\,
            I => \N__34206\
        );

    \I__8545\ : ClkMux
    port map (
            O => \N__34470\,
            I => \N__34206\
        );

    \I__8544\ : ClkMux
    port map (
            O => \N__34469\,
            I => \N__34206\
        );

    \I__8543\ : ClkMux
    port map (
            O => \N__34468\,
            I => \N__34206\
        );

    \I__8542\ : ClkMux
    port map (
            O => \N__34467\,
            I => \N__34206\
        );

    \I__8541\ : GlobalMux
    port map (
            O => \N__34206\,
            I => \N__34203\
        );

    \I__8540\ : gio2CtrlBuf
    port map (
            O => \N__34203\,
            I => clk_0_c_g
        );

    \I__8539\ : CEMux
    port map (
            O => \N__34200\,
            I => \N__34195\
        );

    \I__8538\ : CEMux
    port map (
            O => \N__34199\,
            I => \N__34192\
        );

    \I__8537\ : CEMux
    port map (
            O => \N__34198\,
            I => \N__34189\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__34195\,
            I => \N__34184\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__34192\,
            I => \N__34179\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__34189\,
            I => \N__34179\
        );

    \I__8533\ : CEMux
    port map (
            O => \N__34188\,
            I => \N__34176\
        );

    \I__8532\ : CEMux
    port map (
            O => \N__34187\,
            I => \N__34173\
        );

    \I__8531\ : Span4Mux_v
    port map (
            O => \N__34184\,
            I => \N__34170\
        );

    \I__8530\ : Span4Mux_v
    port map (
            O => \N__34179\,
            I => \N__34167\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__34176\,
            I => \N__34164\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__34173\,
            I => \N__34159\
        );

    \I__8527\ : Span4Mux_h
    port map (
            O => \N__34170\,
            I => \N__34152\
        );

    \I__8526\ : Span4Mux_v
    port map (
            O => \N__34167\,
            I => \N__34152\
        );

    \I__8525\ : Span4Mux_h
    port map (
            O => \N__34164\,
            I => \N__34152\
        );

    \I__8524\ : CEMux
    port map (
            O => \N__34163\,
            I => \N__34149\
        );

    \I__8523\ : CEMux
    port map (
            O => \N__34162\,
            I => \N__34146\
        );

    \I__8522\ : Span4Mux_v
    port map (
            O => \N__34159\,
            I => \N__34143\
        );

    \I__8521\ : Span4Mux_h
    port map (
            O => \N__34152\,
            I => \N__34138\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__34149\,
            I => \N__34138\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__34146\,
            I => \N__34135\
        );

    \I__8518\ : Span4Mux_h
    port map (
            O => \N__34143\,
            I => \N__34130\
        );

    \I__8517\ : Span4Mux_h
    port map (
            O => \N__34138\,
            I => \N__34130\
        );

    \I__8516\ : Odrv12
    port map (
            O => \N__34135\,
            I => \N_1142_0\
        );

    \I__8515\ : Odrv4
    port map (
            O => \N__34130\,
            I => \N_1142_0\
        );

    \I__8514\ : InMux
    port map (
            O => \N__34125\,
            I => \N__34101\
        );

    \I__8513\ : InMux
    port map (
            O => \N__34124\,
            I => \N__34098\
        );

    \I__8512\ : InMux
    port map (
            O => \N__34123\,
            I => \N__34095\
        );

    \I__8511\ : InMux
    port map (
            O => \N__34122\,
            I => \N__34092\
        );

    \I__8510\ : InMux
    port map (
            O => \N__34121\,
            I => \N__34085\
        );

    \I__8509\ : InMux
    port map (
            O => \N__34120\,
            I => \N__34085\
        );

    \I__8508\ : InMux
    port map (
            O => \N__34119\,
            I => \N__34085\
        );

    \I__8507\ : InMux
    port map (
            O => \N__34118\,
            I => \N__34082\
        );

    \I__8506\ : InMux
    port map (
            O => \N__34117\,
            I => \N__34079\
        );

    \I__8505\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34076\
        );

    \I__8504\ : InMux
    port map (
            O => \N__34115\,
            I => \N__34073\
        );

    \I__8503\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34070\
        );

    \I__8502\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34067\
        );

    \I__8501\ : InMux
    port map (
            O => \N__34112\,
            I => \N__34064\
        );

    \I__8500\ : InMux
    port map (
            O => \N__34111\,
            I => \N__34061\
        );

    \I__8499\ : InMux
    port map (
            O => \N__34110\,
            I => \N__34058\
        );

    \I__8498\ : InMux
    port map (
            O => \N__34109\,
            I => \N__34055\
        );

    \I__8497\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34052\
        );

    \I__8496\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34049\
        );

    \I__8495\ : InMux
    port map (
            O => \N__34106\,
            I => \N__34046\
        );

    \I__8494\ : InMux
    port map (
            O => \N__34105\,
            I => \N__34041\
        );

    \I__8493\ : InMux
    port map (
            O => \N__34104\,
            I => \N__34041\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__34101\,
            I => \N__34007\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__34098\,
            I => \N__34004\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__34095\,
            I => \N__34001\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__34092\,
            I => \N__33998\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__34085\,
            I => \N__33995\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__34082\,
            I => \N__33992\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__34079\,
            I => \N__33989\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__34076\,
            I => \N__33986\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__34073\,
            I => \N__33983\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__34070\,
            I => \N__33980\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__34067\,
            I => \N__33977\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__34064\,
            I => \N__33974\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__34061\,
            I => \N__33971\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__34058\,
            I => \N__33968\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__34055\,
            I => \N__33965\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__34052\,
            I => \N__33962\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__34049\,
            I => \N__33959\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__34046\,
            I => \N__33956\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__34041\,
            I => \N__33953\
        );

    \I__8473\ : SRMux
    port map (
            O => \N__34040\,
            I => \N__33852\
        );

    \I__8472\ : SRMux
    port map (
            O => \N__34039\,
            I => \N__33852\
        );

    \I__8471\ : SRMux
    port map (
            O => \N__34038\,
            I => \N__33852\
        );

    \I__8470\ : SRMux
    port map (
            O => \N__34037\,
            I => \N__33852\
        );

    \I__8469\ : SRMux
    port map (
            O => \N__34036\,
            I => \N__33852\
        );

    \I__8468\ : SRMux
    port map (
            O => \N__34035\,
            I => \N__33852\
        );

    \I__8467\ : SRMux
    port map (
            O => \N__34034\,
            I => \N__33852\
        );

    \I__8466\ : SRMux
    port map (
            O => \N__34033\,
            I => \N__33852\
        );

    \I__8465\ : SRMux
    port map (
            O => \N__34032\,
            I => \N__33852\
        );

    \I__8464\ : SRMux
    port map (
            O => \N__34031\,
            I => \N__33852\
        );

    \I__8463\ : SRMux
    port map (
            O => \N__34030\,
            I => \N__33852\
        );

    \I__8462\ : SRMux
    port map (
            O => \N__34029\,
            I => \N__33852\
        );

    \I__8461\ : SRMux
    port map (
            O => \N__34028\,
            I => \N__33852\
        );

    \I__8460\ : SRMux
    port map (
            O => \N__34027\,
            I => \N__33852\
        );

    \I__8459\ : SRMux
    port map (
            O => \N__34026\,
            I => \N__33852\
        );

    \I__8458\ : SRMux
    port map (
            O => \N__34025\,
            I => \N__33852\
        );

    \I__8457\ : SRMux
    port map (
            O => \N__34024\,
            I => \N__33852\
        );

    \I__8456\ : SRMux
    port map (
            O => \N__34023\,
            I => \N__33852\
        );

    \I__8455\ : SRMux
    port map (
            O => \N__34022\,
            I => \N__33852\
        );

    \I__8454\ : SRMux
    port map (
            O => \N__34021\,
            I => \N__33852\
        );

    \I__8453\ : SRMux
    port map (
            O => \N__34020\,
            I => \N__33852\
        );

    \I__8452\ : SRMux
    port map (
            O => \N__34019\,
            I => \N__33852\
        );

    \I__8451\ : SRMux
    port map (
            O => \N__34018\,
            I => \N__33852\
        );

    \I__8450\ : SRMux
    port map (
            O => \N__34017\,
            I => \N__33852\
        );

    \I__8449\ : SRMux
    port map (
            O => \N__34016\,
            I => \N__33852\
        );

    \I__8448\ : SRMux
    port map (
            O => \N__34015\,
            I => \N__33852\
        );

    \I__8447\ : SRMux
    port map (
            O => \N__34014\,
            I => \N__33852\
        );

    \I__8446\ : SRMux
    port map (
            O => \N__34013\,
            I => \N__33852\
        );

    \I__8445\ : SRMux
    port map (
            O => \N__34012\,
            I => \N__33852\
        );

    \I__8444\ : SRMux
    port map (
            O => \N__34011\,
            I => \N__33852\
        );

    \I__8443\ : SRMux
    port map (
            O => \N__34010\,
            I => \N__33852\
        );

    \I__8442\ : Glb2LocalMux
    port map (
            O => \N__34007\,
            I => \N__33852\
        );

    \I__8441\ : Glb2LocalMux
    port map (
            O => \N__34004\,
            I => \N__33852\
        );

    \I__8440\ : Glb2LocalMux
    port map (
            O => \N__34001\,
            I => \N__33852\
        );

    \I__8439\ : Glb2LocalMux
    port map (
            O => \N__33998\,
            I => \N__33852\
        );

    \I__8438\ : Glb2LocalMux
    port map (
            O => \N__33995\,
            I => \N__33852\
        );

    \I__8437\ : Glb2LocalMux
    port map (
            O => \N__33992\,
            I => \N__33852\
        );

    \I__8436\ : Glb2LocalMux
    port map (
            O => \N__33989\,
            I => \N__33852\
        );

    \I__8435\ : Glb2LocalMux
    port map (
            O => \N__33986\,
            I => \N__33852\
        );

    \I__8434\ : Glb2LocalMux
    port map (
            O => \N__33983\,
            I => \N__33852\
        );

    \I__8433\ : Glb2LocalMux
    port map (
            O => \N__33980\,
            I => \N__33852\
        );

    \I__8432\ : Glb2LocalMux
    port map (
            O => \N__33977\,
            I => \N__33852\
        );

    \I__8431\ : Glb2LocalMux
    port map (
            O => \N__33974\,
            I => \N__33852\
        );

    \I__8430\ : Glb2LocalMux
    port map (
            O => \N__33971\,
            I => \N__33852\
        );

    \I__8429\ : Glb2LocalMux
    port map (
            O => \N__33968\,
            I => \N__33852\
        );

    \I__8428\ : Glb2LocalMux
    port map (
            O => \N__33965\,
            I => \N__33852\
        );

    \I__8427\ : Glb2LocalMux
    port map (
            O => \N__33962\,
            I => \N__33852\
        );

    \I__8426\ : Glb2LocalMux
    port map (
            O => \N__33959\,
            I => \N__33852\
        );

    \I__8425\ : Glb2LocalMux
    port map (
            O => \N__33956\,
            I => \N__33852\
        );

    \I__8424\ : Glb2LocalMux
    port map (
            O => \N__33953\,
            I => \N__33852\
        );

    \I__8423\ : GlobalMux
    port map (
            O => \N__33852\,
            I => \N__33849\
        );

    \I__8422\ : gio2CtrlBuf
    port map (
            O => \N__33849\,
            I => \M_this_reset_cond_out_g_0\
        );

    \I__8421\ : InMux
    port map (
            O => \N__33846\,
            I => \N__33843\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__33843\,
            I => \N__33840\
        );

    \I__8419\ : Span4Mux_v
    port map (
            O => \N__33840\,
            I => \N__33837\
        );

    \I__8418\ : Odrv4
    port map (
            O => \N__33837\,
            I => \un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0\
        );

    \I__8417\ : CascadeMux
    port map (
            O => \N__33834\,
            I => \N__33830\
        );

    \I__8416\ : CascadeMux
    port map (
            O => \N__33833\,
            I => \N__33827\
        );

    \I__8415\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33822\
        );

    \I__8414\ : InMux
    port map (
            O => \N__33827\,
            I => \N__33819\
        );

    \I__8413\ : InMux
    port map (
            O => \N__33826\,
            I => \N__33815\
        );

    \I__8412\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33810\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__33822\,
            I => \N__33807\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__33819\,
            I => \N__33804\
        );

    \I__8409\ : CascadeMux
    port map (
            O => \N__33818\,
            I => \N__33801\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__33815\,
            I => \N__33796\
        );

    \I__8407\ : InMux
    port map (
            O => \N__33814\,
            I => \N__33791\
        );

    \I__8406\ : InMux
    port map (
            O => \N__33813\,
            I => \N__33791\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__33810\,
            I => \N__33788\
        );

    \I__8404\ : Span4Mux_v
    port map (
            O => \N__33807\,
            I => \N__33785\
        );

    \I__8403\ : Span4Mux_h
    port map (
            O => \N__33804\,
            I => \N__33782\
        );

    \I__8402\ : InMux
    port map (
            O => \N__33801\,
            I => \N__33779\
        );

    \I__8401\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33776\
        );

    \I__8400\ : InMux
    port map (
            O => \N__33799\,
            I => \N__33773\
        );

    \I__8399\ : Span4Mux_v
    port map (
            O => \N__33796\,
            I => \N__33770\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__33791\,
            I => \N__33767\
        );

    \I__8397\ : Span4Mux_v
    port map (
            O => \N__33788\,
            I => \N__33764\
        );

    \I__8396\ : Span4Mux_h
    port map (
            O => \N__33785\,
            I => \N__33757\
        );

    \I__8395\ : Span4Mux_v
    port map (
            O => \N__33782\,
            I => \N__33757\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__33779\,
            I => \N__33757\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__33776\,
            I => \N__33754\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__33773\,
            I => \N__33751\
        );

    \I__8391\ : Sp12to4
    port map (
            O => \N__33770\,
            I => \N__33745\
        );

    \I__8390\ : Span12Mux_v
    port map (
            O => \N__33767\,
            I => \N__33745\
        );

    \I__8389\ : Span4Mux_v
    port map (
            O => \N__33764\,
            I => \N__33742\
        );

    \I__8388\ : Span4Mux_h
    port map (
            O => \N__33757\,
            I => \N__33739\
        );

    \I__8387\ : Span4Mux_v
    port map (
            O => \N__33754\,
            I => \N__33734\
        );

    \I__8386\ : Span4Mux_v
    port map (
            O => \N__33751\,
            I => \N__33734\
        );

    \I__8385\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33731\
        );

    \I__8384\ : Span12Mux_h
    port map (
            O => \N__33745\,
            I => \N__33728\
        );

    \I__8383\ : Sp12to4
    port map (
            O => \N__33742\,
            I => \N__33725\
        );

    \I__8382\ : Span4Mux_v
    port map (
            O => \N__33739\,
            I => \N__33722\
        );

    \I__8381\ : Span4Mux_h
    port map (
            O => \N__33734\,
            I => \N__33717\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__33731\,
            I => \N__33717\
        );

    \I__8379\ : Span12Mux_v
    port map (
            O => \N__33728\,
            I => \N__33714\
        );

    \I__8378\ : Span12Mux_h
    port map (
            O => \N__33725\,
            I => \N__33711\
        );

    \I__8377\ : Span4Mux_h
    port map (
            O => \N__33722\,
            I => \N__33708\
        );

    \I__8376\ : Sp12to4
    port map (
            O => \N__33717\,
            I => \N__33705\
        );

    \I__8375\ : Odrv12
    port map (
            O => \N__33714\,
            I => port_data_c_0
        );

    \I__8374\ : Odrv12
    port map (
            O => \N__33711\,
            I => port_data_c_0
        );

    \I__8373\ : Odrv4
    port map (
            O => \N__33708\,
            I => port_data_c_0
        );

    \I__8372\ : Odrv12
    port map (
            O => \N__33705\,
            I => port_data_c_0
        );

    \I__8371\ : IoInMux
    port map (
            O => \N__33696\,
            I => \N__33692\
        );

    \I__8370\ : InMux
    port map (
            O => \N__33695\,
            I => \N__33689\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__33692\,
            I => \N__33686\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__33689\,
            I => \N__33683\
        );

    \I__8367\ : Span12Mux_s10_v
    port map (
            O => \N__33686\,
            I => \N__33680\
        );

    \I__8366\ : Span4Mux_h
    port map (
            O => \N__33683\,
            I => \N__33677\
        );

    \I__8365\ : Odrv12
    port map (
            O => \N__33680\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__8364\ : Odrv4
    port map (
            O => \N__33677\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__8363\ : InMux
    port map (
            O => \N__33672\,
            I => \N__33665\
        );

    \I__8362\ : InMux
    port map (
            O => \N__33671\,
            I => \N__33662\
        );

    \I__8361\ : InMux
    port map (
            O => \N__33670\,
            I => \N__33659\
        );

    \I__8360\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33654\
        );

    \I__8359\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33651\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__33665\,
            I => \N__33644\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__33662\,
            I => \N__33644\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__33659\,
            I => \N__33644\
        );

    \I__8355\ : CascadeMux
    port map (
            O => \N__33658\,
            I => \N__33641\
        );

    \I__8354\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33638\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__33654\,
            I => \N__33634\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__33651\,
            I => \N__33631\
        );

    \I__8351\ : Span4Mux_v
    port map (
            O => \N__33644\,
            I => \N__33626\
        );

    \I__8350\ : InMux
    port map (
            O => \N__33641\,
            I => \N__33623\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__33638\,
            I => \N__33620\
        );

    \I__8348\ : CascadeMux
    port map (
            O => \N__33637\,
            I => \N__33617\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__33634\,
            I => \N__33614\
        );

    \I__8346\ : Span4Mux_v
    port map (
            O => \N__33631\,
            I => \N__33611\
        );

    \I__8345\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33608\
        );

    \I__8344\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33605\
        );

    \I__8343\ : Sp12to4
    port map (
            O => \N__33626\,
            I => \N__33600\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__33623\,
            I => \N__33600\
        );

    \I__8341\ : Span12Mux_s10_v
    port map (
            O => \N__33620\,
            I => \N__33597\
        );

    \I__8340\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33594\
        );

    \I__8339\ : Span4Mux_h
    port map (
            O => \N__33614\,
            I => \N__33589\
        );

    \I__8338\ : Span4Mux_h
    port map (
            O => \N__33611\,
            I => \N__33589\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__33608\,
            I => \N__33584\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__33605\,
            I => \N__33584\
        );

    \I__8335\ : Span12Mux_v
    port map (
            O => \N__33600\,
            I => \N__33581\
        );

    \I__8334\ : Span12Mux_v
    port map (
            O => \N__33597\,
            I => \N__33578\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__33594\,
            I => \N__33575\
        );

    \I__8332\ : IoSpan4Mux
    port map (
            O => \N__33589\,
            I => \N__33572\
        );

    \I__8331\ : Span4Mux_v
    port map (
            O => \N__33584\,
            I => \N__33569\
        );

    \I__8330\ : Span12Mux_h
    port map (
            O => \N__33581\,
            I => \N__33566\
        );

    \I__8329\ : Span12Mux_h
    port map (
            O => \N__33578\,
            I => \N__33561\
        );

    \I__8328\ : Span12Mux_v
    port map (
            O => \N__33575\,
            I => \N__33561\
        );

    \I__8327\ : IoSpan4Mux
    port map (
            O => \N__33572\,
            I => \N__33558\
        );

    \I__8326\ : Sp12to4
    port map (
            O => \N__33569\,
            I => \N__33555\
        );

    \I__8325\ : Odrv12
    port map (
            O => \N__33566\,
            I => port_data_c_7
        );

    \I__8324\ : Odrv12
    port map (
            O => \N__33561\,
            I => port_data_c_7
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__33558\,
            I => port_data_c_7
        );

    \I__8322\ : Odrv12
    port map (
            O => \N__33555\,
            I => port_data_c_7
        );

    \I__8321\ : InMux
    port map (
            O => \N__33546\,
            I => \N__33543\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__33543\,
            I => \N__33540\
        );

    \I__8319\ : Span4Mux_h
    port map (
            O => \N__33540\,
            I => \N__33537\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__33537\,
            I => \un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0\
        );

    \I__8317\ : IoInMux
    port map (
            O => \N__33534\,
            I => \N__33531\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__8315\ : Span4Mux_s2_h
    port map (
            O => \N__33528\,
            I => \N__33525\
        );

    \I__8314\ : Span4Mux_h
    port map (
            O => \N__33525\,
            I => \N__33521\
        );

    \I__8313\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33518\
        );

    \I__8312\ : Sp12to4
    port map (
            O => \N__33521\,
            I => \N__33515\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__33518\,
            I => \N__33512\
        );

    \I__8310\ : Span12Mux_v
    port map (
            O => \N__33515\,
            I => \N__33509\
        );

    \I__8309\ : Span4Mux_h
    port map (
            O => \N__33512\,
            I => \N__33506\
        );

    \I__8308\ : Odrv12
    port map (
            O => \N__33509\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__8307\ : Odrv4
    port map (
            O => \N__33506\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__8306\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33498\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__33498\,
            I => \N__33495\
        );

    \I__8304\ : Odrv4
    port map (
            O => \N__33495\,
            I => \un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0\
        );

    \I__8303\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33488\
        );

    \I__8302\ : CascadeMux
    port map (
            O => \N__33491\,
            I => \N__33484\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__33488\,
            I => \N__33479\
        );

    \I__8300\ : InMux
    port map (
            O => \N__33487\,
            I => \N__33476\
        );

    \I__8299\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33473\
        );

    \I__8298\ : CascadeMux
    port map (
            O => \N__33483\,
            I => \N__33468\
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__33482\,
            I => \N__33465\
        );

    \I__8296\ : Span4Mux_h
    port map (
            O => \N__33479\,
            I => \N__33458\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__33476\,
            I => \N__33458\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__33473\,
            I => \N__33458\
        );

    \I__8293\ : InMux
    port map (
            O => \N__33472\,
            I => \N__33455\
        );

    \I__8292\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33451\
        );

    \I__8291\ : InMux
    port map (
            O => \N__33468\,
            I => \N__33448\
        );

    \I__8290\ : InMux
    port map (
            O => \N__33465\,
            I => \N__33445\
        );

    \I__8289\ : Span4Mux_h
    port map (
            O => \N__33458\,
            I => \N__33440\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__33455\,
            I => \N__33437\
        );

    \I__8287\ : InMux
    port map (
            O => \N__33454\,
            I => \N__33434\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__33451\,
            I => \N__33431\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__33448\,
            I => \N__33428\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__33445\,
            I => \N__33425\
        );

    \I__8283\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33422\
        );

    \I__8282\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33417\
        );

    \I__8281\ : Span4Mux_h
    port map (
            O => \N__33440\,
            I => \N__33414\
        );

    \I__8280\ : Span4Mux_h
    port map (
            O => \N__33437\,
            I => \N__33411\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__33434\,
            I => \N__33408\
        );

    \I__8278\ : Span4Mux_v
    port map (
            O => \N__33431\,
            I => \N__33401\
        );

    \I__8277\ : Span4Mux_h
    port map (
            O => \N__33428\,
            I => \N__33401\
        );

    \I__8276\ : Span4Mux_v
    port map (
            O => \N__33425\,
            I => \N__33401\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__33422\,
            I => \N__33398\
        );

    \I__8274\ : CascadeMux
    port map (
            O => \N__33421\,
            I => \N__33395\
        );

    \I__8273\ : CascadeMux
    port map (
            O => \N__33420\,
            I => \N__33391\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__33417\,
            I => \N__33388\
        );

    \I__8271\ : Span4Mux_h
    port map (
            O => \N__33414\,
            I => \N__33383\
        );

    \I__8270\ : Span4Mux_v
    port map (
            O => \N__33411\,
            I => \N__33383\
        );

    \I__8269\ : Span4Mux_h
    port map (
            O => \N__33408\,
            I => \N__33380\
        );

    \I__8268\ : Span4Mux_h
    port map (
            O => \N__33401\,
            I => \N__33375\
        );

    \I__8267\ : Span4Mux_v
    port map (
            O => \N__33398\,
            I => \N__33375\
        );

    \I__8266\ : InMux
    port map (
            O => \N__33395\,
            I => \N__33372\
        );

    \I__8265\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33369\
        );

    \I__8264\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33366\
        );

    \I__8263\ : Span12Mux_h
    port map (
            O => \N__33388\,
            I => \N__33363\
        );

    \I__8262\ : Span4Mux_v
    port map (
            O => \N__33383\,
            I => \N__33360\
        );

    \I__8261\ : Span4Mux_h
    port map (
            O => \N__33380\,
            I => \N__33357\
        );

    \I__8260\ : Span4Mux_h
    port map (
            O => \N__33375\,
            I => \N__33348\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__33372\,
            I => \N__33348\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__33369\,
            I => \N__33348\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__33366\,
            I => \N__33348\
        );

    \I__8256\ : Span12Mux_h
    port map (
            O => \N__33363\,
            I => \N__33345\
        );

    \I__8255\ : Span4Mux_v
    port map (
            O => \N__33360\,
            I => \N__33342\
        );

    \I__8254\ : Sp12to4
    port map (
            O => \N__33357\,
            I => \N__33337\
        );

    \I__8253\ : Sp12to4
    port map (
            O => \N__33348\,
            I => \N__33337\
        );

    \I__8252\ : Odrv12
    port map (
            O => \N__33345\,
            I => port_data_c_2
        );

    \I__8251\ : Odrv4
    port map (
            O => \N__33342\,
            I => port_data_c_2
        );

    \I__8250\ : Odrv12
    port map (
            O => \N__33337\,
            I => port_data_c_2
        );

    \I__8249\ : IoInMux
    port map (
            O => \N__33330\,
            I => \N__33327\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__33327\,
            I => \N__33324\
        );

    \I__8247\ : IoSpan4Mux
    port map (
            O => \N__33324\,
            I => \N__33321\
        );

    \I__8246\ : Span4Mux_s1_v
    port map (
            O => \N__33321\,
            I => \N__33318\
        );

    \I__8245\ : Span4Mux_v
    port map (
            O => \N__33318\,
            I => \N__33314\
        );

    \I__8244\ : InMux
    port map (
            O => \N__33317\,
            I => \N__33311\
        );

    \I__8243\ : Span4Mux_v
    port map (
            O => \N__33314\,
            I => \N__33306\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__33311\,
            I => \N__33306\
        );

    \I__8241\ : Odrv4
    port map (
            O => \N__33306\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__8240\ : InMux
    port map (
            O => \N__33303\,
            I => \N__33300\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__33300\,
            I => \N__33297\
        );

    \I__8238\ : Span4Mux_v
    port map (
            O => \N__33297\,
            I => \N__33293\
        );

    \I__8237\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33290\
        );

    \I__8236\ : Sp12to4
    port map (
            O => \N__33293\,
            I => \N__33285\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__33290\,
            I => \N__33285\
        );

    \I__8234\ : Span12Mux_s11_h
    port map (
            O => \N__33285\,
            I => \N__33282\
        );

    \I__8233\ : Odrv12
    port map (
            O => \N__33282\,
            I => \un1_M_this_state_q_11_0_i\
        );

    \I__8232\ : IoInMux
    port map (
            O => \N__33279\,
            I => \N__33276\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__33276\,
            I => \N__33273\
        );

    \I__8230\ : IoSpan4Mux
    port map (
            O => \N__33273\,
            I => \N__33269\
        );

    \I__8229\ : CascadeMux
    port map (
            O => \N__33272\,
            I => \N__33266\
        );

    \I__8228\ : IoSpan4Mux
    port map (
            O => \N__33269\,
            I => \N__33263\
        );

    \I__8227\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33259\
        );

    \I__8226\ : IoSpan4Mux
    port map (
            O => \N__33263\,
            I => \N__33256\
        );

    \I__8225\ : CascadeMux
    port map (
            O => \N__33262\,
            I => \N__33253\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__33259\,
            I => \N__33250\
        );

    \I__8223\ : Sp12to4
    port map (
            O => \N__33256\,
            I => \N__33247\
        );

    \I__8222\ : InMux
    port map (
            O => \N__33253\,
            I => \N__33244\
        );

    \I__8221\ : Span4Mux_v
    port map (
            O => \N__33250\,
            I => \N__33241\
        );

    \I__8220\ : Odrv12
    port map (
            O => \N__33247\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__33244\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__8218\ : Odrv4
    port map (
            O => \N__33241\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__8217\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33231\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__33231\,
            I => \N__33228\
        );

    \I__8215\ : Span4Mux_h
    port map (
            O => \N__33228\,
            I => \N__33225\
        );

    \I__8214\ : Odrv4
    port map (
            O => \N__33225\,
            I => \un1_M_this_external_address_q_cry_0_THRU_CO\
        );

    \I__8213\ : InMux
    port map (
            O => \N__33222\,
            I => \N__33217\
        );

    \I__8212\ : IoInMux
    port map (
            O => \N__33221\,
            I => \N__33214\
        );

    \I__8211\ : CascadeMux
    port map (
            O => \N__33220\,
            I => \N__33211\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__33217\,
            I => \N__33208\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__33214\,
            I => \N__33205\
        );

    \I__8208\ : InMux
    port map (
            O => \N__33211\,
            I => \N__33202\
        );

    \I__8207\ : Span4Mux_h
    port map (
            O => \N__33208\,
            I => \N__33199\
        );

    \I__8206\ : Odrv12
    port map (
            O => \N__33205\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__33202\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__8204\ : Odrv4
    port map (
            O => \N__33199\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__8203\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33189\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__33189\,
            I => \N__33186\
        );

    \I__8201\ : Span4Mux_h
    port map (
            O => \N__33186\,
            I => \N__33183\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__33183\,
            I => \un1_M_this_external_address_q_cry_1_THRU_CO\
        );

    \I__8199\ : IoInMux
    port map (
            O => \N__33180\,
            I => \N__33177\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__33177\,
            I => \N__33174\
        );

    \I__8197\ : IoSpan4Mux
    port map (
            O => \N__33174\,
            I => \N__33169\
        );

    \I__8196\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33166\
        );

    \I__8195\ : CascadeMux
    port map (
            O => \N__33172\,
            I => \N__33163\
        );

    \I__8194\ : Span4Mux_s2_v
    port map (
            O => \N__33169\,
            I => \N__33160\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__33166\,
            I => \N__33157\
        );

    \I__8192\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33154\
        );

    \I__8191\ : Span4Mux_v
    port map (
            O => \N__33160\,
            I => \N__33149\
        );

    \I__8190\ : Span4Mux_h
    port map (
            O => \N__33157\,
            I => \N__33149\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__33154\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__8188\ : Odrv4
    port map (
            O => \N__33149\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__8187\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33141\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__33141\,
            I => \N__33138\
        );

    \I__8185\ : Span4Mux_h
    port map (
            O => \N__33138\,
            I => \N__33135\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__33135\,
            I => \un1_M_this_external_address_q_cry_2_THRU_CO\
        );

    \I__8183\ : IoInMux
    port map (
            O => \N__33132\,
            I => \N__33129\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__33129\,
            I => \N__33126\
        );

    \I__8181\ : IoSpan4Mux
    port map (
            O => \N__33126\,
            I => \N__33121\
        );

    \I__8180\ : InMux
    port map (
            O => \N__33125\,
            I => \N__33118\
        );

    \I__8179\ : CascadeMux
    port map (
            O => \N__33124\,
            I => \N__33115\
        );

    \I__8178\ : Span4Mux_s1_h
    port map (
            O => \N__33121\,
            I => \N__33112\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__33118\,
            I => \N__33109\
        );

    \I__8176\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33106\
        );

    \I__8175\ : Span4Mux_h
    port map (
            O => \N__33112\,
            I => \N__33101\
        );

    \I__8174\ : Span4Mux_h
    port map (
            O => \N__33109\,
            I => \N__33101\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__33106\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__8172\ : Odrv4
    port map (
            O => \N__33101\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__8171\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33093\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__33093\,
            I => \N__33090\
        );

    \I__8169\ : Span4Mux_v
    port map (
            O => \N__33090\,
            I => \N__33087\
        );

    \I__8168\ : Odrv4
    port map (
            O => \N__33087\,
            I => \un1_M_this_external_address_q_cry_3_THRU_CO\
        );

    \I__8167\ : InMux
    port map (
            O => \N__33084\,
            I => \N__33079\
        );

    \I__8166\ : IoInMux
    port map (
            O => \N__33083\,
            I => \N__33076\
        );

    \I__8165\ : CascadeMux
    port map (
            O => \N__33082\,
            I => \N__33073\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__33079\,
            I => \N__33070\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__33076\,
            I => \N__33067\
        );

    \I__8162\ : InMux
    port map (
            O => \N__33073\,
            I => \N__33064\
        );

    \I__8161\ : Span4Mux_v
    port map (
            O => \N__33070\,
            I => \N__33061\
        );

    \I__8160\ : Odrv12
    port map (
            O => \N__33067\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__33064\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__33061\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__8157\ : InMux
    port map (
            O => \N__33054\,
            I => \N__33051\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__33048\
        );

    \I__8155\ : Span4Mux_v
    port map (
            O => \N__33048\,
            I => \N__33045\
        );

    \I__8154\ : Odrv4
    port map (
            O => \N__33045\,
            I => \un1_M_this_external_address_q_cry_4_THRU_CO\
        );

    \I__8153\ : IoInMux
    port map (
            O => \N__33042\,
            I => \N__33039\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__33039\,
            I => \N__33035\
        );

    \I__8151\ : InMux
    port map (
            O => \N__33038\,
            I => \N__33031\
        );

    \I__8150\ : Span4Mux_s1_h
    port map (
            O => \N__33035\,
            I => \N__33028\
        );

    \I__8149\ : CascadeMux
    port map (
            O => \N__33034\,
            I => \N__33025\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__33031\,
            I => \N__33022\
        );

    \I__8147\ : Span4Mux_h
    port map (
            O => \N__33028\,
            I => \N__33019\
        );

    \I__8146\ : InMux
    port map (
            O => \N__33025\,
            I => \N__33016\
        );

    \I__8145\ : Span4Mux_h
    port map (
            O => \N__33022\,
            I => \N__33013\
        );

    \I__8144\ : Odrv4
    port map (
            O => \N__33019\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__33016\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__8142\ : Odrv4
    port map (
            O => \N__33013\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__8141\ : CascadeMux
    port map (
            O => \N__33006\,
            I => \N__33003\
        );

    \I__8140\ : InMux
    port map (
            O => \N__33003\,
            I => \N__33000\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__33000\,
            I => \N__32997\
        );

    \I__8138\ : Odrv12
    port map (
            O => \N__32997\,
            I => \M_this_data_tmp_qZ0Z_23\
        );

    \I__8137\ : InMux
    port map (
            O => \N__32994\,
            I => \N__32991\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__32991\,
            I => \M_this_oam_ram_write_data_23\
        );

    \I__8135\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32982\
        );

    \I__8134\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32978\
        );

    \I__8133\ : CascadeMux
    port map (
            O => \N__32986\,
            I => \N__32975\
        );

    \I__8132\ : CascadeMux
    port map (
            O => \N__32985\,
            I => \N__32972\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__32982\,
            I => \N__32968\
        );

    \I__8130\ : InMux
    port map (
            O => \N__32981\,
            I => \N__32965\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__32978\,
            I => \N__32962\
        );

    \I__8128\ : InMux
    port map (
            O => \N__32975\,
            I => \N__32959\
        );

    \I__8127\ : InMux
    port map (
            O => \N__32972\,
            I => \N__32956\
        );

    \I__8126\ : CascadeMux
    port map (
            O => \N__32971\,
            I => \N__32951\
        );

    \I__8125\ : Span4Mux_h
    port map (
            O => \N__32968\,
            I => \N__32946\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__32965\,
            I => \N__32946\
        );

    \I__8123\ : Span4Mux_v
    port map (
            O => \N__32962\,
            I => \N__32941\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__32959\,
            I => \N__32941\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__32956\,
            I => \N__32938\
        );

    \I__8120\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32935\
        );

    \I__8119\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32930\
        );

    \I__8118\ : InMux
    port map (
            O => \N__32951\,
            I => \N__32930\
        );

    \I__8117\ : Span4Mux_v
    port map (
            O => \N__32946\,
            I => \N__32927\
        );

    \I__8116\ : Span4Mux_v
    port map (
            O => \N__32941\,
            I => \N__32923\
        );

    \I__8115\ : Span4Mux_v
    port map (
            O => \N__32938\,
            I => \N__32918\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__32935\,
            I => \N__32918\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__32930\,
            I => \N__32913\
        );

    \I__8112\ : Span4Mux_h
    port map (
            O => \N__32927\,
            I => \N__32909\
        );

    \I__8111\ : InMux
    port map (
            O => \N__32926\,
            I => \N__32906\
        );

    \I__8110\ : Span4Mux_h
    port map (
            O => \N__32923\,
            I => \N__32901\
        );

    \I__8109\ : Span4Mux_v
    port map (
            O => \N__32918\,
            I => \N__32901\
        );

    \I__8108\ : InMux
    port map (
            O => \N__32917\,
            I => \N__32898\
        );

    \I__8107\ : InMux
    port map (
            O => \N__32916\,
            I => \N__32895\
        );

    \I__8106\ : Span4Mux_v
    port map (
            O => \N__32913\,
            I => \N__32892\
        );

    \I__8105\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32889\
        );

    \I__8104\ : Sp12to4
    port map (
            O => \N__32909\,
            I => \N__32878\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__32906\,
            I => \N__32878\
        );

    \I__8102\ : Sp12to4
    port map (
            O => \N__32901\,
            I => \N__32878\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__32898\,
            I => \N__32878\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__32895\,
            I => \N__32878\
        );

    \I__8099\ : Span4Mux_h
    port map (
            O => \N__32892\,
            I => \N__32873\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__32889\,
            I => \N__32873\
        );

    \I__8097\ : Span12Mux_h
    port map (
            O => \N__32878\,
            I => \N__32868\
        );

    \I__8096\ : Sp12to4
    port map (
            O => \N__32873\,
            I => \N__32868\
        );

    \I__8095\ : Odrv12
    port map (
            O => \N__32868\,
            I => port_data_c_1
        );

    \I__8094\ : InMux
    port map (
            O => \N__32865\,
            I => \N__32862\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__32862\,
            I => \N_41_0\
        );

    \I__8092\ : CascadeMux
    port map (
            O => \N__32859\,
            I => \N__32856\
        );

    \I__8091\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32853\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__32853\,
            I => \N__32850\
        );

    \I__8089\ : Odrv12
    port map (
            O => \N__32850\,
            I => \M_this_data_tmp_qZ0Z_2\
        );

    \I__8088\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32844\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__32844\,
            I => \N__32841\
        );

    \I__8086\ : Span4Mux_h
    port map (
            O => \N__32841\,
            I => \N__32838\
        );

    \I__8085\ : Odrv4
    port map (
            O => \N__32838\,
            I => \un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0\
        );

    \I__8084\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32827\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__32834\,
            I => \N__32824\
        );

    \I__8082\ : InMux
    port map (
            O => \N__32833\,
            I => \N__32820\
        );

    \I__8081\ : CascadeMux
    port map (
            O => \N__32832\,
            I => \N__32817\
        );

    \I__8080\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32814\
        );

    \I__8079\ : CascadeMux
    port map (
            O => \N__32830\,
            I => \N__32811\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__32827\,
            I => \N__32808\
        );

    \I__8077\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32805\
        );

    \I__8076\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32802\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__32820\,
            I => \N__32796\
        );

    \I__8074\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32793\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__32814\,
            I => \N__32790\
        );

    \I__8072\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32787\
        );

    \I__8071\ : Span4Mux_v
    port map (
            O => \N__32808\,
            I => \N__32782\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__32805\,
            I => \N__32782\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__32802\,
            I => \N__32779\
        );

    \I__8068\ : InMux
    port map (
            O => \N__32801\,
            I => \N__32776\
        );

    \I__8067\ : InMux
    port map (
            O => \N__32800\,
            I => \N__32773\
        );

    \I__8066\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32770\
        );

    \I__8065\ : Span4Mux_v
    port map (
            O => \N__32796\,
            I => \N__32767\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__32793\,
            I => \N__32764\
        );

    \I__8063\ : Span4Mux_h
    port map (
            O => \N__32790\,
            I => \N__32759\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__32787\,
            I => \N__32759\
        );

    \I__8061\ : Span4Mux_h
    port map (
            O => \N__32782\,
            I => \N__32756\
        );

    \I__8060\ : Span4Mux_v
    port map (
            O => \N__32779\,
            I => \N__32751\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__32776\,
            I => \N__32751\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__32773\,
            I => \N__32748\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__32770\,
            I => \N__32745\
        );

    \I__8056\ : Sp12to4
    port map (
            O => \N__32767\,
            I => \N__32742\
        );

    \I__8055\ : Span4Mux_v
    port map (
            O => \N__32764\,
            I => \N__32739\
        );

    \I__8054\ : Span4Mux_v
    port map (
            O => \N__32759\,
            I => \N__32736\
        );

    \I__8053\ : Span4Mux_v
    port map (
            O => \N__32756\,
            I => \N__32731\
        );

    \I__8052\ : Span4Mux_h
    port map (
            O => \N__32751\,
            I => \N__32731\
        );

    \I__8051\ : Span12Mux_h
    port map (
            O => \N__32748\,
            I => \N__32728\
        );

    \I__8050\ : Span12Mux_v
    port map (
            O => \N__32745\,
            I => \N__32725\
        );

    \I__8049\ : Span12Mux_h
    port map (
            O => \N__32742\,
            I => \N__32720\
        );

    \I__8048\ : Sp12to4
    port map (
            O => \N__32739\,
            I => \N__32720\
        );

    \I__8047\ : Sp12to4
    port map (
            O => \N__32736\,
            I => \N__32717\
        );

    \I__8046\ : Span4Mux_v
    port map (
            O => \N__32731\,
            I => \N__32714\
        );

    \I__8045\ : Span12Mux_v
    port map (
            O => \N__32728\,
            I => \N__32709\
        );

    \I__8044\ : Span12Mux_h
    port map (
            O => \N__32725\,
            I => \N__32709\
        );

    \I__8043\ : Span12Mux_h
    port map (
            O => \N__32720\,
            I => \N__32706\
        );

    \I__8042\ : Span12Mux_h
    port map (
            O => \N__32717\,
            I => \N__32703\
        );

    \I__8041\ : Span4Mux_h
    port map (
            O => \N__32714\,
            I => \N__32700\
        );

    \I__8040\ : Odrv12
    port map (
            O => \N__32709\,
            I => port_data_c_3
        );

    \I__8039\ : Odrv12
    port map (
            O => \N__32706\,
            I => port_data_c_3
        );

    \I__8038\ : Odrv12
    port map (
            O => \N__32703\,
            I => port_data_c_3
        );

    \I__8037\ : Odrv4
    port map (
            O => \N__32700\,
            I => port_data_c_3
        );

    \I__8036\ : IoInMux
    port map (
            O => \N__32691\,
            I => \N__32688\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__32688\,
            I => \N__32685\
        );

    \I__8034\ : Span4Mux_s2_v
    port map (
            O => \N__32685\,
            I => \N__32681\
        );

    \I__8033\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32678\
        );

    \I__8032\ : Span4Mux_v
    port map (
            O => \N__32681\,
            I => \N__32675\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__32678\,
            I => \N__32672\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__32675\,
            I => \N__32669\
        );

    \I__8029\ : Span4Mux_h
    port map (
            O => \N__32672\,
            I => \N__32666\
        );

    \I__8028\ : Odrv4
    port map (
            O => \N__32669\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__8027\ : Odrv4
    port map (
            O => \N__32666\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__8026\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32658\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__32658\,
            I => \N__32655\
        );

    \I__8024\ : Odrv4
    port map (
            O => \N__32655\,
            I => \un1_M_this_external_address_q_cry_6_THRU_CO\
        );

    \I__8023\ : IoInMux
    port map (
            O => \N__32652\,
            I => \N__32649\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__32649\,
            I => \N__32646\
        );

    \I__8021\ : IoSpan4Mux
    port map (
            O => \N__32646\,
            I => \N__32643\
        );

    \I__8020\ : Span4Mux_s2_h
    port map (
            O => \N__32643\,
            I => \N__32640\
        );

    \I__8019\ : Span4Mux_h
    port map (
            O => \N__32640\,
            I => \N__32637\
        );

    \I__8018\ : Sp12to4
    port map (
            O => \N__32637\,
            I => \N__32632\
        );

    \I__8017\ : CascadeMux
    port map (
            O => \N__32636\,
            I => \N__32629\
        );

    \I__8016\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32626\
        );

    \I__8015\ : Span12Mux_v
    port map (
            O => \N__32632\,
            I => \N__32623\
        );

    \I__8014\ : InMux
    port map (
            O => \N__32629\,
            I => \N__32620\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32617\
        );

    \I__8012\ : Odrv12
    port map (
            O => \N__32623\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__32620\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__8010\ : Odrv4
    port map (
            O => \N__32617\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__8009\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32607\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__32607\,
            I => \N__32604\
        );

    \I__8007\ : Span4Mux_h
    port map (
            O => \N__32604\,
            I => \N__32601\
        );

    \I__8006\ : Odrv4
    port map (
            O => \N__32601\,
            I => \un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0\
        );

    \I__8005\ : CascadeMux
    port map (
            O => \N__32598\,
            I => \N__32595\
        );

    \I__8004\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32589\
        );

    \I__8003\ : CascadeMux
    port map (
            O => \N__32594\,
            I => \N__32585\
        );

    \I__8002\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32582\
        );

    \I__8001\ : CascadeMux
    port map (
            O => \N__32592\,
            I => \N__32579\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__32589\,
            I => \N__32575\
        );

    \I__7999\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32572\
        );

    \I__7998\ : InMux
    port map (
            O => \N__32585\,
            I => \N__32569\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__32582\,
            I => \N__32565\
        );

    \I__7996\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32562\
        );

    \I__7995\ : InMux
    port map (
            O => \N__32578\,
            I => \N__32559\
        );

    \I__7994\ : Span4Mux_v
    port map (
            O => \N__32575\,
            I => \N__32556\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__32572\,
            I => \N__32551\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__32569\,
            I => \N__32551\
        );

    \I__7991\ : CascadeMux
    port map (
            O => \N__32568\,
            I => \N__32548\
        );

    \I__7990\ : Span4Mux_v
    port map (
            O => \N__32565\,
            I => \N__32544\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__32562\,
            I => \N__32538\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__32559\,
            I => \N__32538\
        );

    \I__7987\ : Span4Mux_v
    port map (
            O => \N__32556\,
            I => \N__32533\
        );

    \I__7986\ : Span4Mux_v
    port map (
            O => \N__32551\,
            I => \N__32533\
        );

    \I__7985\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32530\
        );

    \I__7984\ : CascadeMux
    port map (
            O => \N__32547\,
            I => \N__32526\
        );

    \I__7983\ : Span4Mux_v
    port map (
            O => \N__32544\,
            I => \N__32523\
        );

    \I__7982\ : InMux
    port map (
            O => \N__32543\,
            I => \N__32520\
        );

    \I__7981\ : Span4Mux_v
    port map (
            O => \N__32538\,
            I => \N__32513\
        );

    \I__7980\ : Span4Mux_h
    port map (
            O => \N__32533\,
            I => \N__32513\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__32530\,
            I => \N__32513\
        );

    \I__7978\ : InMux
    port map (
            O => \N__32529\,
            I => \N__32510\
        );

    \I__7977\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32507\
        );

    \I__7976\ : Sp12to4
    port map (
            O => \N__32523\,
            I => \N__32502\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__32520\,
            I => \N__32502\
        );

    \I__7974\ : Sp12to4
    port map (
            O => \N__32513\,
            I => \N__32499\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__32510\,
            I => \N__32494\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__32507\,
            I => \N__32494\
        );

    \I__7971\ : Span12Mux_h
    port map (
            O => \N__32502\,
            I => \N__32489\
        );

    \I__7970\ : Span12Mux_v
    port map (
            O => \N__32499\,
            I => \N__32489\
        );

    \I__7969\ : Span12Mux_v
    port map (
            O => \N__32494\,
            I => \N__32486\
        );

    \I__7968\ : Odrv12
    port map (
            O => \N__32489\,
            I => port_data_c_4
        );

    \I__7967\ : Odrv12
    port map (
            O => \N__32486\,
            I => port_data_c_4
        );

    \I__7966\ : IoInMux
    port map (
            O => \N__32481\,
            I => \N__32477\
        );

    \I__7965\ : InMux
    port map (
            O => \N__32480\,
            I => \N__32474\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__32477\,
            I => \N__32471\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__32474\,
            I => \N__32468\
        );

    \I__7962\ : Span12Mux_s6_h
    port map (
            O => \N__32471\,
            I => \N__32465\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__32468\,
            I => \N__32462\
        );

    \I__7960\ : Odrv12
    port map (
            O => \N__32465\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__7959\ : Odrv4
    port map (
            O => \N__32462\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__7958\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32454\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__32454\,
            I => \N__32451\
        );

    \I__7956\ : Span4Mux_h
    port map (
            O => \N__32451\,
            I => \N__32448\
        );

    \I__7955\ : Odrv4
    port map (
            O => \N__32448\,
            I => \un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0\
        );

    \I__7954\ : IoInMux
    port map (
            O => \N__32445\,
            I => \N__32441\
        );

    \I__7953\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32438\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__32441\,
            I => \N__32435\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__32438\,
            I => \N__32432\
        );

    \I__7950\ : Span12Mux_s6_h
    port map (
            O => \N__32435\,
            I => \N__32429\
        );

    \I__7949\ : Span4Mux_h
    port map (
            O => \N__32432\,
            I => \N__32426\
        );

    \I__7948\ : Odrv12
    port map (
            O => \N__32429\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__32426\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__7946\ : InMux
    port map (
            O => \N__32421\,
            I => \N__32418\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32415\
        );

    \I__7944\ : Span4Mux_h
    port map (
            O => \N__32415\,
            I => \N__32412\
        );

    \I__7943\ : Odrv4
    port map (
            O => \N__32412\,
            I => \un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0\
        );

    \I__7942\ : CascadeMux
    port map (
            O => \N__32409\,
            I => \N__32404\
        );

    \I__7941\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32400\
        );

    \I__7940\ : CascadeMux
    port map (
            O => \N__32407\,
            I => \N__32397\
        );

    \I__7939\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32394\
        );

    \I__7938\ : CascadeMux
    port map (
            O => \N__32403\,
            I => \N__32390\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__32400\,
            I => \N__32385\
        );

    \I__7936\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32382\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__32394\,
            I => \N__32379\
        );

    \I__7934\ : InMux
    port map (
            O => \N__32393\,
            I => \N__32374\
        );

    \I__7933\ : InMux
    port map (
            O => \N__32390\,
            I => \N__32374\
        );

    \I__7932\ : CascadeMux
    port map (
            O => \N__32389\,
            I => \N__32371\
        );

    \I__7931\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32368\
        );

    \I__7930\ : Span4Mux_v
    port map (
            O => \N__32385\,
            I => \N__32365\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__32382\,
            I => \N__32362\
        );

    \I__7928\ : Span4Mux_h
    port map (
            O => \N__32379\,
            I => \N__32359\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__32374\,
            I => \N__32356\
        );

    \I__7926\ : InMux
    port map (
            O => \N__32371\,
            I => \N__32353\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__32368\,
            I => \N__32349\
        );

    \I__7924\ : Sp12to4
    port map (
            O => \N__32365\,
            I => \N__32345\
        );

    \I__7923\ : Span4Mux_v
    port map (
            O => \N__32362\,
            I => \N__32342\
        );

    \I__7922\ : Span4Mux_v
    port map (
            O => \N__32359\,
            I => \N__32335\
        );

    \I__7921\ : Span4Mux_h
    port map (
            O => \N__32356\,
            I => \N__32335\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__32353\,
            I => \N__32335\
        );

    \I__7919\ : CascadeMux
    port map (
            O => \N__32352\,
            I => \N__32332\
        );

    \I__7918\ : Span4Mux_h
    port map (
            O => \N__32349\,
            I => \N__32328\
        );

    \I__7917\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32325\
        );

    \I__7916\ : Span12Mux_h
    port map (
            O => \N__32345\,
            I => \N__32322\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__32342\,
            I => \N__32319\
        );

    \I__7914\ : Span4Mux_h
    port map (
            O => \N__32335\,
            I => \N__32316\
        );

    \I__7913\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32313\
        );

    \I__7912\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32310\
        );

    \I__7911\ : Span4Mux_v
    port map (
            O => \N__32328\,
            I => \N__32305\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__32325\,
            I => \N__32305\
        );

    \I__7909\ : Span12Mux_h
    port map (
            O => \N__32322\,
            I => \N__32302\
        );

    \I__7908\ : Span4Mux_v
    port map (
            O => \N__32319\,
            I => \N__32299\
        );

    \I__7907\ : Sp12to4
    port map (
            O => \N__32316\,
            I => \N__32290\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__32313\,
            I => \N__32290\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__32310\,
            I => \N__32290\
        );

    \I__7904\ : Sp12to4
    port map (
            O => \N__32305\,
            I => \N__32290\
        );

    \I__7903\ : Span12Mux_v
    port map (
            O => \N__32302\,
            I => \N__32287\
        );

    \I__7902\ : Sp12to4
    port map (
            O => \N__32299\,
            I => \N__32282\
        );

    \I__7901\ : Span12Mux_v
    port map (
            O => \N__32290\,
            I => \N__32282\
        );

    \I__7900\ : Odrv12
    port map (
            O => \N__32287\,
            I => port_data_c_6
        );

    \I__7899\ : Odrv12
    port map (
            O => \N__32282\,
            I => port_data_c_6
        );

    \I__7898\ : IoInMux
    port map (
            O => \N__32277\,
            I => \N__32274\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__32274\,
            I => \N__32271\
        );

    \I__7896\ : IoSpan4Mux
    port map (
            O => \N__32271\,
            I => \N__32267\
        );

    \I__7895\ : InMux
    port map (
            O => \N__32270\,
            I => \N__32264\
        );

    \I__7894\ : Span4Mux_s2_h
    port map (
            O => \N__32267\,
            I => \N__32261\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__32264\,
            I => \N__32258\
        );

    \I__7892\ : Span4Mux_v
    port map (
            O => \N__32261\,
            I => \N__32255\
        );

    \I__7891\ : Span4Mux_v
    port map (
            O => \N__32258\,
            I => \N__32252\
        );

    \I__7890\ : Odrv4
    port map (
            O => \N__32255\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__7889\ : Odrv4
    port map (
            O => \N__32252\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__7888\ : InMux
    port map (
            O => \N__32247\,
            I => \N__32244\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__32244\,
            I => \N_63_0\
        );

    \I__7886\ : InMux
    port map (
            O => \N__32241\,
            I => \N__32238\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__32238\,
            I => \N_75_0\
        );

    \I__7884\ : InMux
    port map (
            O => \N__32235\,
            I => \N__32232\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__32232\,
            I => \M_this_oam_ram_write_data_11\
        );

    \I__7882\ : CascadeMux
    port map (
            O => \N__32229\,
            I => \N__32226\
        );

    \I__7881\ : InMux
    port map (
            O => \N__32226\,
            I => \N__32223\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__32223\,
            I => \M_this_data_tmp_qZ0Z_11\
        );

    \I__7879\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32217\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__32217\,
            I => \N__32214\
        );

    \I__7877\ : Odrv4
    port map (
            O => \N__32214\,
            I => \M_this_data_tmp_qZ0Z_12\
        );

    \I__7876\ : CascadeMux
    port map (
            O => \N__32211\,
            I => \N__32208\
        );

    \I__7875\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32205\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__32205\,
            I => \M_this_data_tmp_qZ0Z_9\
        );

    \I__7873\ : CascadeMux
    port map (
            O => \N__32202\,
            I => \N__32199\
        );

    \I__7872\ : InMux
    port map (
            O => \N__32199\,
            I => \N__32196\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__32196\,
            I => \N__32193\
        );

    \I__7870\ : Odrv4
    port map (
            O => \N__32193\,
            I => \M_this_data_tmp_qZ0Z_14\
        );

    \I__7869\ : CEMux
    port map (
            O => \N__32190\,
            I => \N__32185\
        );

    \I__7868\ : CEMux
    port map (
            O => \N__32189\,
            I => \N__32180\
        );

    \I__7867\ : CEMux
    port map (
            O => \N__32188\,
            I => \N__32177\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__32185\,
            I => \N__32174\
        );

    \I__7865\ : CEMux
    port map (
            O => \N__32184\,
            I => \N__32171\
        );

    \I__7864\ : CEMux
    port map (
            O => \N__32183\,
            I => \N__32168\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__32180\,
            I => \N__32165\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__32177\,
            I => \N__32162\
        );

    \I__7861\ : Span4Mux_v
    port map (
            O => \N__32174\,
            I => \N__32159\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__32171\,
            I => \N__32156\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__32168\,
            I => \N__32153\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__32165\,
            I => \N__32150\
        );

    \I__7857\ : Span4Mux_v
    port map (
            O => \N__32162\,
            I => \N__32143\
        );

    \I__7856\ : Span4Mux_h
    port map (
            O => \N__32159\,
            I => \N__32143\
        );

    \I__7855\ : Span4Mux_v
    port map (
            O => \N__32156\,
            I => \N__32143\
        );

    \I__7854\ : Span4Mux_h
    port map (
            O => \N__32153\,
            I => \N__32140\
        );

    \I__7853\ : Sp12to4
    port map (
            O => \N__32150\,
            I => \N__32137\
        );

    \I__7852\ : Span4Mux_h
    port map (
            O => \N__32143\,
            I => \N__32134\
        );

    \I__7851\ : Odrv4
    port map (
            O => \N__32140\,
            I => \N_1134_0\
        );

    \I__7850\ : Odrv12
    port map (
            O => \N__32137\,
            I => \N_1134_0\
        );

    \I__7849\ : Odrv4
    port map (
            O => \N__32134\,
            I => \N_1134_0\
        );

    \I__7848\ : InMux
    port map (
            O => \N__32127\,
            I => \N__32124\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__32124\,
            I => \N_39_0\
        );

    \I__7846\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32118\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__32118\,
            I => \M_this_oam_ram_write_data_27\
        );

    \I__7844\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32112\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__32112\,
            I => \M_this_oam_ram_write_data_8\
        );

    \I__7842\ : CascadeMux
    port map (
            O => \N__32109\,
            I => \N__32106\
        );

    \I__7841\ : InMux
    port map (
            O => \N__32106\,
            I => \N__32103\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__32103\,
            I => \M_this_data_tmp_qZ0Z_8\
        );

    \I__7839\ : InMux
    port map (
            O => \N__32100\,
            I => \N__32097\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__32097\,
            I => \N_79_0\
        );

    \I__7837\ : CascadeMux
    port map (
            O => \N__32094\,
            I => \N__32091\
        );

    \I__7836\ : InMux
    port map (
            O => \N__32091\,
            I => \N__32088\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__32088\,
            I => \M_this_data_tmp_qZ0Z_0\
        );

    \I__7834\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32082\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__32082\,
            I => \N__32079\
        );

    \I__7832\ : Span4Mux_v
    port map (
            O => \N__32079\,
            I => \N__32076\
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__32076\,
            I => \N_43_0\
        );

    \I__7830\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32070\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__32070\,
            I => \N__32067\
        );

    \I__7828\ : Odrv4
    port map (
            O => \N__32067\,
            I => \N_77_0\
        );

    \I__7827\ : InMux
    port map (
            O => \N__32064\,
            I => \N__32061\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__32061\,
            I => \M_this_data_tmp_qZ0Z_1\
        );

    \I__7825\ : InMux
    port map (
            O => \N__32058\,
            I => \N__32055\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__32055\,
            I => \N_58_0\
        );

    \I__7823\ : InMux
    port map (
            O => \N__32052\,
            I => \N__32049\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__32049\,
            I => \M_this_oam_ram_write_data_14\
        );

    \I__7821\ : InMux
    port map (
            O => \N__32046\,
            I => \bfn_24_23_0_\
        );

    \I__7820\ : IoInMux
    port map (
            O => \N__32043\,
            I => \N__32040\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__32040\,
            I => \N__32037\
        );

    \I__7818\ : Span4Mux_s1_v
    port map (
            O => \N__32037\,
            I => \N__32034\
        );

    \I__7817\ : Span4Mux_v
    port map (
            O => \N__32034\,
            I => \N__32030\
        );

    \I__7816\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32027\
        );

    \I__7815\ : Span4Mux_v
    port map (
            O => \N__32030\,
            I => \N__32022\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__32027\,
            I => \N__32022\
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__32022\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__7812\ : InMux
    port map (
            O => \N__32019\,
            I => \N__32016\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__32016\,
            I => \N__32013\
        );

    \I__7810\ : Odrv12
    port map (
            O => \N__32013\,
            I => \un1_M_this_external_address_q_cry_8_c_RNI09PBZ0\
        );

    \I__7809\ : InMux
    port map (
            O => \N__32010\,
            I => \un1_M_this_external_address_q_cry_8\
        );

    \I__7808\ : InMux
    port map (
            O => \N__32007\,
            I => \un1_M_this_external_address_q_cry_9\
        );

    \I__7807\ : InMux
    port map (
            O => \N__32004\,
            I => \un1_M_this_external_address_q_cry_10\
        );

    \I__7806\ : InMux
    port map (
            O => \N__32001\,
            I => \un1_M_this_external_address_q_cry_11\
        );

    \I__7805\ : InMux
    port map (
            O => \N__31998\,
            I => \un1_M_this_external_address_q_cry_12\
        );

    \I__7804\ : InMux
    port map (
            O => \N__31995\,
            I => \un1_M_this_external_address_q_cry_13\
        );

    \I__7803\ : InMux
    port map (
            O => \N__31992\,
            I => \un1_M_this_external_address_q_cry_14\
        );

    \I__7802\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31985\
        );

    \I__7801\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31980\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__31985\,
            I => \N__31977\
        );

    \I__7799\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31974\
        );

    \I__7798\ : InMux
    port map (
            O => \N__31983\,
            I => \N__31971\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__31980\,
            I => \N__31964\
        );

    \I__7796\ : Span4Mux_v
    port map (
            O => \N__31977\,
            I => \N__31961\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__31974\,
            I => \N__31958\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__31971\,
            I => \N__31955\
        );

    \I__7793\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31952\
        );

    \I__7792\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31949\
        );

    \I__7791\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31944\
        );

    \I__7790\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31941\
        );

    \I__7789\ : Span4Mux_v
    port map (
            O => \N__31964\,
            I => \N__31937\
        );

    \I__7788\ : Span4Mux_v
    port map (
            O => \N__31961\,
            I => \N__31932\
        );

    \I__7787\ : Span4Mux_v
    port map (
            O => \N__31958\,
            I => \N__31932\
        );

    \I__7786\ : Span4Mux_v
    port map (
            O => \N__31955\,
            I => \N__31929\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__31952\,
            I => \N__31924\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__31949\,
            I => \N__31924\
        );

    \I__7783\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31921\
        );

    \I__7782\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31918\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__31944\,
            I => \N__31915\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__31941\,
            I => \N__31912\
        );

    \I__7779\ : InMux
    port map (
            O => \N__31940\,
            I => \N__31909\
        );

    \I__7778\ : Odrv4
    port map (
            O => \N__31937\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7777\ : Odrv4
    port map (
            O => \N__31932\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__31929\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7775\ : Odrv12
    port map (
            O => \N__31924\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__31921\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__31918\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7772\ : Odrv4
    port map (
            O => \N__31915\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7771\ : Odrv4
    port map (
            O => \N__31912\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__31909\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7769\ : InMux
    port map (
            O => \N__31890\,
            I => \N__31887\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__31887\,
            I => \N__31882\
        );

    \I__7767\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31879\
        );

    \I__7766\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31876\
        );

    \I__7765\ : Span4Mux_v
    port map (
            O => \N__31882\,
            I => \N__31870\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__31879\,
            I => \N__31870\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__31876\,
            I => \N__31867\
        );

    \I__7762\ : InMux
    port map (
            O => \N__31875\,
            I => \N__31864\
        );

    \I__7761\ : Span4Mux_h
    port map (
            O => \N__31870\,
            I => \N__31858\
        );

    \I__7760\ : Span4Mux_h
    port map (
            O => \N__31867\,
            I => \N__31853\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__31864\,
            I => \N__31853\
        );

    \I__7758\ : InMux
    port map (
            O => \N__31863\,
            I => \N__31850\
        );

    \I__7757\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31847\
        );

    \I__7756\ : CascadeMux
    port map (
            O => \N__31861\,
            I => \N__31840\
        );

    \I__7755\ : Span4Mux_v
    port map (
            O => \N__31858\,
            I => \N__31835\
        );

    \I__7754\ : Span4Mux_h
    port map (
            O => \N__31853\,
            I => \N__31835\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__31850\,
            I => \N__31830\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__31847\,
            I => \N__31830\
        );

    \I__7751\ : InMux
    port map (
            O => \N__31846\,
            I => \N__31827\
        );

    \I__7750\ : InMux
    port map (
            O => \N__31845\,
            I => \N__31824\
        );

    \I__7749\ : InMux
    port map (
            O => \N__31844\,
            I => \N__31821\
        );

    \I__7748\ : InMux
    port map (
            O => \N__31843\,
            I => \N__31818\
        );

    \I__7747\ : InMux
    port map (
            O => \N__31840\,
            I => \N__31815\
        );

    \I__7746\ : Odrv4
    port map (
            O => \N__31835\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7745\ : Odrv12
    port map (
            O => \N__31830\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__31827\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__31824\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__31821\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__31818\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__31815\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7739\ : CascadeMux
    port map (
            O => \N__31800\,
            I => \N__31796\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__31799\,
            I => \N__31792\
        );

    \I__7737\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31787\
        );

    \I__7736\ : CascadeMux
    port map (
            O => \N__31795\,
            I => \N__31784\
        );

    \I__7735\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31780\
        );

    \I__7734\ : CascadeMux
    port map (
            O => \N__31791\,
            I => \N__31776\
        );

    \I__7733\ : CascadeMux
    port map (
            O => \N__31790\,
            I => \N__31773\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__31787\,
            I => \N__31770\
        );

    \I__7731\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31767\
        );

    \I__7730\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31764\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__31780\,
            I => \N__31761\
        );

    \I__7728\ : CascadeMux
    port map (
            O => \N__31779\,
            I => \N__31758\
        );

    \I__7727\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31755\
        );

    \I__7726\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31750\
        );

    \I__7725\ : Span4Mux_v
    port map (
            O => \N__31770\,
            I => \N__31746\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__31767\,
            I => \N__31743\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__31764\,
            I => \N__31740\
        );

    \I__7722\ : Span4Mux_v
    port map (
            O => \N__31761\,
            I => \N__31737\
        );

    \I__7721\ : InMux
    port map (
            O => \N__31758\,
            I => \N__31734\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__31755\,
            I => \N__31731\
        );

    \I__7719\ : CascadeMux
    port map (
            O => \N__31754\,
            I => \N__31728\
        );

    \I__7718\ : CascadeMux
    port map (
            O => \N__31753\,
            I => \N__31725\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__31750\,
            I => \N__31721\
        );

    \I__7716\ : InMux
    port map (
            O => \N__31749\,
            I => \N__31718\
        );

    \I__7715\ : Span4Mux_v
    port map (
            O => \N__31746\,
            I => \N__31711\
        );

    \I__7714\ : Span4Mux_v
    port map (
            O => \N__31743\,
            I => \N__31711\
        );

    \I__7713\ : Span4Mux_h
    port map (
            O => \N__31740\,
            I => \N__31711\
        );

    \I__7712\ : Span4Mux_v
    port map (
            O => \N__31737\,
            I => \N__31708\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__31734\,
            I => \N__31705\
        );

    \I__7710\ : Span4Mux_v
    port map (
            O => \N__31731\,
            I => \N__31702\
        );

    \I__7709\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31699\
        );

    \I__7708\ : InMux
    port map (
            O => \N__31725\,
            I => \N__31696\
        );

    \I__7707\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31693\
        );

    \I__7706\ : Span4Mux_v
    port map (
            O => \N__31721\,
            I => \N__31686\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__31718\,
            I => \N__31686\
        );

    \I__7704\ : Span4Mux_h
    port map (
            O => \N__31711\,
            I => \N__31686\
        );

    \I__7703\ : Odrv4
    port map (
            O => \N__31708\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7702\ : Odrv12
    port map (
            O => \N__31705\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7701\ : Odrv4
    port map (
            O => \N__31702\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__31699\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__31696\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__31693\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__31686\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7696\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31668\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__31668\,
            I => \N__31664\
        );

    \I__7694\ : InMux
    port map (
            O => \N__31667\,
            I => \N__31661\
        );

    \I__7693\ : Span4Mux_v
    port map (
            O => \N__31664\,
            I => \N__31656\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__31661\,
            I => \N__31653\
        );

    \I__7691\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31650\
        );

    \I__7690\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31646\
        );

    \I__7689\ : Span4Mux_v
    port map (
            O => \N__31656\,
            I => \N__31640\
        );

    \I__7688\ : Span4Mux_v
    port map (
            O => \N__31653\,
            I => \N__31640\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__31650\,
            I => \N__31637\
        );

    \I__7686\ : InMux
    port map (
            O => \N__31649\,
            I => \N__31634\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__31646\,
            I => \N__31631\
        );

    \I__7684\ : InMux
    port map (
            O => \N__31645\,
            I => \N__31628\
        );

    \I__7683\ : Span4Mux_h
    port map (
            O => \N__31640\,
            I => \N__31621\
        );

    \I__7682\ : Span4Mux_v
    port map (
            O => \N__31637\,
            I => \N__31621\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__31634\,
            I => \N__31618\
        );

    \I__7680\ : Span4Mux_v
    port map (
            O => \N__31631\,
            I => \N__31615\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__31628\,
            I => \N__31612\
        );

    \I__7678\ : InMux
    port map (
            O => \N__31627\,
            I => \N__31609\
        );

    \I__7677\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31606\
        );

    \I__7676\ : Odrv4
    port map (
            O => \N__31621\,
            I => \M_this_sprites_ram_write_en_0_0\
        );

    \I__7675\ : Odrv12
    port map (
            O => \N__31618\,
            I => \M_this_sprites_ram_write_en_0_0\
        );

    \I__7674\ : Odrv4
    port map (
            O => \N__31615\,
            I => \M_this_sprites_ram_write_en_0_0\
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__31612\,
            I => \M_this_sprites_ram_write_en_0_0\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__31609\,
            I => \M_this_sprites_ram_write_en_0_0\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__31606\,
            I => \M_this_sprites_ram_write_en_0_0\
        );

    \I__7670\ : CEMux
    port map (
            O => \N__31593\,
            I => \N__31589\
        );

    \I__7669\ : CEMux
    port map (
            O => \N__31592\,
            I => \N__31586\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__31589\,
            I => \N__31581\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__31586\,
            I => \N__31581\
        );

    \I__7666\ : Odrv4
    port map (
            O => \N__31581\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__7665\ : InMux
    port map (
            O => \N__31578\,
            I => \N__31575\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__31575\,
            I => \N__31572\
        );

    \I__7663\ : Span4Mux_v
    port map (
            O => \N__31572\,
            I => \N__31569\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__31569\,
            I => \M_this_oam_ram_write_data_30\
        );

    \I__7661\ : InMux
    port map (
            O => \N__31566\,
            I => \un1_M_this_external_address_q_cry_0\
        );

    \I__7660\ : InMux
    port map (
            O => \N__31563\,
            I => \un1_M_this_external_address_q_cry_1\
        );

    \I__7659\ : InMux
    port map (
            O => \N__31560\,
            I => \un1_M_this_external_address_q_cry_2\
        );

    \I__7658\ : InMux
    port map (
            O => \N__31557\,
            I => \un1_M_this_external_address_q_cry_3\
        );

    \I__7657\ : InMux
    port map (
            O => \N__31554\,
            I => \un1_M_this_external_address_q_cry_4\
        );

    \I__7656\ : InMux
    port map (
            O => \N__31551\,
            I => \un1_M_this_external_address_q_cry_5\
        );

    \I__7655\ : InMux
    port map (
            O => \N__31548\,
            I => \un1_M_this_external_address_q_cry_6\
        );

    \I__7654\ : InMux
    port map (
            O => \N__31545\,
            I => \N__31542\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__31542\,
            I => \N__31537\
        );

    \I__7652\ : InMux
    port map (
            O => \N__31541\,
            I => \N__31529\
        );

    \I__7651\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31529\
        );

    \I__7650\ : Span4Mux_h
    port map (
            O => \N__31537\,
            I => \N__31526\
        );

    \I__7649\ : InMux
    port map (
            O => \N__31536\,
            I => \N__31519\
        );

    \I__7648\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31519\
        );

    \I__7647\ : InMux
    port map (
            O => \N__31534\,
            I => \N__31519\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31516\
        );

    \I__7645\ : Odrv4
    port map (
            O => \N__31526\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__31519\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__31516\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__7642\ : CascadeMux
    port map (
            O => \N__31509\,
            I => \N__31506\
        );

    \I__7641\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31503\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__31503\,
            I => \N__31500\
        );

    \I__7639\ : Span4Mux_v
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__7638\ : Odrv4
    port map (
            O => \N__31497\,
            I => \M_this_oam_ram_read_data_i_19\
        );

    \I__7637\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31491\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__31491\,
            I => \M_this_data_tmp_qZ0Z_16\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__31488\,
            I => \N__31485\
        );

    \I__7634\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31482\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__31482\,
            I => \M_this_data_tmp_qZ0Z_19\
        );

    \I__7632\ : CascadeMux
    port map (
            O => \N__31479\,
            I => \N__31476\
        );

    \I__7631\ : InMux
    port map (
            O => \N__31476\,
            I => \N__31473\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__31473\,
            I => \M_this_data_tmp_qZ0Z_18\
        );

    \I__7629\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31467\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__31467\,
            I => \M_this_data_tmp_qZ0Z_22\
        );

    \I__7627\ : CascadeMux
    port map (
            O => \N__31464\,
            I => \N__31461\
        );

    \I__7626\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31458\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__31458\,
            I => \M_this_data_tmp_qZ0Z_17\
        );

    \I__7624\ : InMux
    port map (
            O => \N__31455\,
            I => \N__31452\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__31452\,
            I => \N_54_0\
        );

    \I__7622\ : CEMux
    port map (
            O => \N__31449\,
            I => \N__31446\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__31446\,
            I => \N__31442\
        );

    \I__7620\ : CEMux
    port map (
            O => \N__31445\,
            I => \N__31439\
        );

    \I__7619\ : Span4Mux_v
    port map (
            O => \N__31442\,
            I => \N__31433\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__31439\,
            I => \N__31433\
        );

    \I__7617\ : CEMux
    port map (
            O => \N__31438\,
            I => \N__31430\
        );

    \I__7616\ : Span4Mux_h
    port map (
            O => \N__31433\,
            I => \N__31427\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__31430\,
            I => \N__31424\
        );

    \I__7614\ : Span4Mux_h
    port map (
            O => \N__31427\,
            I => \N__31421\
        );

    \I__7613\ : Odrv12
    port map (
            O => \N__31424\,
            I => \N_1126_0\
        );

    \I__7612\ : Odrv4
    port map (
            O => \N__31421\,
            I => \N_1126_0\
        );

    \I__7611\ : CascadeMux
    port map (
            O => \N__31416\,
            I => \N__31412\
        );

    \I__7610\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31409\
        );

    \I__7609\ : InMux
    port map (
            O => \N__31412\,
            I => \N__31406\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__31409\,
            I => \N__31401\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__31406\,
            I => \N__31401\
        );

    \I__7606\ : Span4Mux_v
    port map (
            O => \N__31401\,
            I => \N__31398\
        );

    \I__7605\ : Odrv4
    port map (
            O => \N__31398\,
            I => \M_this_oam_ram_read_data_23\
        );

    \I__7604\ : CascadeMux
    port map (
            O => \N__31395\,
            I => \this_ppu.un1_oam_data_c2_cascade_\
        );

    \I__7603\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31389\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__31389\,
            I => \N__31386\
        );

    \I__7601\ : Span4Mux_h
    port map (
            O => \N__31386\,
            I => \N__31383\
        );

    \I__7600\ : Odrv4
    port map (
            O => \N__31383\,
            I => \this_ppu.un1_M_vaddress_q_3_7\
        );

    \I__7599\ : InMux
    port map (
            O => \N__31380\,
            I => \N__31377\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__31377\,
            I => \M_this_oam_ram_write_data_22\
        );

    \I__7597\ : InMux
    port map (
            O => \N__31374\,
            I => \N__31369\
        );

    \I__7596\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31366\
        );

    \I__7595\ : CascadeMux
    port map (
            O => \N__31372\,
            I => \N__31363\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__31369\,
            I => \N__31358\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__31366\,
            I => \N__31358\
        );

    \I__7592\ : InMux
    port map (
            O => \N__31363\,
            I => \N__31355\
        );

    \I__7591\ : Span4Mux_v
    port map (
            O => \N__31358\,
            I => \N__31352\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__31355\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__7589\ : Odrv4
    port map (
            O => \N__31352\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__31347\,
            I => \N__31344\
        );

    \I__7587\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31341\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__31341\,
            I => \N__31338\
        );

    \I__7585\ : Span4Mux_h
    port map (
            O => \N__31338\,
            I => \N__31335\
        );

    \I__7584\ : Odrv4
    port map (
            O => \N__31335\,
            I => \this_ppu.un1_M_vaddress_q_3_6\
        );

    \I__7583\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31329\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__31329\,
            I => \M_this_oam_ram_write_data_31\
        );

    \I__7581\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31323\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__31323\,
            I => \N_52_0\
        );

    \I__7579\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31317\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__31317\,
            I => \M_this_oam_ram_write_data_16\
        );

    \I__7577\ : CEMux
    port map (
            O => \N__31314\,
            I => \N__31311\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__31311\,
            I => \N__31307\
        );

    \I__7575\ : CEMux
    port map (
            O => \N__31310\,
            I => \N__31304\
        );

    \I__7574\ : Span4Mux_h
    port map (
            O => \N__31307\,
            I => \N__31299\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__31304\,
            I => \N__31299\
        );

    \I__7572\ : Span4Mux_v
    port map (
            O => \N__31299\,
            I => \N__31296\
        );

    \I__7571\ : Span4Mux_v
    port map (
            O => \N__31296\,
            I => \N__31293\
        );

    \I__7570\ : Odrv4
    port map (
            O => \N__31293\,
            I => \N_158_0\
        );

    \I__7569\ : InMux
    port map (
            O => \N__31290\,
            I => \N__31286\
        );

    \I__7568\ : InMux
    port map (
            O => \N__31289\,
            I => \N__31283\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__31286\,
            I => \N__31279\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__31283\,
            I => \N__31275\
        );

    \I__7565\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31272\
        );

    \I__7564\ : Span4Mux_h
    port map (
            O => \N__31279\,
            I => \N__31269\
        );

    \I__7563\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31266\
        );

    \I__7562\ : Odrv4
    port map (
            O => \N__31275\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__31272\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__31269\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__31266\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__7558\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31253\
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__31256\,
            I => \N__31250\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__31253\,
            I => \N__31244\
        );

    \I__7555\ : InMux
    port map (
            O => \N__31250\,
            I => \N__31239\
        );

    \I__7554\ : InMux
    port map (
            O => \N__31249\,
            I => \N__31239\
        );

    \I__7553\ : InMux
    port map (
            O => \N__31248\,
            I => \N__31234\
        );

    \I__7552\ : InMux
    port map (
            O => \N__31247\,
            I => \N__31234\
        );

    \I__7551\ : Span4Mux_h
    port map (
            O => \N__31244\,
            I => \N__31231\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__31239\,
            I => \N__31228\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__31234\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__31231\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__7547\ : Odrv4
    port map (
            O => \N__31228\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__7546\ : CascadeMux
    port map (
            O => \N__31221\,
            I => \N__31218\
        );

    \I__7545\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31215\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__31215\,
            I => \N__31212\
        );

    \I__7543\ : Span4Mux_h
    port map (
            O => \N__31212\,
            I => \N__31209\
        );

    \I__7542\ : Odrv4
    port map (
            O => \N__31209\,
            I => \this_ppu.un1_M_vaddress_q_3_5\
        );

    \I__7541\ : CascadeMux
    port map (
            O => \N__31206\,
            I => \N__31202\
        );

    \I__7540\ : CascadeMux
    port map (
            O => \N__31205\,
            I => \N__31198\
        );

    \I__7539\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31195\
        );

    \I__7538\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31192\
        );

    \I__7537\ : InMux
    port map (
            O => \N__31198\,
            I => \N__31189\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__31195\,
            I => \N__31186\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__31192\,
            I => \N__31183\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__31189\,
            I => \N__31180\
        );

    \I__7533\ : Span4Mux_h
    port map (
            O => \N__31186\,
            I => \N__31177\
        );

    \I__7532\ : Span4Mux_v
    port map (
            O => \N__31183\,
            I => \N__31172\
        );

    \I__7531\ : Span4Mux_h
    port map (
            O => \N__31180\,
            I => \N__31172\
        );

    \I__7530\ : Odrv4
    port map (
            O => \N__31177\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__7529\ : Odrv4
    port map (
            O => \N__31172\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__7528\ : InMux
    port map (
            O => \N__31167\,
            I => \N__31164\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__31164\,
            I => \M_this_oam_ram_read_data_i_17\
        );

    \I__7526\ : InMux
    port map (
            O => \N__31161\,
            I => \N__31158\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__31158\,
            I => \N__31155\
        );

    \I__7524\ : Span4Mux_h
    port map (
            O => \N__31155\,
            I => \N__31152\
        );

    \I__7523\ : Span4Mux_h
    port map (
            O => \N__31152\,
            I => \N__31149\
        );

    \I__7522\ : Span4Mux_h
    port map (
            O => \N__31149\,
            I => \N__31145\
        );

    \I__7521\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31142\
        );

    \I__7520\ : Odrv4
    port map (
            O => \N__31145\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__31142\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__7518\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__7516\ : Span4Mux_v
    port map (
            O => \N__31131\,
            I => \N__31128\
        );

    \I__7515\ : Sp12to4
    port map (
            O => \N__31128\,
            I => \N__31124\
        );

    \I__7514\ : InMux
    port map (
            O => \N__31127\,
            I => \N__31121\
        );

    \I__7513\ : Odrv12
    port map (
            O => \N__31124\,
            I => \M_this_oam_ram_read_data_1\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__31121\,
            I => \M_this_oam_ram_read_data_1\
        );

    \I__7511\ : InMux
    port map (
            O => \N__31116\,
            I => \N__31113\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__31113\,
            I => \N__31110\
        );

    \I__7509\ : Span4Mux_v
    port map (
            O => \N__31110\,
            I => \N__31106\
        );

    \I__7508\ : CascadeMux
    port map (
            O => \N__31109\,
            I => \N__31103\
        );

    \I__7507\ : Span4Mux_h
    port map (
            O => \N__31106\,
            I => \N__31100\
        );

    \I__7506\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31097\
        );

    \I__7505\ : Span4Mux_h
    port map (
            O => \N__31100\,
            I => \N__31094\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__31097\,
            I => \M_this_oam_ram_read_data_0\
        );

    \I__7503\ : Odrv4
    port map (
            O => \N__31094\,
            I => \M_this_oam_ram_read_data_0\
        );

    \I__7502\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31086\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__31086\,
            I => \N__31083\
        );

    \I__7500\ : Span12Mux_v
    port map (
            O => \N__31083\,
            I => \N__31080\
        );

    \I__7499\ : Span12Mux_h
    port map (
            O => \N__31080\,
            I => \N__31076\
        );

    \I__7498\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31073\
        );

    \I__7497\ : Odrv12
    port map (
            O => \N__31076\,
            I => \M_this_oam_ram_read_data_3\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__31073\,
            I => \M_this_oam_ram_read_data_3\
        );

    \I__7495\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31065\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__31065\,
            I => \N__31062\
        );

    \I__7493\ : Span4Mux_v
    port map (
            O => \N__31062\,
            I => \N__31059\
        );

    \I__7492\ : Odrv4
    port map (
            O => \N__31059\,
            I => \this_ppu.un9lto7Z0Z_5\
        );

    \I__7491\ : CascadeMux
    port map (
            O => \N__31056\,
            I => \N__31053\
        );

    \I__7490\ : InMux
    port map (
            O => \N__31053\,
            I => \N__31050\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__31050\,
            I => \N__31047\
        );

    \I__7488\ : Span4Mux_h
    port map (
            O => \N__31047\,
            I => \N__31044\
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__31044\,
            I => \this_ppu.un1_M_haddress_q_2_6\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__31041\,
            I => \N__31038\
        );

    \I__7485\ : InMux
    port map (
            O => \N__31038\,
            I => \N__31035\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__31035\,
            I => \N__31032\
        );

    \I__7483\ : Span4Mux_h
    port map (
            O => \N__31032\,
            I => \N__31028\
        );

    \I__7482\ : InMux
    port map (
            O => \N__31031\,
            I => \N__31025\
        );

    \I__7481\ : Odrv4
    port map (
            O => \N__31028\,
            I => \M_this_oam_ram_read_data_4\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__31025\,
            I => \M_this_oam_ram_read_data_4\
        );

    \I__7479\ : InMux
    port map (
            O => \N__31020\,
            I => \N__31017\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__31017\,
            I => \N__31014\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__31014\,
            I => \N__31010\
        );

    \I__7476\ : InMux
    port map (
            O => \N__31013\,
            I => \N__31007\
        );

    \I__7475\ : Odrv4
    port map (
            O => \N__31010\,
            I => \M_this_oam_ram_read_data_6\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__31007\,
            I => \M_this_oam_ram_read_data_6\
        );

    \I__7473\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30999\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__30999\,
            I => \N__30996\
        );

    \I__7471\ : Span4Mux_v
    port map (
            O => \N__30996\,
            I => \N__30992\
        );

    \I__7470\ : CascadeMux
    port map (
            O => \N__30995\,
            I => \N__30989\
        );

    \I__7469\ : Span4Mux_h
    port map (
            O => \N__30992\,
            I => \N__30986\
        );

    \I__7468\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30983\
        );

    \I__7467\ : Odrv4
    port map (
            O => \N__30986\,
            I => \M_this_oam_ram_read_data_7\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__30983\,
            I => \M_this_oam_ram_read_data_7\
        );

    \I__7465\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30975\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__30975\,
            I => \N__30972\
        );

    \I__7463\ : Span4Mux_h
    port map (
            O => \N__30972\,
            I => \N__30969\
        );

    \I__7462\ : Span4Mux_h
    port map (
            O => \N__30969\,
            I => \N__30965\
        );

    \I__7461\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30962\
        );

    \I__7460\ : Odrv4
    port map (
            O => \N__30965\,
            I => \M_this_oam_ram_read_data_5\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__30962\,
            I => \M_this_oam_ram_read_data_5\
        );

    \I__7458\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30954\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__30954\,
            I => \N__30951\
        );

    \I__7456\ : Span4Mux_h
    port map (
            O => \N__30951\,
            I => \N__30948\
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__30948\,
            I => \this_ppu.un9lto7Z0Z_4\
        );

    \I__7454\ : CascadeMux
    port map (
            O => \N__30945\,
            I => \N__30942\
        );

    \I__7453\ : InMux
    port map (
            O => \N__30942\,
            I => \N__30939\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__30939\,
            I => \N__30936\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__30936\,
            I => \N__30933\
        );

    \I__7450\ : Odrv4
    port map (
            O => \N__30933\,
            I => \this_ppu.un1_M_vaddress_q_3_4\
        );

    \I__7449\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30924\
        );

    \I__7448\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30921\
        );

    \I__7447\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30916\
        );

    \I__7446\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30916\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__30924\,
            I => \N__30912\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__30921\,
            I => \N__30909\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30906\
        );

    \I__7442\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30902\
        );

    \I__7441\ : Span4Mux_v
    port map (
            O => \N__30912\,
            I => \N__30899\
        );

    \I__7440\ : Span4Mux_h
    port map (
            O => \N__30909\,
            I => \N__30896\
        );

    \I__7439\ : Span4Mux_h
    port map (
            O => \N__30906\,
            I => \N__30893\
        );

    \I__7438\ : InMux
    port map (
            O => \N__30905\,
            I => \N__30890\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__30902\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7436\ : Odrv4
    port map (
            O => \N__30899\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7435\ : Odrv4
    port map (
            O => \N__30896\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__30893\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__30890\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7432\ : InMux
    port map (
            O => \N__30879\,
            I => \N__30875\
        );

    \I__7431\ : InMux
    port map (
            O => \N__30878\,
            I => \N__30872\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__30875\,
            I => \N__30865\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__30872\,
            I => \N__30865\
        );

    \I__7428\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30862\
        );

    \I__7427\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30858\
        );

    \I__7426\ : Span4Mux_v
    port map (
            O => \N__30865\,
            I => \N__30855\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__30862\,
            I => \N__30852\
        );

    \I__7424\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30849\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__30858\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__7422\ : Odrv4
    port map (
            O => \N__30855\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__7421\ : Odrv12
    port map (
            O => \N__30852\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__30849\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__7419\ : CascadeMux
    port map (
            O => \N__30840\,
            I => \N__30837\
        );

    \I__7418\ : InMux
    port map (
            O => \N__30837\,
            I => \N__30834\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__30834\,
            I => \N__30831\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__30831\,
            I => \N__30827\
        );

    \I__7415\ : InMux
    port map (
            O => \N__30830\,
            I => \N__30824\
        );

    \I__7414\ : Odrv4
    port map (
            O => \N__30827\,
            I => \M_this_oam_ram_read_data_15\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__30824\,
            I => \M_this_oam_ram_read_data_15\
        );

    \I__7412\ : CascadeMux
    port map (
            O => \N__30819\,
            I => \N__30816\
        );

    \I__7411\ : InMux
    port map (
            O => \N__30816\,
            I => \N__30812\
        );

    \I__7410\ : CascadeMux
    port map (
            O => \N__30815\,
            I => \N__30808\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__30812\,
            I => \N__30805\
        );

    \I__7408\ : InMux
    port map (
            O => \N__30811\,
            I => \N__30802\
        );

    \I__7407\ : InMux
    port map (
            O => \N__30808\,
            I => \N__30799\
        );

    \I__7406\ : Span4Mux_h
    port map (
            O => \N__30805\,
            I => \N__30796\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__30802\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__30799\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__7403\ : Odrv4
    port map (
            O => \N__30796\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__7402\ : CascadeMux
    port map (
            O => \N__30789\,
            I => \this_ppu.un1_oam_data_1_c2_cascade_\
        );

    \I__7401\ : CascadeMux
    port map (
            O => \N__30786\,
            I => \N__30783\
        );

    \I__7400\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30779\
        );

    \I__7399\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30776\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30771\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__30776\,
            I => \N__30768\
        );

    \I__7396\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30765\
        );

    \I__7395\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30762\
        );

    \I__7394\ : Span4Mux_v
    port map (
            O => \N__30771\,
            I => \N__30759\
        );

    \I__7393\ : Span4Mux_h
    port map (
            O => \N__30768\,
            I => \N__30756\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__30765\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__30762\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__30759\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__30756\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__7388\ : InMux
    port map (
            O => \N__30747\,
            I => \N__30744\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__30744\,
            I => \N__30741\
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__30741\,
            I => \this_ppu.un1_M_haddress_q_2_7\
        );

    \I__7385\ : CascadeMux
    port map (
            O => \N__30738\,
            I => \N__30735\
        );

    \I__7384\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30732\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__30732\,
            I => \N__30729\
        );

    \I__7382\ : Span4Mux_v
    port map (
            O => \N__30729\,
            I => \N__30726\
        );

    \I__7381\ : Odrv4
    port map (
            O => \N__30726\,
            I => \M_this_data_tmp_qZ0Z_6\
        );

    \I__7380\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30720\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__30720\,
            I => \N_67_0\
        );

    \I__7378\ : CascadeMux
    port map (
            O => \N__30717\,
            I => \N__30714\
        );

    \I__7377\ : CascadeBuf
    port map (
            O => \N__30714\,
            I => \N__30711\
        );

    \I__7376\ : CascadeMux
    port map (
            O => \N__30711\,
            I => \N__30707\
        );

    \I__7375\ : CascadeMux
    port map (
            O => \N__30710\,
            I => \N__30704\
        );

    \I__7374\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30701\
        );

    \I__7373\ : InMux
    port map (
            O => \N__30704\,
            I => \N__30698\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__30701\,
            I => \N__30695\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__30698\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__7370\ : Odrv12
    port map (
            O => \N__30695\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__7369\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30686\
        );

    \I__7368\ : InMux
    port map (
            O => \N__30689\,
            I => \N__30679\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__30686\,
            I => \N__30676\
        );

    \I__7366\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30671\
        );

    \I__7365\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30671\
        );

    \I__7364\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30668\
        );

    \I__7363\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30665\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__30679\,
            I => \N__30662\
        );

    \I__7361\ : Span4Mux_v
    port map (
            O => \N__30676\,
            I => \N__30655\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__30671\,
            I => \N__30655\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__30668\,
            I => \N__30655\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__30665\,
            I => \N__30652\
        );

    \I__7357\ : Span12Mux_v
    port map (
            O => \N__30662\,
            I => \N__30649\
        );

    \I__7356\ : Span4Mux_h
    port map (
            O => \N__30655\,
            I => \N__30646\
        );

    \I__7355\ : Odrv12
    port map (
            O => \N__30652\,
            I => \N_1152_0\
        );

    \I__7354\ : Odrv12
    port map (
            O => \N__30649\,
            I => \N_1152_0\
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__30646\,
            I => \N_1152_0\
        );

    \I__7352\ : CascadeMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__7351\ : CascadeBuf
    port map (
            O => \N__30636\,
            I => \N__30631\
        );

    \I__7350\ : CascadeMux
    port map (
            O => \N__30635\,
            I => \N__30628\
        );

    \I__7349\ : InMux
    port map (
            O => \N__30634\,
            I => \N__30625\
        );

    \I__7348\ : CascadeMux
    port map (
            O => \N__30631\,
            I => \N__30622\
        );

    \I__7347\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30618\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__30625\,
            I => \N__30615\
        );

    \I__7345\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30612\
        );

    \I__7344\ : InMux
    port map (
            O => \N__30621\,
            I => \N__30609\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__30618\,
            I => \N__30602\
        );

    \I__7342\ : Span12Mux_v
    port map (
            O => \N__30615\,
            I => \N__30602\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__30612\,
            I => \N__30602\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__30609\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__7339\ : Odrv12
    port map (
            O => \N__30602\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__7338\ : CascadeMux
    port map (
            O => \N__30597\,
            I => \N__30594\
        );

    \I__7337\ : CascadeBuf
    port map (
            O => \N__30594\,
            I => \N__30591\
        );

    \I__7336\ : CascadeMux
    port map (
            O => \N__30591\,
            I => \N__30587\
        );

    \I__7335\ : InMux
    port map (
            O => \N__30590\,
            I => \N__30582\
        );

    \I__7334\ : InMux
    port map (
            O => \N__30587\,
            I => \N__30578\
        );

    \I__7333\ : InMux
    port map (
            O => \N__30586\,
            I => \N__30575\
        );

    \I__7332\ : InMux
    port map (
            O => \N__30585\,
            I => \N__30572\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__30582\,
            I => \N__30569\
        );

    \I__7330\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30566\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__30578\,
            I => \N__30563\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__30575\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__30572\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__7326\ : Odrv12
    port map (
            O => \N__30569\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__30566\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__7324\ : Odrv12
    port map (
            O => \N__30563\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__7323\ : InMux
    port map (
            O => \N__30552\,
            I => \N__30547\
        );

    \I__7322\ : InMux
    port map (
            O => \N__30551\,
            I => \N__30542\
        );

    \I__7321\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30542\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__30547\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__30542\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__7318\ : InMux
    port map (
            O => \N__30537\,
            I => \N__30534\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__30534\,
            I => \un1_M_this_oam_address_q_c4\
        );

    \I__7316\ : InMux
    port map (
            O => \N__30531\,
            I => \N__30528\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__30528\,
            I => \N__30525\
        );

    \I__7314\ : Odrv12
    port map (
            O => \N__30525\,
            I => \N_50_0\
        );

    \I__7313\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30519\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__30519\,
            I => \N__30516\
        );

    \I__7311\ : Span4Mux_v
    port map (
            O => \N__30516\,
            I => \N__30513\
        );

    \I__7310\ : Odrv4
    port map (
            O => \N__30513\,
            I => \N_46_0\
        );

    \I__7309\ : CascadeMux
    port map (
            O => \N__30510\,
            I => \N__30507\
        );

    \I__7308\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30504\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__30504\,
            I => \M_this_data_tmp_qZ0Z_21\
        );

    \I__7306\ : CascadeMux
    port map (
            O => \N__30501\,
            I => \N__30498\
        );

    \I__7305\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30495\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__30495\,
            I => \N__30492\
        );

    \I__7303\ : Odrv4
    port map (
            O => \N__30492\,
            I => \M_this_data_tmp_qZ0Z_10\
        );

    \I__7302\ : InMux
    port map (
            O => \N__30489\,
            I => \N__30486\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__30486\,
            I => \N__30483\
        );

    \I__7300\ : Span4Mux_v
    port map (
            O => \N__30483\,
            I => \N__30480\
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__30480\,
            I => \this_sprites_ram.mem_out_bus5_3\
        );

    \I__7298\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30474\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__30474\,
            I => \N__30471\
        );

    \I__7296\ : Span4Mux_v
    port map (
            O => \N__30471\,
            I => \N__30468\
        );

    \I__7295\ : Odrv4
    port map (
            O => \N__30468\,
            I => \this_sprites_ram.mem_out_bus1_3\
        );

    \I__7294\ : InMux
    port map (
            O => \N__30465\,
            I => \N__30461\
        );

    \I__7293\ : InMux
    port map (
            O => \N__30464\,
            I => \N__30450\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__30461\,
            I => \N__30446\
        );

    \I__7291\ : InMux
    port map (
            O => \N__30460\,
            I => \N__30443\
        );

    \I__7290\ : InMux
    port map (
            O => \N__30459\,
            I => \N__30440\
        );

    \I__7289\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30431\
        );

    \I__7288\ : InMux
    port map (
            O => \N__30457\,
            I => \N__30431\
        );

    \I__7287\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30431\
        );

    \I__7286\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30431\
        );

    \I__7285\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30426\
        );

    \I__7284\ : InMux
    port map (
            O => \N__30453\,
            I => \N__30426\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__30450\,
            I => \N__30420\
        );

    \I__7282\ : InMux
    port map (
            O => \N__30449\,
            I => \N__30415\
        );

    \I__7281\ : Span4Mux_h
    port map (
            O => \N__30446\,
            I => \N__30404\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__30443\,
            I => \N__30404\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__30440\,
            I => \N__30404\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__30431\,
            I => \N__30404\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__30426\,
            I => \N__30404\
        );

    \I__7276\ : InMux
    port map (
            O => \N__30425\,
            I => \N__30397\
        );

    \I__7275\ : InMux
    port map (
            O => \N__30424\,
            I => \N__30397\
        );

    \I__7274\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30397\
        );

    \I__7273\ : Span4Mux_h
    port map (
            O => \N__30420\,
            I => \N__30394\
        );

    \I__7272\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30389\
        );

    \I__7271\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30389\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__30415\,
            I => \N__30386\
        );

    \I__7269\ : Span4Mux_h
    port map (
            O => \N__30404\,
            I => \N__30383\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__30397\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7267\ : Odrv4
    port map (
            O => \N__30394\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__30389\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7265\ : Odrv4
    port map (
            O => \N__30386\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7264\ : Odrv4
    port map (
            O => \N__30383\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7263\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30369\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__30369\,
            I => \N__30366\
        );

    \I__7261\ : Span4Mux_h
    port map (
            O => \N__30366\,
            I => \N__30363\
        );

    \I__7260\ : Span4Mux_h
    port map (
            O => \N__30363\,
            I => \N__30360\
        );

    \I__7259\ : Odrv4
    port map (
            O => \N__30360\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\
        );

    \I__7258\ : CEMux
    port map (
            O => \N__30357\,
            I => \N__30353\
        );

    \I__7257\ : CEMux
    port map (
            O => \N__30356\,
            I => \N__30350\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30347\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__30350\,
            I => \N__30344\
        );

    \I__7254\ : Span4Mux_v
    port map (
            O => \N__30347\,
            I => \N__30339\
        );

    \I__7253\ : Span4Mux_h
    port map (
            O => \N__30344\,
            I => \N__30339\
        );

    \I__7252\ : Odrv4
    port map (
            O => \N__30339\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__7251\ : CascadeMux
    port map (
            O => \N__30336\,
            I => \N__30333\
        );

    \I__7250\ : InMux
    port map (
            O => \N__30333\,
            I => \N__30329\
        );

    \I__7249\ : InMux
    port map (
            O => \N__30332\,
            I => \N__30326\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__30329\,
            I => \N__30323\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__30326\,
            I => \this_ppu.M_this_ppu_map_addr_i_5\
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__30323\,
            I => \this_ppu.M_this_ppu_map_addr_i_5\
        );

    \I__7245\ : CascadeMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__7244\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30311\
        );

    \I__7243\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30308\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__30311\,
            I => \N__30305\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__30308\,
            I => \this_ppu.M_this_ppu_map_addr_i_6\
        );

    \I__7240\ : Odrv4
    port map (
            O => \N__30305\,
            I => \this_ppu.M_this_ppu_map_addr_i_6\
        );

    \I__7239\ : CascadeMux
    port map (
            O => \N__30300\,
            I => \N__30297\
        );

    \I__7238\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30293\
        );

    \I__7237\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30290\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__30293\,
            I => \N__30287\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__30290\,
            I => \this_ppu.M_this_ppu_map_addr_i_7\
        );

    \I__7234\ : Odrv4
    port map (
            O => \N__30287\,
            I => \this_ppu.M_this_ppu_map_addr_i_7\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__30282\,
            I => \N__30279\
        );

    \I__7232\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30275\
        );

    \I__7231\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30272\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__30275\,
            I => \N__30269\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__30272\,
            I => \this_ppu.M_this_ppu_map_addr_i_8\
        );

    \I__7228\ : Odrv4
    port map (
            O => \N__30269\,
            I => \this_ppu.M_this_ppu_map_addr_i_8\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__30264\,
            I => \N__30260\
        );

    \I__7226\ : InMux
    port map (
            O => \N__30263\,
            I => \N__30257\
        );

    \I__7225\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30254\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__30257\,
            I => \N__30251\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__30254\,
            I => \this_ppu.M_this_ppu_map_addr_i_9\
        );

    \I__7222\ : Odrv4
    port map (
            O => \N__30251\,
            I => \this_ppu.M_this_ppu_map_addr_i_9\
        );

    \I__7221\ : InMux
    port map (
            O => \N__30246\,
            I => \bfn_23_20_0_\
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__7219\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30237\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__30237\,
            I => \this_ppu.un1_M_vaddress_q_cry_7_THRU_CO\
        );

    \I__7217\ : InMux
    port map (
            O => \N__30234\,
            I => \N__30231\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__30231\,
            I => \N__30228\
        );

    \I__7215\ : Span12Mux_s9_h
    port map (
            O => \N__30228\,
            I => \N__30225\
        );

    \I__7214\ : Odrv12
    port map (
            O => \N__30225\,
            I => \N_61_0\
        );

    \I__7213\ : InMux
    port map (
            O => \N__30222\,
            I => \N__30219\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__30219\,
            I => \N__30216\
        );

    \I__7211\ : Span4Mux_v
    port map (
            O => \N__30216\,
            I => \N__30213\
        );

    \I__7210\ : Odrv4
    port map (
            O => \N__30213\,
            I => \M_this_data_tmp_qZ0Z_3\
        );

    \I__7209\ : InMux
    port map (
            O => \N__30210\,
            I => \N__30207\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__30207\,
            I => \N__30204\
        );

    \I__7207\ : Span4Mux_v
    port map (
            O => \N__30204\,
            I => \N__30201\
        );

    \I__7206\ : Odrv4
    port map (
            O => \N__30201\,
            I => \N_73_0\
        );

    \I__7205\ : CascadeMux
    port map (
            O => \N__30198\,
            I => \N__30195\
        );

    \I__7204\ : CascadeBuf
    port map (
            O => \N__30195\,
            I => \N__30192\
        );

    \I__7203\ : CascadeMux
    port map (
            O => \N__30192\,
            I => \N__30188\
        );

    \I__7202\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30185\
        );

    \I__7201\ : InMux
    port map (
            O => \N__30188\,
            I => \N__30182\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__30185\,
            I => \N__30176\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__30182\,
            I => \N__30176\
        );

    \I__7198\ : InMux
    port map (
            O => \N__30181\,
            I => \N__30173\
        );

    \I__7197\ : Span4Mux_h
    port map (
            O => \N__30176\,
            I => \N__30170\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__30173\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__7195\ : Odrv4
    port map (
            O => \N__30170\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__7194\ : CascadeMux
    port map (
            O => \N__30165\,
            I => \N__30157\
        );

    \I__7193\ : CascadeMux
    port map (
            O => \N__30164\,
            I => \N__30154\
        );

    \I__7192\ : CascadeMux
    port map (
            O => \N__30163\,
            I => \N__30149\
        );

    \I__7191\ : CascadeMux
    port map (
            O => \N__30162\,
            I => \N__30146\
        );

    \I__7190\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30142\
        );

    \I__7189\ : InMux
    port map (
            O => \N__30160\,
            I => \N__30137\
        );

    \I__7188\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30137\
        );

    \I__7187\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30133\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__30153\,
            I => \N__30130\
        );

    \I__7185\ : InMux
    port map (
            O => \N__30152\,
            I => \N__30127\
        );

    \I__7184\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30124\
        );

    \I__7183\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30121\
        );

    \I__7182\ : CascadeMux
    port map (
            O => \N__30145\,
            I => \N__30118\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__30142\,
            I => \N__30113\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__30137\,
            I => \N__30113\
        );

    \I__7179\ : CascadeMux
    port map (
            O => \N__30136\,
            I => \N__30109\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__30133\,
            I => \N__30105\
        );

    \I__7177\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30102\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__30127\,
            I => \N__30097\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__30124\,
            I => \N__30097\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__30121\,
            I => \N__30094\
        );

    \I__7173\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30091\
        );

    \I__7172\ : Span4Mux_v
    port map (
            O => \N__30113\,
            I => \N__30088\
        );

    \I__7171\ : InMux
    port map (
            O => \N__30112\,
            I => \N__30083\
        );

    \I__7170\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30083\
        );

    \I__7169\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30078\
        );

    \I__7168\ : Span4Mux_h
    port map (
            O => \N__30105\,
            I => \N__30075\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__30102\,
            I => \N__30072\
        );

    \I__7166\ : Span4Mux_v
    port map (
            O => \N__30097\,
            I => \N__30069\
        );

    \I__7165\ : Span4Mux_h
    port map (
            O => \N__30094\,
            I => \N__30064\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__30091\,
            I => \N__30064\
        );

    \I__7163\ : Span4Mux_h
    port map (
            O => \N__30088\,
            I => \N__30059\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__30083\,
            I => \N__30059\
        );

    \I__7161\ : CascadeMux
    port map (
            O => \N__30082\,
            I => \N__30056\
        );

    \I__7160\ : InMux
    port map (
            O => \N__30081\,
            I => \N__30052\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__30078\,
            I => \N__30045\
        );

    \I__7158\ : Span4Mux_h
    port map (
            O => \N__30075\,
            I => \N__30045\
        );

    \I__7157\ : Span4Mux_h
    port map (
            O => \N__30072\,
            I => \N__30045\
        );

    \I__7156\ : Span4Mux_h
    port map (
            O => \N__30069\,
            I => \N__30038\
        );

    \I__7155\ : Span4Mux_h
    port map (
            O => \N__30064\,
            I => \N__30038\
        );

    \I__7154\ : Span4Mux_h
    port map (
            O => \N__30059\,
            I => \N__30038\
        );

    \I__7153\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30033\
        );

    \I__7152\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30033\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__30052\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__7150\ : Odrv4
    port map (
            O => \N__30045\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__7149\ : Odrv4
    port map (
            O => \N__30038\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__30033\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__7147\ : CascadeMux
    port map (
            O => \N__30024\,
            I => \this_ppu.un2_vscroll_axb_0_cascade_\
        );

    \I__7146\ : InMux
    port map (
            O => \N__30021\,
            I => \N__30013\
        );

    \I__7145\ : InMux
    port map (
            O => \N__30020\,
            I => \N__30010\
        );

    \I__7144\ : InMux
    port map (
            O => \N__30019\,
            I => \N__30007\
        );

    \I__7143\ : CascadeMux
    port map (
            O => \N__30018\,
            I => \N__30003\
        );

    \I__7142\ : InMux
    port map (
            O => \N__30017\,
            I => \N__29992\
        );

    \I__7141\ : InMux
    port map (
            O => \N__30016\,
            I => \N__29992\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__30013\,
            I => \N__29987\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__30010\,
            I => \N__29982\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__30007\,
            I => \N__29982\
        );

    \I__7137\ : InMux
    port map (
            O => \N__30006\,
            I => \N__29979\
        );

    \I__7136\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29975\
        );

    \I__7135\ : InMux
    port map (
            O => \N__30002\,
            I => \N__29972\
        );

    \I__7134\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29969\
        );

    \I__7133\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29966\
        );

    \I__7132\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29963\
        );

    \I__7131\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29958\
        );

    \I__7130\ : InMux
    port map (
            O => \N__29997\,
            I => \N__29958\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__29992\,
            I => \N__29955\
        );

    \I__7128\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29952\
        );

    \I__7127\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29949\
        );

    \I__7126\ : Span4Mux_v
    port map (
            O => \N__29987\,
            I => \N__29942\
        );

    \I__7125\ : Span4Mux_h
    port map (
            O => \N__29982\,
            I => \N__29942\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__29979\,
            I => \N__29942\
        );

    \I__7123\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29938\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__29975\,
            I => \N__29931\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__29972\,
            I => \N__29931\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__29969\,
            I => \N__29931\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__29966\,
            I => \N__29928\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__29963\,
            I => \N__29919\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__29958\,
            I => \N__29919\
        );

    \I__7116\ : Span4Mux_v
    port map (
            O => \N__29955\,
            I => \N__29919\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__29952\,
            I => \N__29919\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__29949\,
            I => \N__29916\
        );

    \I__7113\ : Span4Mux_h
    port map (
            O => \N__29942\,
            I => \N__29913\
        );

    \I__7112\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29910\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__29938\,
            I => \N__29907\
        );

    \I__7110\ : Span12Mux_h
    port map (
            O => \N__29931\,
            I => \N__29904\
        );

    \I__7109\ : Span4Mux_v
    port map (
            O => \N__29928\,
            I => \N__29899\
        );

    \I__7108\ : Span4Mux_h
    port map (
            O => \N__29919\,
            I => \N__29899\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__29916\,
            I => \N__29896\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__29913\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__29910\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__29907\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7103\ : Odrv12
    port map (
            O => \N__29904\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7102\ : Odrv4
    port map (
            O => \N__29899\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7101\ : Odrv4
    port map (
            O => \N__29896\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7100\ : CascadeMux
    port map (
            O => \N__29883\,
            I => \N__29879\
        );

    \I__7099\ : CascadeMux
    port map (
            O => \N__29882\,
            I => \N__29876\
        );

    \I__7098\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29871\
        );

    \I__7097\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29866\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__29875\,
            I => \N__29863\
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__29874\,
            I => \N__29859\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__29871\,
            I => \N__29855\
        );

    \I__7093\ : CascadeMux
    port map (
            O => \N__29870\,
            I => \N__29852\
        );

    \I__7092\ : CascadeMux
    port map (
            O => \N__29869\,
            I => \N__29848\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29844\
        );

    \I__7090\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29841\
        );

    \I__7089\ : CascadeMux
    port map (
            O => \N__29862\,
            I => \N__29838\
        );

    \I__7088\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29835\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__29858\,
            I => \N__29832\
        );

    \I__7086\ : Span4Mux_h
    port map (
            O => \N__29855\,
            I => \N__29829\
        );

    \I__7085\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29826\
        );

    \I__7084\ : CascadeMux
    port map (
            O => \N__29851\,
            I => \N__29823\
        );

    \I__7083\ : InMux
    port map (
            O => \N__29848\,
            I => \N__29819\
        );

    \I__7082\ : CascadeMux
    port map (
            O => \N__29847\,
            I => \N__29816\
        );

    \I__7081\ : Span4Mux_v
    port map (
            O => \N__29844\,
            I => \N__29809\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__29841\,
            I => \N__29809\
        );

    \I__7079\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29805\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__29835\,
            I => \N__29802\
        );

    \I__7077\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29799\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__29829\,
            I => \N__29793\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__29826\,
            I => \N__29793\
        );

    \I__7074\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29790\
        );

    \I__7073\ : CascadeMux
    port map (
            O => \N__29822\,
            I => \N__29787\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__29819\,
            I => \N__29784\
        );

    \I__7071\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29781\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__29815\,
            I => \N__29778\
        );

    \I__7069\ : CascadeMux
    port map (
            O => \N__29814\,
            I => \N__29774\
        );

    \I__7068\ : Span4Mux_h
    port map (
            O => \N__29809\,
            I => \N__29771\
        );

    \I__7067\ : CascadeMux
    port map (
            O => \N__29808\,
            I => \N__29768\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__29805\,
            I => \N__29765\
        );

    \I__7065\ : Span4Mux_h
    port map (
            O => \N__29802\,
            I => \N__29762\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__29799\,
            I => \N__29759\
        );

    \I__7063\ : CascadeMux
    port map (
            O => \N__29798\,
            I => \N__29756\
        );

    \I__7062\ : Span4Mux_h
    port map (
            O => \N__29793\,
            I => \N__29753\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__29790\,
            I => \N__29750\
        );

    \I__7060\ : InMux
    port map (
            O => \N__29787\,
            I => \N__29747\
        );

    \I__7059\ : Span4Mux_h
    port map (
            O => \N__29784\,
            I => \N__29744\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__29781\,
            I => \N__29741\
        );

    \I__7057\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29738\
        );

    \I__7056\ : CascadeMux
    port map (
            O => \N__29777\,
            I => \N__29735\
        );

    \I__7055\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29732\
        );

    \I__7054\ : Sp12to4
    port map (
            O => \N__29771\,
            I => \N__29729\
        );

    \I__7053\ : InMux
    port map (
            O => \N__29768\,
            I => \N__29726\
        );

    \I__7052\ : Span4Mux_h
    port map (
            O => \N__29765\,
            I => \N__29723\
        );

    \I__7051\ : Span4Mux_v
    port map (
            O => \N__29762\,
            I => \N__29718\
        );

    \I__7050\ : Span4Mux_h
    port map (
            O => \N__29759\,
            I => \N__29718\
        );

    \I__7049\ : InMux
    port map (
            O => \N__29756\,
            I => \N__29715\
        );

    \I__7048\ : Span4Mux_h
    port map (
            O => \N__29753\,
            I => \N__29712\
        );

    \I__7047\ : Span4Mux_h
    port map (
            O => \N__29750\,
            I => \N__29709\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__29747\,
            I => \N__29706\
        );

    \I__7045\ : Span4Mux_v
    port map (
            O => \N__29744\,
            I => \N__29701\
        );

    \I__7044\ : Span4Mux_h
    port map (
            O => \N__29741\,
            I => \N__29701\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__29738\,
            I => \N__29698\
        );

    \I__7042\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29695\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__29732\,
            I => \N__29692\
        );

    \I__7040\ : Span12Mux_h
    port map (
            O => \N__29729\,
            I => \N__29687\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__29726\,
            I => \N__29687\
        );

    \I__7038\ : Span4Mux_v
    port map (
            O => \N__29723\,
            I => \N__29684\
        );

    \I__7037\ : Span4Mux_v
    port map (
            O => \N__29718\,
            I => \N__29681\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29678\
        );

    \I__7035\ : Span4Mux_h
    port map (
            O => \N__29712\,
            I => \N__29675\
        );

    \I__7034\ : Span4Mux_v
    port map (
            O => \N__29709\,
            I => \N__29670\
        );

    \I__7033\ : Span4Mux_h
    port map (
            O => \N__29706\,
            I => \N__29670\
        );

    \I__7032\ : Span4Mux_v
    port map (
            O => \N__29701\,
            I => \N__29665\
        );

    \I__7031\ : Span4Mux_h
    port map (
            O => \N__29698\,
            I => \N__29665\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__29695\,
            I => \N__29662\
        );

    \I__7029\ : Span12Mux_s9_h
    port map (
            O => \N__29692\,
            I => \N__29657\
        );

    \I__7028\ : Span12Mux_s9_h
    port map (
            O => \N__29687\,
            I => \N__29657\
        );

    \I__7027\ : Span4Mux_v
    port map (
            O => \N__29684\,
            I => \N__29650\
        );

    \I__7026\ : Span4Mux_v
    port map (
            O => \N__29681\,
            I => \N__29650\
        );

    \I__7025\ : Span4Mux_h
    port map (
            O => \N__29678\,
            I => \N__29650\
        );

    \I__7024\ : Span4Mux_h
    port map (
            O => \N__29675\,
            I => \N__29641\
        );

    \I__7023\ : Span4Mux_v
    port map (
            O => \N__29670\,
            I => \N__29641\
        );

    \I__7022\ : Span4Mux_v
    port map (
            O => \N__29665\,
            I => \N__29641\
        );

    \I__7021\ : Span4Mux_h
    port map (
            O => \N__29662\,
            I => \N__29641\
        );

    \I__7020\ : Odrv12
    port map (
            O => \N__29657\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__29650\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__7018\ : Odrv4
    port map (
            O => \N__29641\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__7017\ : InMux
    port map (
            O => \N__29634\,
            I => \N__29619\
        );

    \I__7016\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29619\
        );

    \I__7015\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29619\
        );

    \I__7014\ : InMux
    port map (
            O => \N__29631\,
            I => \N__29619\
        );

    \I__7013\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29616\
        );

    \I__7012\ : InMux
    port map (
            O => \N__29629\,
            I => \N__29613\
        );

    \I__7011\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29610\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__29619\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__29616\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__29613\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__29610\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7006\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29595\
        );

    \I__7005\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29595\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__29595\,
            I => \N__29591\
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__29594\,
            I => \N__29588\
        );

    \I__7002\ : Span4Mux_h
    port map (
            O => \N__29591\,
            I => \N__29585\
        );

    \I__7001\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29582\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__29585\,
            I => \this_ppu.un1_M_vaddress_q_2_c2\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__29582\,
            I => \this_ppu.un1_M_vaddress_q_2_c2\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__29577\,
            I => \N__29574\
        );

    \I__6997\ : CascadeBuf
    port map (
            O => \N__29574\,
            I => \N__29571\
        );

    \I__6996\ : CascadeMux
    port map (
            O => \N__29571\,
            I => \N__29568\
        );

    \I__6995\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__29565\,
            I => \N__29561\
        );

    \I__6993\ : CascadeMux
    port map (
            O => \N__29564\,
            I => \N__29558\
        );

    \I__6992\ : Span12Mux_s10_h
    port map (
            O => \N__29561\,
            I => \N__29552\
        );

    \I__6991\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29547\
        );

    \I__6990\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29547\
        );

    \I__6989\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29544\
        );

    \I__6988\ : InMux
    port map (
            O => \N__29555\,
            I => \N__29541\
        );

    \I__6987\ : Span12Mux_h
    port map (
            O => \N__29552\,
            I => \N__29538\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__29547\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__29544\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__29541\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__6983\ : Odrv12
    port map (
            O => \N__29538\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__6982\ : CascadeMux
    port map (
            O => \N__29529\,
            I => \N__29526\
        );

    \I__6981\ : CascadeBuf
    port map (
            O => \N__29526\,
            I => \N__29523\
        );

    \I__6980\ : CascadeMux
    port map (
            O => \N__29523\,
            I => \N__29520\
        );

    \I__6979\ : InMux
    port map (
            O => \N__29520\,
            I => \N__29517\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__29517\,
            I => \N__29514\
        );

    \I__6977\ : Span4Mux_h
    port map (
            O => \N__29514\,
            I => \N__29511\
        );

    \I__6976\ : Sp12to4
    port map (
            O => \N__29511\,
            I => \N__29508\
        );

    \I__6975\ : Span12Mux_s10_v
    port map (
            O => \N__29508\,
            I => \N__29502\
        );

    \I__6974\ : InMux
    port map (
            O => \N__29507\,
            I => \N__29499\
        );

    \I__6973\ : InMux
    port map (
            O => \N__29506\,
            I => \N__29496\
        );

    \I__6972\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29493\
        );

    \I__6971\ : Span12Mux_h
    port map (
            O => \N__29502\,
            I => \N__29490\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__29499\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__29496\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__29493\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__6967\ : Odrv12
    port map (
            O => \N__29490\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__6966\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__29478\,
            I => \N__29475\
        );

    \I__6964\ : Span4Mux_v
    port map (
            O => \N__29475\,
            I => \N__29468\
        );

    \I__6963\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29465\
        );

    \I__6962\ : InMux
    port map (
            O => \N__29473\,
            I => \N__29460\
        );

    \I__6961\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29460\
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__29471\,
            I => \N__29457\
        );

    \I__6959\ : Span4Mux_h
    port map (
            O => \N__29468\,
            I => \N__29451\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__29465\,
            I => \N__29451\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__29460\,
            I => \N__29448\
        );

    \I__6956\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29443\
        );

    \I__6955\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29443\
        );

    \I__6954\ : Odrv4
    port map (
            O => \N__29451\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__6953\ : Odrv4
    port map (
            O => \N__29448\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__29443\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__29436\,
            I => \N__29431\
        );

    \I__6950\ : CascadeMux
    port map (
            O => \N__29435\,
            I => \N__29428\
        );

    \I__6949\ : CascadeMux
    port map (
            O => \N__29434\,
            I => \N__29424\
        );

    \I__6948\ : InMux
    port map (
            O => \N__29431\,
            I => \N__29421\
        );

    \I__6947\ : InMux
    port map (
            O => \N__29428\,
            I => \N__29418\
        );

    \I__6946\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29413\
        );

    \I__6945\ : InMux
    port map (
            O => \N__29424\,
            I => \N__29413\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__29421\,
            I => \N__29410\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__29418\,
            I => \N__29407\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__29413\,
            I => \N__29404\
        );

    \I__6941\ : Sp12to4
    port map (
            O => \N__29410\,
            I => \N__29399\
        );

    \I__6940\ : Span4Mux_h
    port map (
            O => \N__29407\,
            I => \N__29396\
        );

    \I__6939\ : Span4Mux_v
    port map (
            O => \N__29404\,
            I => \N__29393\
        );

    \I__6938\ : InMux
    port map (
            O => \N__29403\,
            I => \N__29388\
        );

    \I__6937\ : InMux
    port map (
            O => \N__29402\,
            I => \N__29388\
        );

    \I__6936\ : Odrv12
    port map (
            O => \N__29399\,
            I => \this_ppu.M_last_q\
        );

    \I__6935\ : Odrv4
    port map (
            O => \N__29396\,
            I => \this_ppu.M_last_q\
        );

    \I__6934\ : Odrv4
    port map (
            O => \N__29393\,
            I => \this_ppu.M_last_q\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__29388\,
            I => \this_ppu.M_last_q\
        );

    \I__6932\ : InMux
    port map (
            O => \N__29379\,
            I => \N__29376\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__29376\,
            I => \N__29373\
        );

    \I__6930\ : Span4Mux_v
    port map (
            O => \N__29373\,
            I => \N__29367\
        );

    \I__6929\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29364\
        );

    \I__6928\ : InMux
    port map (
            O => \N__29371\,
            I => \N__29359\
        );

    \I__6927\ : InMux
    port map (
            O => \N__29370\,
            I => \N__29359\
        );

    \I__6926\ : Span4Mux_h
    port map (
            O => \N__29367\,
            I => \N__29352\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__29364\,
            I => \N__29352\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__29359\,
            I => \N__29349\
        );

    \I__6923\ : InMux
    port map (
            O => \N__29358\,
            I => \N__29344\
        );

    \I__6922\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29344\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__29352\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__29349\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__29344\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__6918\ : CascadeMux
    port map (
            O => \N__29337\,
            I => \N__29334\
        );

    \I__6917\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29331\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__29328\,
            I => \N__29323\
        );

    \I__6914\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29320\
        );

    \I__6913\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29316\
        );

    \I__6912\ : Sp12to4
    port map (
            O => \N__29323\,
            I => \N__29313\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__29320\,
            I => \N__29310\
        );

    \I__6910\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29307\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__29316\,
            I => \N__29299\
        );

    \I__6908\ : Span12Mux_h
    port map (
            O => \N__29313\,
            I => \N__29296\
        );

    \I__6907\ : Span4Mux_h
    port map (
            O => \N__29310\,
            I => \N__29291\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__29307\,
            I => \N__29291\
        );

    \I__6905\ : InMux
    port map (
            O => \N__29306\,
            I => \N__29284\
        );

    \I__6904\ : InMux
    port map (
            O => \N__29305\,
            I => \N__29284\
        );

    \I__6903\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29284\
        );

    \I__6902\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29281\
        );

    \I__6901\ : InMux
    port map (
            O => \N__29302\,
            I => \N__29278\
        );

    \I__6900\ : Odrv4
    port map (
            O => \N__29299\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6899\ : Odrv12
    port map (
            O => \N__29296\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__29291\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__29284\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__29281\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__29278\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6894\ : SRMux
    port map (
            O => \N__29265\,
            I => \N__29261\
        );

    \I__6893\ : SRMux
    port map (
            O => \N__29264\,
            I => \N__29258\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__29261\,
            I => \N__29255\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__29258\,
            I => \N__29252\
        );

    \I__6890\ : Span4Mux_h
    port map (
            O => \N__29255\,
            I => \N__29249\
        );

    \I__6889\ : Span4Mux_h
    port map (
            O => \N__29252\,
            I => \N__29246\
        );

    \I__6888\ : Odrv4
    port map (
            O => \N__29249\,
            I => \this_ppu.M_state_q_RNI42KTAZ0Z_0\
        );

    \I__6887\ : Odrv4
    port map (
            O => \N__29246\,
            I => \this_ppu.M_state_q_RNI42KTAZ0Z_0\
        );

    \I__6886\ : CascadeMux
    port map (
            O => \N__29241\,
            I => \N__29238\
        );

    \I__6885\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29235\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__6883\ : Span4Mux_h
    port map (
            O => \N__29232\,
            I => \N__29229\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__29229\,
            I => \M_this_data_tmp_qZ0Z_4\
        );

    \I__6881\ : InMux
    port map (
            O => \N__29226\,
            I => \N__29223\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__29223\,
            I => \N__29220\
        );

    \I__6879\ : Span4Mux_h
    port map (
            O => \N__29220\,
            I => \N__29217\
        );

    \I__6878\ : Odrv4
    port map (
            O => \N__29217\,
            I => \N_71_0\
        );

    \I__6877\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29210\
        );

    \I__6876\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29207\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__29210\,
            I => \N__29204\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__29207\,
            I => \this_ppu.M_this_ppu_vram_addr_i_7\
        );

    \I__6873\ : Odrv4
    port map (
            O => \N__29204\,
            I => \this_ppu.M_this_ppu_vram_addr_i_7\
        );

    \I__6872\ : InMux
    port map (
            O => \N__29199\,
            I => \N__29194\
        );

    \I__6871\ : CascadeMux
    port map (
            O => \N__29198\,
            I => \N__29190\
        );

    \I__6870\ : CascadeMux
    port map (
            O => \N__29197\,
            I => \N__29187\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__29194\,
            I => \N__29184\
        );

    \I__6868\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29181\
        );

    \I__6867\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29178\
        );

    \I__6866\ : InMux
    port map (
            O => \N__29187\,
            I => \N__29175\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__29184\,
            I => \N__29172\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__29181\,
            I => \N__29167\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__29178\,
            I => \N__29167\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__29175\,
            I => \N__29164\
        );

    \I__6861\ : Span4Mux_v
    port map (
            O => \N__29172\,
            I => \N__29161\
        );

    \I__6860\ : Span4Mux_h
    port map (
            O => \N__29167\,
            I => \N__29158\
        );

    \I__6859\ : Span4Mux_h
    port map (
            O => \N__29164\,
            I => \N__29155\
        );

    \I__6858\ : Odrv4
    port map (
            O => \N__29161\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__6857\ : Odrv4
    port map (
            O => \N__29158\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__6856\ : Odrv4
    port map (
            O => \N__29155\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__6855\ : InMux
    port map (
            O => \N__29148\,
            I => \N__29144\
        );

    \I__6854\ : InMux
    port map (
            O => \N__29147\,
            I => \N__29141\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__29144\,
            I => \N__29138\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__29141\,
            I => \this_ppu.M_vaddress_q_i_1\
        );

    \I__6851\ : Odrv4
    port map (
            O => \N__29138\,
            I => \this_ppu.M_vaddress_q_i_1\
        );

    \I__6850\ : InMux
    port map (
            O => \N__29133\,
            I => \N__29129\
        );

    \I__6849\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29126\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__29129\,
            I => \N__29123\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__29126\,
            I => \this_ppu.M_vaddress_q_i_2\
        );

    \I__6846\ : Odrv4
    port map (
            O => \N__29123\,
            I => \this_ppu.M_vaddress_q_i_2\
        );

    \I__6845\ : CascadeMux
    port map (
            O => \N__29118\,
            I => \N__29113\
        );

    \I__6844\ : CascadeMux
    port map (
            O => \N__29117\,
            I => \N__29110\
        );

    \I__6843\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29107\
        );

    \I__6842\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29104\
        );

    \I__6841\ : InMux
    port map (
            O => \N__29110\,
            I => \N__29101\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__29107\,
            I => \N__29098\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__29104\,
            I => \N__29095\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__29101\,
            I => \N__29092\
        );

    \I__6837\ : Span4Mux_h
    port map (
            O => \N__29098\,
            I => \N__29089\
        );

    \I__6836\ : Span4Mux_v
    port map (
            O => \N__29095\,
            I => \N__29086\
        );

    \I__6835\ : Span4Mux_h
    port map (
            O => \N__29092\,
            I => \N__29083\
        );

    \I__6834\ : Odrv4
    port map (
            O => \N__29089\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__29086\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__29083\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__6831\ : CascadeMux
    port map (
            O => \N__29076\,
            I => \N__29073\
        );

    \I__6830\ : InMux
    port map (
            O => \N__29073\,
            I => \N__29070\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__29070\,
            I => \N__29067\
        );

    \I__6828\ : Odrv4
    port map (
            O => \N__29067\,
            I => \M_this_data_tmp_qZ0Z_15\
        );

    \I__6827\ : InMux
    port map (
            O => \N__29064\,
            I => \N__29061\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__29061\,
            I => \N__29058\
        );

    \I__6825\ : Span4Mux_v
    port map (
            O => \N__29058\,
            I => \N__29055\
        );

    \I__6824\ : Sp12to4
    port map (
            O => \N__29055\,
            I => \N__29052\
        );

    \I__6823\ : Odrv12
    port map (
            O => \N__29052\,
            I => \M_this_oam_ram_write_data_15\
        );

    \I__6822\ : CascadeMux
    port map (
            O => \N__29049\,
            I => \N__29046\
        );

    \I__6821\ : InMux
    port map (
            O => \N__29046\,
            I => \N__29043\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__29043\,
            I => \this_ppu.M_this_oam_ram_read_data_i_16\
        );

    \I__6819\ : InMux
    port map (
            O => \N__29040\,
            I => \N__29037\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__29037\,
            I => \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0\
        );

    \I__6817\ : InMux
    port map (
            O => \N__29034\,
            I => \this_ppu.un2_vscroll_cry_0\
        );

    \I__6816\ : InMux
    port map (
            O => \N__29031\,
            I => \this_ppu.un2_vscroll_cry_1\
        );

    \I__6815\ : CascadeMux
    port map (
            O => \N__29028\,
            I => \N__29025\
        );

    \I__6814\ : InMux
    port map (
            O => \N__29025\,
            I => \N__29022\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__29022\,
            I => \N__29019\
        );

    \I__6812\ : Span4Mux_v
    port map (
            O => \N__29019\,
            I => \N__29016\
        );

    \I__6811\ : Sp12to4
    port map (
            O => \N__29016\,
            I => \N__29013\
        );

    \I__6810\ : Span12Mux_h
    port map (
            O => \N__29013\,
            I => \N__29010\
        );

    \I__6809\ : Span12Mux_v
    port map (
            O => \N__29010\,
            I => \N__29007\
        );

    \I__6808\ : Odrv12
    port map (
            O => \N__29007\,
            I => \M_this_map_ram_read_data_6\
        );

    \I__6807\ : CascadeMux
    port map (
            O => \N__29004\,
            I => \N__29000\
        );

    \I__6806\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28996\
        );

    \I__6805\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28993\
        );

    \I__6804\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28990\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__28996\,
            I => \N__28986\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__28993\,
            I => \N__28983\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__28990\,
            I => \N__28980\
        );

    \I__6800\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28977\
        );

    \I__6799\ : Span4Mux_h
    port map (
            O => \N__28986\,
            I => \N__28974\
        );

    \I__6798\ : Span4Mux_v
    port map (
            O => \N__28983\,
            I => \N__28967\
        );

    \I__6797\ : Span4Mux_h
    port map (
            O => \N__28980\,
            I => \N__28967\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__28977\,
            I => \N__28967\
        );

    \I__6795\ : Span4Mux_h
    port map (
            O => \N__28974\,
            I => \N__28964\
        );

    \I__6794\ : Span4Mux_h
    port map (
            O => \N__28967\,
            I => \N__28961\
        );

    \I__6793\ : Odrv4
    port map (
            O => \N__28964\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__6792\ : Odrv4
    port map (
            O => \N__28961\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__6791\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28953\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__28953\,
            I => \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0\
        );

    \I__6789\ : CascadeMux
    port map (
            O => \N__28950\,
            I => \N__28945\
        );

    \I__6788\ : CascadeMux
    port map (
            O => \N__28949\,
            I => \N__28941\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__28948\,
            I => \N__28938\
        );

    \I__6786\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28934\
        );

    \I__6785\ : CascadeMux
    port map (
            O => \N__28944\,
            I => \N__28931\
        );

    \I__6784\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28927\
        );

    \I__6783\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28924\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__28937\,
            I => \N__28921\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__28934\,
            I => \N__28915\
        );

    \I__6780\ : InMux
    port map (
            O => \N__28931\,
            I => \N__28912\
        );

    \I__6779\ : CascadeMux
    port map (
            O => \N__28930\,
            I => \N__28909\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__28927\,
            I => \N__28906\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__28924\,
            I => \N__28903\
        );

    \I__6776\ : InMux
    port map (
            O => \N__28921\,
            I => \N__28900\
        );

    \I__6775\ : CascadeMux
    port map (
            O => \N__28920\,
            I => \N__28897\
        );

    \I__6774\ : CascadeMux
    port map (
            O => \N__28919\,
            I => \N__28893\
        );

    \I__6773\ : CascadeMux
    port map (
            O => \N__28918\,
            I => \N__28890\
        );

    \I__6772\ : Span4Mux_h
    port map (
            O => \N__28915\,
            I => \N__28885\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__28912\,
            I => \N__28882\
        );

    \I__6770\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28879\
        );

    \I__6769\ : Span4Mux_h
    port map (
            O => \N__28906\,
            I => \N__28875\
        );

    \I__6768\ : Span4Mux_v
    port map (
            O => \N__28903\,
            I => \N__28870\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__28900\,
            I => \N__28870\
        );

    \I__6766\ : InMux
    port map (
            O => \N__28897\,
            I => \N__28867\
        );

    \I__6765\ : CascadeMux
    port map (
            O => \N__28896\,
            I => \N__28864\
        );

    \I__6764\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28861\
        );

    \I__6763\ : InMux
    port map (
            O => \N__28890\,
            I => \N__28858\
        );

    \I__6762\ : CascadeMux
    port map (
            O => \N__28889\,
            I => \N__28855\
        );

    \I__6761\ : CascadeMux
    port map (
            O => \N__28888\,
            I => \N__28852\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__28885\,
            I => \N__28845\
        );

    \I__6759\ : Span4Mux_h
    port map (
            O => \N__28882\,
            I => \N__28845\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__28879\,
            I => \N__28842\
        );

    \I__6757\ : CascadeMux
    port map (
            O => \N__28878\,
            I => \N__28838\
        );

    \I__6756\ : Span4Mux_h
    port map (
            O => \N__28875\,
            I => \N__28835\
        );

    \I__6755\ : Span4Mux_v
    port map (
            O => \N__28870\,
            I => \N__28830\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28830\
        );

    \I__6753\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28827\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__28861\,
            I => \N__28822\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28822\
        );

    \I__6750\ : InMux
    port map (
            O => \N__28855\,
            I => \N__28819\
        );

    \I__6749\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28816\
        );

    \I__6748\ : CascadeMux
    port map (
            O => \N__28851\,
            I => \N__28813\
        );

    \I__6747\ : CascadeMux
    port map (
            O => \N__28850\,
            I => \N__28810\
        );

    \I__6746\ : Span4Mux_v
    port map (
            O => \N__28845\,
            I => \N__28805\
        );

    \I__6745\ : Span4Mux_h
    port map (
            O => \N__28842\,
            I => \N__28805\
        );

    \I__6744\ : CascadeMux
    port map (
            O => \N__28841\,
            I => \N__28802\
        );

    \I__6743\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28799\
        );

    \I__6742\ : Span4Mux_h
    port map (
            O => \N__28835\,
            I => \N__28796\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__28830\,
            I => \N__28791\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__28827\,
            I => \N__28791\
        );

    \I__6739\ : Span4Mux_v
    port map (
            O => \N__28822\,
            I => \N__28784\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__28819\,
            I => \N__28784\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__28816\,
            I => \N__28784\
        );

    \I__6736\ : InMux
    port map (
            O => \N__28813\,
            I => \N__28781\
        );

    \I__6735\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28778\
        );

    \I__6734\ : Span4Mux_h
    port map (
            O => \N__28805\,
            I => \N__28775\
        );

    \I__6733\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28772\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__28799\,
            I => \N__28769\
        );

    \I__6731\ : Span4Mux_h
    port map (
            O => \N__28796\,
            I => \N__28766\
        );

    \I__6730\ : Span4Mux_v
    port map (
            O => \N__28791\,
            I => \N__28763\
        );

    \I__6729\ : Span4Mux_v
    port map (
            O => \N__28784\,
            I => \N__28758\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__28781\,
            I => \N__28758\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__28778\,
            I => \N__28755\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__28775\,
            I => \N__28752\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__28772\,
            I => \N__28749\
        );

    \I__6724\ : Span12Mux_s9_h
    port map (
            O => \N__28769\,
            I => \N__28746\
        );

    \I__6723\ : Span4Mux_v
    port map (
            O => \N__28766\,
            I => \N__28739\
        );

    \I__6722\ : Span4Mux_v
    port map (
            O => \N__28763\,
            I => \N__28739\
        );

    \I__6721\ : Span4Mux_v
    port map (
            O => \N__28758\,
            I => \N__28739\
        );

    \I__6720\ : Span4Mux_h
    port map (
            O => \N__28755\,
            I => \N__28736\
        );

    \I__6719\ : Span4Mux_h
    port map (
            O => \N__28752\,
            I => \N__28731\
        );

    \I__6718\ : Span4Mux_h
    port map (
            O => \N__28749\,
            I => \N__28731\
        );

    \I__6717\ : Odrv12
    port map (
            O => \N__28746\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__6716\ : Odrv4
    port map (
            O => \N__28739\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__28736\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__28731\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__28722\,
            I => \N__28717\
        );

    \I__6712\ : CascadeMux
    port map (
            O => \N__28721\,
            I => \N__28712\
        );

    \I__6711\ : InMux
    port map (
            O => \N__28720\,
            I => \N__28708\
        );

    \I__6710\ : InMux
    port map (
            O => \N__28717\,
            I => \N__28705\
        );

    \I__6709\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28702\
        );

    \I__6708\ : InMux
    port map (
            O => \N__28715\,
            I => \N__28699\
        );

    \I__6707\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28694\
        );

    \I__6706\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28694\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__28708\,
            I => \N__28689\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28689\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__28702\,
            I => \N__28686\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__28699\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__28694\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6700\ : Odrv4
    port map (
            O => \N__28689\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6699\ : Odrv4
    port map (
            O => \N__28686\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6698\ : CascadeMux
    port map (
            O => \N__28677\,
            I => \N__28673\
        );

    \I__6697\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28669\
        );

    \I__6696\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28665\
        );

    \I__6695\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28660\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__28669\,
            I => \N__28657\
        );

    \I__6693\ : CascadeMux
    port map (
            O => \N__28668\,
            I => \N__28654\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__28665\,
            I => \N__28651\
        );

    \I__6691\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28646\
        );

    \I__6690\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28646\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__28660\,
            I => \N__28643\
        );

    \I__6688\ : Span4Mux_h
    port map (
            O => \N__28657\,
            I => \N__28639\
        );

    \I__6687\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28636\
        );

    \I__6686\ : Span4Mux_h
    port map (
            O => \N__28651\,
            I => \N__28633\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__28646\,
            I => \N__28628\
        );

    \I__6684\ : Span4Mux_h
    port map (
            O => \N__28643\,
            I => \N__28628\
        );

    \I__6683\ : InMux
    port map (
            O => \N__28642\,
            I => \N__28625\
        );

    \I__6682\ : Span4Mux_h
    port map (
            O => \N__28639\,
            I => \N__28622\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__28636\,
            I => \N__28617\
        );

    \I__6680\ : Span4Mux_h
    port map (
            O => \N__28633\,
            I => \N__28617\
        );

    \I__6679\ : Span4Mux_h
    port map (
            O => \N__28628\,
            I => \N__28614\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__28625\,
            I => \this_ppu.N_132_0\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__28622\,
            I => \this_ppu.N_132_0\
        );

    \I__6676\ : Odrv4
    port map (
            O => \N__28617\,
            I => \this_ppu.N_132_0\
        );

    \I__6675\ : Odrv4
    port map (
            O => \N__28614\,
            I => \this_ppu.N_132_0\
        );

    \I__6674\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28602\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__28602\,
            I => \N__28599\
        );

    \I__6672\ : Span4Mux_h
    port map (
            O => \N__28599\,
            I => \N__28596\
        );

    \I__6671\ : Odrv4
    port map (
            O => \N__28596\,
            I => \N_56_0\
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__28593\,
            I => \N__28590\
        );

    \I__6669\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28587\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__28587\,
            I => \M_this_data_tmp_qZ0Z_13\
        );

    \I__6667\ : CascadeMux
    port map (
            O => \N__28584\,
            I => \N__28580\
        );

    \I__6666\ : CascadeMux
    port map (
            O => \N__28583\,
            I => \N__28576\
        );

    \I__6665\ : InMux
    port map (
            O => \N__28580\,
            I => \N__28571\
        );

    \I__6664\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28571\
        );

    \I__6663\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28568\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__28571\,
            I => \N__28562\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__28568\,
            I => \N__28562\
        );

    \I__6660\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28558\
        );

    \I__6659\ : Span4Mux_v
    port map (
            O => \N__28562\,
            I => \N__28554\
        );

    \I__6658\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28551\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__28558\,
            I => \N__28548\
        );

    \I__6656\ : InMux
    port map (
            O => \N__28557\,
            I => \N__28545\
        );

    \I__6655\ : Span4Mux_h
    port map (
            O => \N__28554\,
            I => \N__28542\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__28551\,
            I => \N__28539\
        );

    \I__6653\ : Span4Mux_h
    port map (
            O => \N__28548\,
            I => \N__28534\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__28545\,
            I => \N__28534\
        );

    \I__6651\ : Odrv4
    port map (
            O => \N__28542\,
            I => \M_this_state_d21_1\
        );

    \I__6650\ : Odrv12
    port map (
            O => \N__28539\,
            I => \M_this_state_d21_1\
        );

    \I__6649\ : Odrv4
    port map (
            O => \N__28534\,
            I => \M_this_state_d21_1\
        );

    \I__6648\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__6646\ : Span4Mux_v
    port map (
            O => \N__28521\,
            I => \N__28516\
        );

    \I__6645\ : InMux
    port map (
            O => \N__28520\,
            I => \N__28511\
        );

    \I__6644\ : InMux
    port map (
            O => \N__28519\,
            I => \N__28511\
        );

    \I__6643\ : Sp12to4
    port map (
            O => \N__28516\,
            I => \N__28506\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__28511\,
            I => \N__28506\
        );

    \I__6641\ : Odrv12
    port map (
            O => \N__28506\,
            I => port_address_in_4
        );

    \I__6640\ : InMux
    port map (
            O => \N__28503\,
            I => \N__28495\
        );

    \I__6639\ : InMux
    port map (
            O => \N__28502\,
            I => \N__28495\
        );

    \I__6638\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28490\
        );

    \I__6637\ : InMux
    port map (
            O => \N__28500\,
            I => \N__28490\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__28495\,
            I => \N__28485\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__28490\,
            I => \N__28485\
        );

    \I__6634\ : Sp12to4
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__6633\ : Odrv12
    port map (
            O => \N__28482\,
            I => port_address_in_2
        );

    \I__6632\ : CascadeMux
    port map (
            O => \N__28479\,
            I => \N__28475\
        );

    \I__6631\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28470\
        );

    \I__6630\ : InMux
    port map (
            O => \N__28475\,
            I => \N__28470\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__28470\,
            I => \N__28467\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__28467\,
            I => \M_this_state_d21_6_x\
        );

    \I__6627\ : InMux
    port map (
            O => \N__28464\,
            I => \N__28461\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__28461\,
            I => \N__28458\
        );

    \I__6625\ : Odrv4
    port map (
            O => \N__28458\,
            I => \M_this_substate_q_RNOZ0Z_2\
        );

    \I__6624\ : CascadeMux
    port map (
            O => \N__28455\,
            I => \N__28451\
        );

    \I__6623\ : InMux
    port map (
            O => \N__28454\,
            I => \N__28447\
        );

    \I__6622\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28442\
        );

    \I__6621\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28442\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__28447\,
            I => \N__28436\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__28442\,
            I => \N__28436\
        );

    \I__6618\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28433\
        );

    \I__6617\ : Span4Mux_v
    port map (
            O => \N__28436\,
            I => \N__28428\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__28433\,
            I => \N__28428\
        );

    \I__6615\ : Span4Mux_h
    port map (
            O => \N__28428\,
            I => \N__28425\
        );

    \I__6614\ : Span4Mux_v
    port map (
            O => \N__28425\,
            I => \N__28422\
        );

    \I__6613\ : Span4Mux_h
    port map (
            O => \N__28422\,
            I => \N__28419\
        );

    \I__6612\ : Odrv4
    port map (
            O => \N__28419\,
            I => port_address_in_3
        );

    \I__6611\ : CascadeMux
    port map (
            O => \N__28416\,
            I => \N__28411\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__28415\,
            I => \N__28408\
        );

    \I__6609\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28404\
        );

    \I__6608\ : InMux
    port map (
            O => \N__28411\,
            I => \N__28399\
        );

    \I__6607\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28399\
        );

    \I__6606\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28396\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__28404\,
            I => \N__28391\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__28399\,
            I => \N__28386\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__28396\,
            I => \N__28386\
        );

    \I__6602\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28383\
        );

    \I__6601\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28379\
        );

    \I__6600\ : Span4Mux_h
    port map (
            O => \N__28391\,
            I => \N__28374\
        );

    \I__6599\ : Span4Mux_h
    port map (
            O => \N__28386\,
            I => \N__28374\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__28383\,
            I => \N__28371\
        );

    \I__6597\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28368\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__28379\,
            I => \N__28365\
        );

    \I__6595\ : Span4Mux_h
    port map (
            O => \N__28374\,
            I => \N__28357\
        );

    \I__6594\ : Span4Mux_v
    port map (
            O => \N__28371\,
            I => \N__28357\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28357\
        );

    \I__6592\ : Span4Mux_v
    port map (
            O => \N__28365\,
            I => \N__28354\
        );

    \I__6591\ : InMux
    port map (
            O => \N__28364\,
            I => \N__28351\
        );

    \I__6590\ : Span4Mux_h
    port map (
            O => \N__28357\,
            I => \N__28348\
        );

    \I__6589\ : Sp12to4
    port map (
            O => \N__28354\,
            I => \N__28343\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__28351\,
            I => \N__28343\
        );

    \I__6587\ : Span4Mux_v
    port map (
            O => \N__28348\,
            I => \N__28340\
        );

    \I__6586\ : Span12Mux_h
    port map (
            O => \N__28343\,
            I => \N__28337\
        );

    \I__6585\ : Span4Mux_v
    port map (
            O => \N__28340\,
            I => \N__28334\
        );

    \I__6584\ : Odrv12
    port map (
            O => \N__28337\,
            I => port_address_in_1
        );

    \I__6583\ : Odrv4
    port map (
            O => \N__28334\,
            I => port_address_in_1
        );

    \I__6582\ : CascadeMux
    port map (
            O => \N__28329\,
            I => \N__28326\
        );

    \I__6581\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28323\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__28323\,
            I => \N__28320\
        );

    \I__6579\ : Span4Mux_v
    port map (
            O => \N__28320\,
            I => \N__28317\
        );

    \I__6578\ : Odrv4
    port map (
            O => \N__28317\,
            I => \this_vga_signals.M_this_state_d24Z0Z_1\
        );

    \I__6577\ : CEMux
    port map (
            O => \N__28314\,
            I => \N__28310\
        );

    \I__6576\ : CEMux
    port map (
            O => \N__28313\,
            I => \N__28307\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__28310\,
            I => \N__28304\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__28307\,
            I => \N__28301\
        );

    \I__6573\ : Span4Mux_h
    port map (
            O => \N__28304\,
            I => \N__28298\
        );

    \I__6572\ : Span4Mux_h
    port map (
            O => \N__28301\,
            I => \N__28295\
        );

    \I__6571\ : Span4Mux_v
    port map (
            O => \N__28298\,
            I => \N__28292\
        );

    \I__6570\ : Span4Mux_v
    port map (
            O => \N__28295\,
            I => \N__28289\
        );

    \I__6569\ : Odrv4
    port map (
            O => \N__28292\,
            I => \this_sprites_ram.mem_WE_0\
        );

    \I__6568\ : Odrv4
    port map (
            O => \N__28289\,
            I => \this_sprites_ram.mem_WE_0\
        );

    \I__6567\ : CascadeMux
    port map (
            O => \N__28284\,
            I => \N__28280\
        );

    \I__6566\ : InMux
    port map (
            O => \N__28283\,
            I => \N__28277\
        );

    \I__6565\ : InMux
    port map (
            O => \N__28280\,
            I => \N__28274\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__28277\,
            I => \this_ppu.M_this_ppu_map_addr_i_1\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__28274\,
            I => \this_ppu.M_this_ppu_map_addr_i_1\
        );

    \I__6562\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28265\
        );

    \I__6561\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28262\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__28265\,
            I => \this_ppu.M_this_ppu_map_addr_i_2\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__28262\,
            I => \this_ppu.M_this_ppu_map_addr_i_2\
        );

    \I__6558\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28253\
        );

    \I__6557\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28250\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__28253\,
            I => \this_ppu.M_this_ppu_map_addr_i_3\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__28250\,
            I => \this_ppu.M_this_ppu_map_addr_i_3\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__28245\,
            I => \N__28242\
        );

    \I__6553\ : InMux
    port map (
            O => \N__28242\,
            I => \N__28238\
        );

    \I__6552\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28235\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__28238\,
            I => \this_ppu.M_this_ppu_map_addr_i_4\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__28235\,
            I => \this_ppu.M_this_ppu_map_addr_i_4\
        );

    \I__6549\ : InMux
    port map (
            O => \N__28230\,
            I => \bfn_22_20_0_\
        );

    \I__6548\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28224\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__28224\,
            I => \this_ppu.vscroll8_1\
        );

    \I__6546\ : InMux
    port map (
            O => \N__28221\,
            I => \N__28218\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__28218\,
            I => \N__28215\
        );

    \I__6544\ : Span4Mux_h
    port map (
            O => \N__28215\,
            I => \N__28211\
        );

    \I__6543\ : InMux
    port map (
            O => \N__28214\,
            I => \N__28208\
        );

    \I__6542\ : Span4Mux_h
    port map (
            O => \N__28211\,
            I => \N__28205\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__28208\,
            I => \N__28202\
        );

    \I__6540\ : IoSpan4Mux
    port map (
            O => \N__28205\,
            I => \N__28199\
        );

    \I__6539\ : Span12Mux_h
    port map (
            O => \N__28202\,
            I => \N__28196\
        );

    \I__6538\ : Odrv4
    port map (
            O => \N__28199\,
            I => port_address_in_5
        );

    \I__6537\ : Odrv12
    port map (
            O => \N__28196\,
            I => port_address_in_5
        );

    \I__6536\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28188\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__28188\,
            I => \N__28184\
        );

    \I__6534\ : InMux
    port map (
            O => \N__28187\,
            I => \N__28181\
        );

    \I__6533\ : Span4Mux_h
    port map (
            O => \N__28184\,
            I => \N__28176\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__28181\,
            I => \N__28176\
        );

    \I__6531\ : Span4Mux_v
    port map (
            O => \N__28176\,
            I => \N__28173\
        );

    \I__6530\ : Sp12to4
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__6529\ : Odrv12
    port map (
            O => \N__28170\,
            I => port_address_in_6
        );

    \I__6528\ : CascadeMux
    port map (
            O => \N__28167\,
            I => \N__28164\
        );

    \I__6527\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28161\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__28161\,
            I => \N__28157\
        );

    \I__6525\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28154\
        );

    \I__6524\ : Span4Mux_v
    port map (
            O => \N__28157\,
            I => \N__28151\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__28154\,
            I => \N__28148\
        );

    \I__6522\ : Sp12to4
    port map (
            O => \N__28151\,
            I => \N__28143\
        );

    \I__6521\ : Span12Mux_v
    port map (
            O => \N__28148\,
            I => \N__28143\
        );

    \I__6520\ : Span12Mux_v
    port map (
            O => \N__28143\,
            I => \N__28140\
        );

    \I__6519\ : Odrv12
    port map (
            O => \N__28140\,
            I => port_address_in_7
        );

    \I__6518\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28134\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__28134\,
            I => \N__28130\
        );

    \I__6516\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28127\
        );

    \I__6515\ : Span4Mux_h
    port map (
            O => \N__28130\,
            I => \N__28121\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__28127\,
            I => \N__28121\
        );

    \I__6513\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28115\
        );

    \I__6512\ : Span4Mux_h
    port map (
            O => \N__28121\,
            I => \N__28112\
        );

    \I__6511\ : InMux
    port map (
            O => \N__28120\,
            I => \N__28109\
        );

    \I__6510\ : InMux
    port map (
            O => \N__28119\,
            I => \N__28106\
        );

    \I__6509\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28103\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__28115\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6507\ : Odrv4
    port map (
            O => \N__28112\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__28109\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__28106\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__28103\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6503\ : InMux
    port map (
            O => \N__28092\,
            I => \bfn_22_18_0_\
        );

    \I__6502\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28086\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__28086\,
            I => \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO\
        );

    \I__6500\ : CascadeMux
    port map (
            O => \N__28083\,
            I => \N__28080\
        );

    \I__6499\ : InMux
    port map (
            O => \N__28080\,
            I => \N__28077\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__28077\,
            I => \N__28074\
        );

    \I__6497\ : Odrv4
    port map (
            O => \N__28074\,
            I => \this_ppu.un1_M_haddress_q_2_5\
        );

    \I__6496\ : CascadeMux
    port map (
            O => \N__28071\,
            I => \un1_M_this_oam_address_q_c3_cascade_\
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__28068\,
            I => \N__28065\
        );

    \I__6494\ : InMux
    port map (
            O => \N__28065\,
            I => \N__28062\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__28062\,
            I => \N__28059\
        );

    \I__6492\ : Odrv12
    port map (
            O => \N__28059\,
            I => \M_this_data_tmp_qZ0Z_7\
        );

    \I__6491\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28053\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28050\
        );

    \I__6489\ : Span4Mux_h
    port map (
            O => \N__28050\,
            I => \N__28047\
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__28047\,
            I => \N_65_0\
        );

    \I__6487\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28040\
        );

    \I__6486\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28037\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__28040\,
            I => \this_ppu.M_this_ppu_vram_addr_i_0\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__28037\,
            I => \this_ppu.M_this_ppu_vram_addr_i_0\
        );

    \I__6483\ : CascadeMux
    port map (
            O => \N__28032\,
            I => \N__28027\
        );

    \I__6482\ : InMux
    port map (
            O => \N__28031\,
            I => \N__28023\
        );

    \I__6481\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28020\
        );

    \I__6480\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28017\
        );

    \I__6479\ : CascadeMux
    port map (
            O => \N__28026\,
            I => \N__28014\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__28023\,
            I => \N__28007\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__28020\,
            I => \N__28007\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__28017\,
            I => \N__28007\
        );

    \I__6475\ : InMux
    port map (
            O => \N__28014\,
            I => \N__28004\
        );

    \I__6474\ : Span4Mux_v
    port map (
            O => \N__28007\,
            I => \N__27999\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__28004\,
            I => \N__27999\
        );

    \I__6472\ : Span4Mux_h
    port map (
            O => \N__27999\,
            I => \N__27996\
        );

    \I__6471\ : Odrv4
    port map (
            O => \N__27996\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__6470\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27989\
        );

    \I__6469\ : InMux
    port map (
            O => \N__27992\,
            I => \N__27986\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__27989\,
            I => \this_ppu.M_this_ppu_vram_addr_i_1\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__27986\,
            I => \this_ppu.M_this_ppu_vram_addr_i_1\
        );

    \I__6466\ : CascadeMux
    port map (
            O => \N__27981\,
            I => \N__27977\
        );

    \I__6465\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27973\
        );

    \I__6464\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27970\
        );

    \I__6463\ : CascadeMux
    port map (
            O => \N__27976\,
            I => \N__27967\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__27973\,
            I => \N__27962\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__27970\,
            I => \N__27962\
        );

    \I__6460\ : InMux
    port map (
            O => \N__27967\,
            I => \N__27959\
        );

    \I__6459\ : Span4Mux_v
    port map (
            O => \N__27962\,
            I => \N__27954\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__27959\,
            I => \N__27954\
        );

    \I__6457\ : Span4Mux_h
    port map (
            O => \N__27954\,
            I => \N__27951\
        );

    \I__6456\ : Odrv4
    port map (
            O => \N__27951\,
            I => \M_this_oam_ram_read_data_9\
        );

    \I__6455\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27944\
        );

    \I__6454\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27941\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__27944\,
            I => \this_ppu.M_this_ppu_vram_addr_i_2\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__27941\,
            I => \this_ppu.M_this_ppu_vram_addr_i_2\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__27936\,
            I => \N__27933\
        );

    \I__6450\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27928\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__27932\,
            I => \N__27925\
        );

    \I__6448\ : InMux
    port map (
            O => \N__27931\,
            I => \N__27922\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__27928\,
            I => \N__27919\
        );

    \I__6446\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27916\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__27922\,
            I => \N__27913\
        );

    \I__6444\ : Span4Mux_v
    port map (
            O => \N__27919\,
            I => \N__27908\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__27916\,
            I => \N__27908\
        );

    \I__6442\ : Span4Mux_h
    port map (
            O => \N__27913\,
            I => \N__27905\
        );

    \I__6441\ : Span4Mux_h
    port map (
            O => \N__27908\,
            I => \N__27902\
        );

    \I__6440\ : Odrv4
    port map (
            O => \N__27905\,
            I => \M_this_oam_ram_read_data_10\
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__27902\,
            I => \M_this_oam_ram_read_data_10\
        );

    \I__6438\ : CascadeMux
    port map (
            O => \N__27897\,
            I => \N__27893\
        );

    \I__6437\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27890\
        );

    \I__6436\ : InMux
    port map (
            O => \N__27893\,
            I => \N__27887\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__27890\,
            I => \this_ppu.M_this_ppu_map_addr_i_0\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__27887\,
            I => \this_ppu.M_this_ppu_map_addr_i_0\
        );

    \I__6433\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27873\
        );

    \I__6432\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27873\
        );

    \I__6431\ : InMux
    port map (
            O => \N__27880\,
            I => \N__27873\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__27873\,
            I => \this_ppu.un1_M_vaddress_q_2_c5\
        );

    \I__6429\ : CascadeMux
    port map (
            O => \N__27870\,
            I => \N__27867\
        );

    \I__6428\ : CascadeBuf
    port map (
            O => \N__27867\,
            I => \N__27864\
        );

    \I__6427\ : CascadeMux
    port map (
            O => \N__27864\,
            I => \N__27861\
        );

    \I__6426\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27858\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27854\
        );

    \I__6424\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27848\
        );

    \I__6423\ : Span12Mux_h
    port map (
            O => \N__27854\,
            I => \N__27845\
        );

    \I__6422\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27838\
        );

    \I__6421\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27838\
        );

    \I__6420\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27838\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__27848\,
            I => \N__27835\
        );

    \I__6418\ : Span12Mux_v
    port map (
            O => \N__27845\,
            I => \N__27832\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__27838\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__6416\ : Odrv4
    port map (
            O => \N__27835\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__6415\ : Odrv12
    port map (
            O => \N__27832\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__27825\,
            I => \N__27822\
        );

    \I__6413\ : CascadeBuf
    port map (
            O => \N__27822\,
            I => \N__27819\
        );

    \I__6412\ : CascadeMux
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__6411\ : InMux
    port map (
            O => \N__27816\,
            I => \N__27813\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__27813\,
            I => \N__27810\
        );

    \I__6409\ : Sp12to4
    port map (
            O => \N__27810\,
            I => \N__27805\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__27809\,
            I => \N__27802\
        );

    \I__6407\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27798\
        );

    \I__6406\ : Span12Mux_h
    port map (
            O => \N__27805\,
            I => \N__27795\
        );

    \I__6405\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27790\
        );

    \I__6404\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27790\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__27798\,
            I => \N__27787\
        );

    \I__6402\ : Span12Mux_v
    port map (
            O => \N__27795\,
            I => \N__27784\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__27790\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__6400\ : Odrv4
    port map (
            O => \N__27787\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__6399\ : Odrv12
    port map (
            O => \N__27784\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__27777\,
            I => \N__27774\
        );

    \I__6397\ : CascadeBuf
    port map (
            O => \N__27774\,
            I => \N__27771\
        );

    \I__6396\ : CascadeMux
    port map (
            O => \N__27771\,
            I => \N__27768\
        );

    \I__6395\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__27765\,
            I => \N__27761\
        );

    \I__6393\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27757\
        );

    \I__6392\ : Span12Mux_h
    port map (
            O => \N__27761\,
            I => \N__27754\
        );

    \I__6391\ : InMux
    port map (
            O => \N__27760\,
            I => \N__27751\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__27757\,
            I => \N__27748\
        );

    \I__6389\ : Span12Mux_v
    port map (
            O => \N__27754\,
            I => \N__27745\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__27751\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__6387\ : Odrv4
    port map (
            O => \N__27748\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__6386\ : Odrv12
    port map (
            O => \N__27745\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__6385\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27735\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27732\
        );

    \I__6383\ : Odrv4
    port map (
            O => \N__27732\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4\
        );

    \I__6382\ : InMux
    port map (
            O => \N__27729\,
            I => \N__27716\
        );

    \I__6381\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27716\
        );

    \I__6380\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27707\
        );

    \I__6379\ : InMux
    port map (
            O => \N__27726\,
            I => \N__27707\
        );

    \I__6378\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27707\
        );

    \I__6377\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27707\
        );

    \I__6376\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27704\
        );

    \I__6375\ : InMux
    port map (
            O => \N__27722\,
            I => \N__27697\
        );

    \I__6374\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27697\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__27716\,
            I => \N__27692\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__27707\,
            I => \N__27692\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27689\
        );

    \I__6370\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27686\
        );

    \I__6369\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27680\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__27697\,
            I => \N__27677\
        );

    \I__6367\ : Span4Mux_v
    port map (
            O => \N__27692\,
            I => \N__27670\
        );

    \I__6366\ : Span4Mux_h
    port map (
            O => \N__27689\,
            I => \N__27670\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__27686\,
            I => \N__27670\
        );

    \I__6364\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27663\
        );

    \I__6363\ : InMux
    port map (
            O => \N__27684\,
            I => \N__27663\
        );

    \I__6362\ : InMux
    port map (
            O => \N__27683\,
            I => \N__27663\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__27680\,
            I => \this_vga_signals.un1_M_this_state_q_14_0\
        );

    \I__6360\ : Odrv4
    port map (
            O => \N__27677\,
            I => \this_vga_signals.un1_M_this_state_q_14_0\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__27670\,
            I => \this_vga_signals.un1_M_this_state_q_14_0\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__27663\,
            I => \this_vga_signals.un1_M_this_state_q_14_0\
        );

    \I__6357\ : CascadeMux
    port map (
            O => \N__27654\,
            I => \N__27651\
        );

    \I__6356\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27648\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__27648\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_4\
        );

    \I__6354\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27642\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__27642\,
            I => \N__27639\
        );

    \I__6352\ : Span4Mux_h
    port map (
            O => \N__27639\,
            I => \N__27636\
        );

    \I__6351\ : Odrv4
    port map (
            O => \N__27636\,
            I => \un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0\
        );

    \I__6350\ : CascadeMux
    port map (
            O => \N__27633\,
            I => \N__27630\
        );

    \I__6349\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27626\
        );

    \I__6348\ : CascadeMux
    port map (
            O => \N__27629\,
            I => \N__27623\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__27626\,
            I => \N__27619\
        );

    \I__6346\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27616\
        );

    \I__6345\ : CascadeMux
    port map (
            O => \N__27622\,
            I => \N__27613\
        );

    \I__6344\ : Span4Mux_h
    port map (
            O => \N__27619\,
            I => \N__27606\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__27616\,
            I => \N__27606\
        );

    \I__6342\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27603\
        );

    \I__6341\ : CascadeMux
    port map (
            O => \N__27612\,
            I => \N__27600\
        );

    \I__6340\ : CascadeMux
    port map (
            O => \N__27611\,
            I => \N__27596\
        );

    \I__6339\ : Span4Mux_v
    port map (
            O => \N__27606\,
            I => \N__27591\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__27603\,
            I => \N__27591\
        );

    \I__6337\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27588\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__27599\,
            I => \N__27585\
        );

    \I__6335\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27581\
        );

    \I__6334\ : Span4Mux_h
    port map (
            O => \N__27591\,
            I => \N__27575\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27575\
        );

    \I__6332\ : InMux
    port map (
            O => \N__27585\,
            I => \N__27572\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__27584\,
            I => \N__27569\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__27581\,
            I => \N__27565\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__27580\,
            I => \N__27562\
        );

    \I__6328\ : Span4Mux_v
    port map (
            O => \N__27575\,
            I => \N__27556\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__27572\,
            I => \N__27556\
        );

    \I__6326\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27553\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__27568\,
            I => \N__27550\
        );

    \I__6324\ : Span4Mux_h
    port map (
            O => \N__27565\,
            I => \N__27545\
        );

    \I__6323\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27542\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__27561\,
            I => \N__27539\
        );

    \I__6321\ : Span4Mux_h
    port map (
            O => \N__27556\,
            I => \N__27533\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__27553\,
            I => \N__27533\
        );

    \I__6319\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27530\
        );

    \I__6318\ : CascadeMux
    port map (
            O => \N__27549\,
            I => \N__27526\
        );

    \I__6317\ : CascadeMux
    port map (
            O => \N__27548\,
            I => \N__27523\
        );

    \I__6316\ : Span4Mux_v
    port map (
            O => \N__27545\,
            I => \N__27517\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__27542\,
            I => \N__27517\
        );

    \I__6314\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27514\
        );

    \I__6313\ : CascadeMux
    port map (
            O => \N__27538\,
            I => \N__27511\
        );

    \I__6312\ : Span4Mux_v
    port map (
            O => \N__27533\,
            I => \N__27506\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__27530\,
            I => \N__27506\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__27529\,
            I => \N__27503\
        );

    \I__6309\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27500\
        );

    \I__6308\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27497\
        );

    \I__6307\ : CascadeMux
    port map (
            O => \N__27522\,
            I => \N__27494\
        );

    \I__6306\ : Span4Mux_h
    port map (
            O => \N__27517\,
            I => \N__27488\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__27514\,
            I => \N__27488\
        );

    \I__6304\ : InMux
    port map (
            O => \N__27511\,
            I => \N__27485\
        );

    \I__6303\ : Span4Mux_h
    port map (
            O => \N__27506\,
            I => \N__27482\
        );

    \I__6302\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27479\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__27500\,
            I => \N__27476\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__27497\,
            I => \N__27473\
        );

    \I__6299\ : InMux
    port map (
            O => \N__27494\,
            I => \N__27470\
        );

    \I__6298\ : CascadeMux
    port map (
            O => \N__27493\,
            I => \N__27467\
        );

    \I__6297\ : Span4Mux_v
    port map (
            O => \N__27488\,
            I => \N__27461\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__27485\,
            I => \N__27461\
        );

    \I__6295\ : Span4Mux_v
    port map (
            O => \N__27482\,
            I => \N__27456\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__27479\,
            I => \N__27456\
        );

    \I__6293\ : Span4Mux_v
    port map (
            O => \N__27476\,
            I => \N__27449\
        );

    \I__6292\ : Span4Mux_h
    port map (
            O => \N__27473\,
            I => \N__27449\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__27470\,
            I => \N__27449\
        );

    \I__6290\ : InMux
    port map (
            O => \N__27467\,
            I => \N__27446\
        );

    \I__6289\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27442\
        );

    \I__6288\ : Sp12to4
    port map (
            O => \N__27461\,
            I => \N__27438\
        );

    \I__6287\ : Span4Mux_v
    port map (
            O => \N__27456\,
            I => \N__27431\
        );

    \I__6286\ : Span4Mux_v
    port map (
            O => \N__27449\,
            I => \N__27431\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__27446\,
            I => \N__27431\
        );

    \I__6284\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27428\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27425\
        );

    \I__6282\ : InMux
    port map (
            O => \N__27441\,
            I => \N__27422\
        );

    \I__6281\ : Span12Mux_h
    port map (
            O => \N__27438\,
            I => \N__27415\
        );

    \I__6280\ : Sp12to4
    port map (
            O => \N__27431\,
            I => \N__27415\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__27428\,
            I => \N__27415\
        );

    \I__6278\ : Span4Mux_h
    port map (
            O => \N__27425\,
            I => \N__27412\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__27422\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__6276\ : Odrv12
    port map (
            O => \N__27415\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__6275\ : Odrv4
    port map (
            O => \N__27412\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__6274\ : InMux
    port map (
            O => \N__27405\,
            I => \N__27401\
        );

    \I__6273\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27396\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__27401\,
            I => \N__27393\
        );

    \I__6271\ : InMux
    port map (
            O => \N__27400\,
            I => \N__27390\
        );

    \I__6270\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27387\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__27396\,
            I => \N__27384\
        );

    \I__6268\ : Span4Mux_v
    port map (
            O => \N__27393\,
            I => \N__27379\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__27390\,
            I => \N__27379\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__27387\,
            I => \N__27376\
        );

    \I__6265\ : Odrv4
    port map (
            O => \N__27384\,
            I => \this_vga_signals.M_this_state_q_ns_8\
        );

    \I__6264\ : Odrv4
    port map (
            O => \N__27379\,
            I => \this_vga_signals.M_this_state_q_ns_8\
        );

    \I__6263\ : Odrv4
    port map (
            O => \N__27376\,
            I => \this_vga_signals.M_this_state_q_ns_8\
        );

    \I__6262\ : InMux
    port map (
            O => \N__27369\,
            I => \N__27365\
        );

    \I__6261\ : InMux
    port map (
            O => \N__27368\,
            I => \N__27362\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__27365\,
            I => \N__27357\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27354\
        );

    \I__6258\ : InMux
    port map (
            O => \N__27361\,
            I => \N__27351\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__27360\,
            I => \N__27347\
        );

    \I__6256\ : Span4Mux_h
    port map (
            O => \N__27357\,
            I => \N__27344\
        );

    \I__6255\ : Span4Mux_v
    port map (
            O => \N__27354\,
            I => \N__27341\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__27351\,
            I => \N__27338\
        );

    \I__6253\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27335\
        );

    \I__6252\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27332\
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__27344\,
            I => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\
        );

    \I__6250\ : Odrv4
    port map (
            O => \N__27341\,
            I => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\
        );

    \I__6249\ : Odrv12
    port map (
            O => \N__27338\,
            I => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__27335\,
            I => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__27332\,
            I => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\
        );

    \I__6246\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27318\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__27318\,
            I => \N__27313\
        );

    \I__6244\ : InMux
    port map (
            O => \N__27317\,
            I => \N__27310\
        );

    \I__6243\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27306\
        );

    \I__6242\ : Span4Mux_h
    port map (
            O => \N__27313\,
            I => \N__27302\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__27310\,
            I => \N__27299\
        );

    \I__6240\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27296\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__27306\,
            I => \N__27292\
        );

    \I__6238\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27289\
        );

    \I__6237\ : Span4Mux_v
    port map (
            O => \N__27302\,
            I => \N__27284\
        );

    \I__6236\ : Span4Mux_h
    port map (
            O => \N__27299\,
            I => \N__27284\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__27296\,
            I => \N__27281\
        );

    \I__6234\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27278\
        );

    \I__6233\ : Span4Mux_v
    port map (
            O => \N__27292\,
            I => \N__27273\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__27289\,
            I => \N__27273\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__27284\,
            I => \N__27268\
        );

    \I__6230\ : Span4Mux_h
    port map (
            O => \N__27281\,
            I => \N__27268\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__27278\,
            I => \N__27265\
        );

    \I__6228\ : Span4Mux_v
    port map (
            O => \N__27273\,
            I => \N__27260\
        );

    \I__6227\ : Span4Mux_v
    port map (
            O => \N__27268\,
            I => \N__27255\
        );

    \I__6226\ : Span4Mux_h
    port map (
            O => \N__27265\,
            I => \N__27255\
        );

    \I__6225\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27252\
        );

    \I__6224\ : InMux
    port map (
            O => \N__27263\,
            I => \N__27249\
        );

    \I__6223\ : Span4Mux_h
    port map (
            O => \N__27260\,
            I => \N__27246\
        );

    \I__6222\ : Span4Mux_v
    port map (
            O => \N__27255\,
            I => \N__27243\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__27252\,
            I => \N__27240\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__27249\,
            I => \N__27237\
        );

    \I__6219\ : Sp12to4
    port map (
            O => \N__27246\,
            I => \N__27234\
        );

    \I__6218\ : Span4Mux_v
    port map (
            O => \N__27243\,
            I => \N__27227\
        );

    \I__6217\ : Span4Mux_h
    port map (
            O => \N__27240\,
            I => \N__27227\
        );

    \I__6216\ : Span4Mux_h
    port map (
            O => \N__27237\,
            I => \N__27227\
        );

    \I__6215\ : Odrv12
    port map (
            O => \N__27234\,
            I => \M_this_sprites_ram_write_data_1\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__27227\,
            I => \M_this_sprites_ram_write_data_1\
        );

    \I__6213\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27219\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__27219\,
            I => \N__27216\
        );

    \I__6211\ : Span12Mux_v
    port map (
            O => \N__27216\,
            I => \N__27213\
        );

    \I__6210\ : Span12Mux_h
    port map (
            O => \N__27213\,
            I => \N__27210\
        );

    \I__6209\ : Span12Mux_v
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__6208\ : Odrv12
    port map (
            O => \N__27207\,
            I => \M_this_map_ram_read_data_4\
        );

    \I__6207\ : CascadeMux
    port map (
            O => \N__27204\,
            I => \N__27197\
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__27203\,
            I => \N__27193\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__27202\,
            I => \N__27190\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__27201\,
            I => \N__27186\
        );

    \I__6203\ : CascadeMux
    port map (
            O => \N__27200\,
            I => \N__27183\
        );

    \I__6202\ : InMux
    port map (
            O => \N__27197\,
            I => \N__27179\
        );

    \I__6201\ : CascadeMux
    port map (
            O => \N__27196\,
            I => \N__27176\
        );

    \I__6200\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27172\
        );

    \I__6199\ : InMux
    port map (
            O => \N__27190\,
            I => \N__27169\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__27189\,
            I => \N__27166\
        );

    \I__6197\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27161\
        );

    \I__6196\ : InMux
    port map (
            O => \N__27183\,
            I => \N__27158\
        );

    \I__6195\ : CascadeMux
    port map (
            O => \N__27182\,
            I => \N__27155\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__27179\,
            I => \N__27151\
        );

    \I__6193\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27148\
        );

    \I__6192\ : CascadeMux
    port map (
            O => \N__27175\,
            I => \N__27145\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__27172\,
            I => \N__27141\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__27169\,
            I => \N__27138\
        );

    \I__6189\ : InMux
    port map (
            O => \N__27166\,
            I => \N__27135\
        );

    \I__6188\ : CascadeMux
    port map (
            O => \N__27165\,
            I => \N__27132\
        );

    \I__6187\ : CascadeMux
    port map (
            O => \N__27164\,
            I => \N__27128\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__27161\,
            I => \N__27123\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__27158\,
            I => \N__27123\
        );

    \I__6184\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27120\
        );

    \I__6183\ : CascadeMux
    port map (
            O => \N__27154\,
            I => \N__27116\
        );

    \I__6182\ : Span4Mux_v
    port map (
            O => \N__27151\,
            I => \N__27111\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__27148\,
            I => \N__27111\
        );

    \I__6180\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27108\
        );

    \I__6179\ : CascadeMux
    port map (
            O => \N__27144\,
            I => \N__27105\
        );

    \I__6178\ : Span4Mux_v
    port map (
            O => \N__27141\,
            I => \N__27098\
        );

    \I__6177\ : Span4Mux_h
    port map (
            O => \N__27138\,
            I => \N__27098\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__27135\,
            I => \N__27098\
        );

    \I__6175\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27095\
        );

    \I__6174\ : CascadeMux
    port map (
            O => \N__27131\,
            I => \N__27092\
        );

    \I__6173\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27089\
        );

    \I__6172\ : Span4Mux_v
    port map (
            O => \N__27123\,
            I => \N__27084\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__27120\,
            I => \N__27084\
        );

    \I__6170\ : CascadeMux
    port map (
            O => \N__27119\,
            I => \N__27081\
        );

    \I__6169\ : InMux
    port map (
            O => \N__27116\,
            I => \N__27077\
        );

    \I__6168\ : Span4Mux_h
    port map (
            O => \N__27111\,
            I => \N__27072\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__27108\,
            I => \N__27072\
        );

    \I__6166\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27069\
        );

    \I__6165\ : Span4Mux_v
    port map (
            O => \N__27098\,
            I => \N__27064\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__27095\,
            I => \N__27064\
        );

    \I__6163\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27061\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__27089\,
            I => \N__27058\
        );

    \I__6161\ : Span4Mux_v
    port map (
            O => \N__27084\,
            I => \N__27055\
        );

    \I__6160\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27052\
        );

    \I__6159\ : CascadeMux
    port map (
            O => \N__27080\,
            I => \N__27049\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__27077\,
            I => \N__27046\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__27072\,
            I => \N__27041\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__27069\,
            I => \N__27041\
        );

    \I__6155\ : Span4Mux_h
    port map (
            O => \N__27064\,
            I => \N__27038\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__27061\,
            I => \N__27035\
        );

    \I__6153\ : Span12Mux_h
    port map (
            O => \N__27058\,
            I => \N__27032\
        );

    \I__6152\ : Sp12to4
    port map (
            O => \N__27055\,
            I => \N__27027\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__27052\,
            I => \N__27027\
        );

    \I__6150\ : InMux
    port map (
            O => \N__27049\,
            I => \N__27024\
        );

    \I__6149\ : Span12Mux_s10_h
    port map (
            O => \N__27046\,
            I => \N__27021\
        );

    \I__6148\ : Span4Mux_h
    port map (
            O => \N__27041\,
            I => \N__27018\
        );

    \I__6147\ : Span4Mux_v
    port map (
            O => \N__27038\,
            I => \N__27013\
        );

    \I__6146\ : Span4Mux_h
    port map (
            O => \N__27035\,
            I => \N__27013\
        );

    \I__6145\ : Span12Mux_v
    port map (
            O => \N__27032\,
            I => \N__27006\
        );

    \I__6144\ : Span12Mux_h
    port map (
            O => \N__27027\,
            I => \N__27006\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__27006\
        );

    \I__6142\ : Odrv12
    port map (
            O => \N__27021\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__6141\ : Odrv4
    port map (
            O => \N__27018\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__6140\ : Odrv4
    port map (
            O => \N__27013\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__6139\ : Odrv12
    port map (
            O => \N__27006\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__6138\ : CascadeMux
    port map (
            O => \N__26997\,
            I => \N__26993\
        );

    \I__6137\ : CascadeMux
    port map (
            O => \N__26996\,
            I => \N__26987\
        );

    \I__6136\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26982\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__26992\,
            I => \N__26979\
        );

    \I__6134\ : CascadeMux
    port map (
            O => \N__26991\,
            I => \N__26974\
        );

    \I__6133\ : CascadeMux
    port map (
            O => \N__26990\,
            I => \N__26971\
        );

    \I__6132\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26967\
        );

    \I__6131\ : CascadeMux
    port map (
            O => \N__26986\,
            I => \N__26964\
        );

    \I__6130\ : CascadeMux
    port map (
            O => \N__26985\,
            I => \N__26961\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__26982\,
            I => \N__26957\
        );

    \I__6128\ : InMux
    port map (
            O => \N__26979\,
            I => \N__26954\
        );

    \I__6127\ : CascadeMux
    port map (
            O => \N__26978\,
            I => \N__26951\
        );

    \I__6126\ : CascadeMux
    port map (
            O => \N__26977\,
            I => \N__26948\
        );

    \I__6125\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26943\
        );

    \I__6124\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26940\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__26970\,
            I => \N__26937\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__26967\,
            I => \N__26934\
        );

    \I__6121\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26931\
        );

    \I__6120\ : InMux
    port map (
            O => \N__26961\,
            I => \N__26928\
        );

    \I__6119\ : CascadeMux
    port map (
            O => \N__26960\,
            I => \N__26925\
        );

    \I__6118\ : Span4Mux_h
    port map (
            O => \N__26957\,
            I => \N__26920\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__26954\,
            I => \N__26920\
        );

    \I__6116\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26917\
        );

    \I__6115\ : InMux
    port map (
            O => \N__26948\,
            I => \N__26914\
        );

    \I__6114\ : CascadeMux
    port map (
            O => \N__26947\,
            I => \N__26911\
        );

    \I__6113\ : CascadeMux
    port map (
            O => \N__26946\,
            I => \N__26908\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__26943\,
            I => \N__26904\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__26940\,
            I => \N__26901\
        );

    \I__6110\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26898\
        );

    \I__6109\ : Span4Mux_v
    port map (
            O => \N__26934\,
            I => \N__26892\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__26931\,
            I => \N__26892\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__26928\,
            I => \N__26889\
        );

    \I__6106\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26886\
        );

    \I__6105\ : Span4Mux_v
    port map (
            O => \N__26920\,
            I => \N__26879\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__26917\,
            I => \N__26879\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__26914\,
            I => \N__26879\
        );

    \I__6102\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26876\
        );

    \I__6101\ : InMux
    port map (
            O => \N__26908\,
            I => \N__26873\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__26907\,
            I => \N__26870\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__26904\,
            I => \N__26863\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__26901\,
            I => \N__26863\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__26898\,
            I => \N__26863\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__26897\,
            I => \N__26860\
        );

    \I__6095\ : Span4Mux_h
    port map (
            O => \N__26892\,
            I => \N__26856\
        );

    \I__6094\ : Span4Mux_v
    port map (
            O => \N__26889\,
            I => \N__26851\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__26886\,
            I => \N__26851\
        );

    \I__6092\ : Span4Mux_v
    port map (
            O => \N__26879\,
            I => \N__26846\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__26876\,
            I => \N__26846\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__26873\,
            I => \N__26843\
        );

    \I__6089\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26840\
        );

    \I__6088\ : Span4Mux_v
    port map (
            O => \N__26863\,
            I => \N__26837\
        );

    \I__6087\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26834\
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__26859\,
            I => \N__26831\
        );

    \I__6085\ : Span4Mux_v
    port map (
            O => \N__26856\,
            I => \N__26826\
        );

    \I__6084\ : Span4Mux_h
    port map (
            O => \N__26851\,
            I => \N__26826\
        );

    \I__6083\ : Span4Mux_h
    port map (
            O => \N__26846\,
            I => \N__26823\
        );

    \I__6082\ : Span4Mux_v
    port map (
            O => \N__26843\,
            I => \N__26818\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26818\
        );

    \I__6080\ : Sp12to4
    port map (
            O => \N__26837\,
            I => \N__26813\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__26834\,
            I => \N__26813\
        );

    \I__6078\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26810\
        );

    \I__6077\ : Span4Mux_v
    port map (
            O => \N__26826\,
            I => \N__26803\
        );

    \I__6076\ : Span4Mux_v
    port map (
            O => \N__26823\,
            I => \N__26803\
        );

    \I__6075\ : Span4Mux_h
    port map (
            O => \N__26818\,
            I => \N__26803\
        );

    \I__6074\ : Span12Mux_h
    port map (
            O => \N__26813\,
            I => \N__26798\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__26810\,
            I => \N__26798\
        );

    \I__6072\ : Odrv4
    port map (
            O => \N__26803\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__6071\ : Odrv12
    port map (
            O => \N__26798\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__6070\ : CEMux
    port map (
            O => \N__26793\,
            I => \N__26790\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__6068\ : Span4Mux_v
    port map (
            O => \N__26787\,
            I => \N__26783\
        );

    \I__6067\ : CEMux
    port map (
            O => \N__26786\,
            I => \N__26780\
        );

    \I__6066\ : Span4Mux_h
    port map (
            O => \N__26783\,
            I => \N__26777\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__26780\,
            I => \N__26774\
        );

    \I__6064\ : Span4Mux_h
    port map (
            O => \N__26777\,
            I => \N__26771\
        );

    \I__6063\ : Span4Mux_v
    port map (
            O => \N__26774\,
            I => \N__26768\
        );

    \I__6062\ : Span4Mux_h
    port map (
            O => \N__26771\,
            I => \N__26763\
        );

    \I__6061\ : Span4Mux_h
    port map (
            O => \N__26768\,
            I => \N__26763\
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__26763\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__6059\ : CascadeMux
    port map (
            O => \N__26760\,
            I => \N__26757\
        );

    \I__6058\ : InMux
    port map (
            O => \N__26757\,
            I => \N__26754\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__6056\ : Odrv12
    port map (
            O => \N__26751\,
            I => \M_this_state_d22\
        );

    \I__6055\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26745\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__26745\,
            I => \N__26742\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__26742\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11\
        );

    \I__6052\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26736\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__26736\,
            I => \N__26732\
        );

    \I__6050\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26728\
        );

    \I__6049\ : Span4Mux_v
    port map (
            O => \N__26732\,
            I => \N__26722\
        );

    \I__6048\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26719\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__26728\,
            I => \N__26716\
        );

    \I__6046\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26709\
        );

    \I__6045\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26709\
        );

    \I__6044\ : InMux
    port map (
            O => \N__26725\,
            I => \N__26709\
        );

    \I__6043\ : Sp12to4
    port map (
            O => \N__26722\,
            I => \N__26703\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26703\
        );

    \I__6041\ : Span4Mux_h
    port map (
            O => \N__26716\,
            I => \N__26698\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__26709\,
            I => \N__26698\
        );

    \I__6039\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26695\
        );

    \I__6038\ : Span12Mux_h
    port map (
            O => \N__26703\,
            I => \N__26690\
        );

    \I__6037\ : Sp12to4
    port map (
            O => \N__26698\,
            I => \N__26690\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__26695\,
            I => \N__26687\
        );

    \I__6035\ : Odrv12
    port map (
            O => \N__26690\,
            I => port_address_in_0
        );

    \I__6034\ : Odrv12
    port map (
            O => \N__26687\,
            I => port_address_in_0
        );

    \I__6033\ : CascadeMux
    port map (
            O => \N__26682\,
            I => \N__26678\
        );

    \I__6032\ : InMux
    port map (
            O => \N__26681\,
            I => \N__26673\
        );

    \I__6031\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26673\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__26673\,
            I => \this_vga_signals.M_this_state_d21Z0Z_6\
        );

    \I__6029\ : CascadeMux
    port map (
            O => \N__26670\,
            I => \N__26667\
        );

    \I__6028\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26663\
        );

    \I__6027\ : CascadeMux
    port map (
            O => \N__26666\,
            I => \N__26660\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__26663\,
            I => \N__26657\
        );

    \I__6025\ : InMux
    port map (
            O => \N__26660\,
            I => \N__26654\
        );

    \I__6024\ : Span4Mux_v
    port map (
            O => \N__26657\,
            I => \N__26651\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__26654\,
            I => \N__26648\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__26651\,
            I => \N__26643\
        );

    \I__6021\ : Span4Mux_v
    port map (
            O => \N__26648\,
            I => \N__26643\
        );

    \I__6020\ : Odrv4
    port map (
            O => \N__26643\,
            I => \this_vga_signals.M_this_state_dZ0Z24\
        );

    \I__6019\ : InMux
    port map (
            O => \N__26640\,
            I => \N__26637\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__26637\,
            I => \N__26634\
        );

    \I__6017\ : Odrv4
    port map (
            O => \N__26634\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8\
        );

    \I__6016\ : CascadeMux
    port map (
            O => \N__26631\,
            I => \N__26628\
        );

    \I__6015\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26625\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__26625\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_8\
        );

    \I__6013\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26619\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__26619\,
            I => \N__26616\
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__26616\,
            I => \un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0\
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__26613\,
            I => \N__26610\
        );

    \I__6009\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26605\
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__26609\,
            I => \N__26602\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__26608\,
            I => \N__26599\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__26605\,
            I => \N__26594\
        );

    \I__6005\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26591\
        );

    \I__6004\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26588\
        );

    \I__6003\ : CascadeMux
    port map (
            O => \N__26598\,
            I => \N__26585\
        );

    \I__6002\ : CascadeMux
    port map (
            O => \N__26597\,
            I => \N__26581\
        );

    \I__6001\ : Span4Mux_h
    port map (
            O => \N__26594\,
            I => \N__26573\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26573\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__26588\,
            I => \N__26570\
        );

    \I__5998\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26567\
        );

    \I__5997\ : CascadeMux
    port map (
            O => \N__26584\,
            I => \N__26564\
        );

    \I__5996\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26558\
        );

    \I__5995\ : CascadeMux
    port map (
            O => \N__26580\,
            I => \N__26555\
        );

    \I__5994\ : CascadeMux
    port map (
            O => \N__26579\,
            I => \N__26552\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__26578\,
            I => \N__26549\
        );

    \I__5992\ : Span4Mux_v
    port map (
            O => \N__26573\,
            I => \N__26542\
        );

    \I__5991\ : Span4Mux_h
    port map (
            O => \N__26570\,
            I => \N__26542\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__26567\,
            I => \N__26542\
        );

    \I__5989\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26539\
        );

    \I__5988\ : CascadeMux
    port map (
            O => \N__26563\,
            I => \N__26536\
        );

    \I__5987\ : CascadeMux
    port map (
            O => \N__26562\,
            I => \N__26532\
        );

    \I__5986\ : CascadeMux
    port map (
            O => \N__26561\,
            I => \N__26529\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__26558\,
            I => \N__26524\
        );

    \I__5984\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26521\
        );

    \I__5983\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26518\
        );

    \I__5982\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26515\
        );

    \I__5981\ : Span4Mux_v
    port map (
            O => \N__26542\,
            I => \N__26510\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__26539\,
            I => \N__26510\
        );

    \I__5979\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26507\
        );

    \I__5978\ : CascadeMux
    port map (
            O => \N__26535\,
            I => \N__26504\
        );

    \I__5977\ : InMux
    port map (
            O => \N__26532\,
            I => \N__26501\
        );

    \I__5976\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26498\
        );

    \I__5975\ : CascadeMux
    port map (
            O => \N__26528\,
            I => \N__26495\
        );

    \I__5974\ : CascadeMux
    port map (
            O => \N__26527\,
            I => \N__26492\
        );

    \I__5973\ : Span4Mux_v
    port map (
            O => \N__26524\,
            I => \N__26486\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__26521\,
            I => \N__26486\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__26518\,
            I => \N__26481\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__26515\,
            I => \N__26481\
        );

    \I__5969\ : Span4Mux_h
    port map (
            O => \N__26510\,
            I => \N__26476\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__26507\,
            I => \N__26476\
        );

    \I__5967\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26473\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__26501\,
            I => \N__26470\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__26498\,
            I => \N__26467\
        );

    \I__5964\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26464\
        );

    \I__5963\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26461\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__26491\,
            I => \N__26458\
        );

    \I__5961\ : Span4Mux_v
    port map (
            O => \N__26486\,
            I => \N__26453\
        );

    \I__5960\ : Span4Mux_v
    port map (
            O => \N__26481\,
            I => \N__26453\
        );

    \I__5959\ : Span4Mux_v
    port map (
            O => \N__26476\,
            I => \N__26448\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__26473\,
            I => \N__26448\
        );

    \I__5957\ : Span4Mux_v
    port map (
            O => \N__26470\,
            I => \N__26441\
        );

    \I__5956\ : Span4Mux_h
    port map (
            O => \N__26467\,
            I => \N__26441\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__26464\,
            I => \N__26441\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__26461\,
            I => \N__26438\
        );

    \I__5953\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26435\
        );

    \I__5952\ : Sp12to4
    port map (
            O => \N__26453\,
            I => \N__26430\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__26448\,
            I => \N__26427\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__26441\,
            I => \N__26420\
        );

    \I__5949\ : Span4Mux_v
    port map (
            O => \N__26438\,
            I => \N__26420\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__26435\,
            I => \N__26420\
        );

    \I__5947\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26416\
        );

    \I__5946\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26413\
        );

    \I__5945\ : Span12Mux_h
    port map (
            O => \N__26430\,
            I => \N__26410\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__26427\,
            I => \N__26405\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__26420\,
            I => \N__26405\
        );

    \I__5942\ : InMux
    port map (
            O => \N__26419\,
            I => \N__26402\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__26416\,
            I => \N__26399\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__26413\,
            I => \N__26396\
        );

    \I__5939\ : Odrv12
    port map (
            O => \N__26410\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__5938\ : Odrv4
    port map (
            O => \N__26405\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__26402\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__26399\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__5935\ : Odrv4
    port map (
            O => \N__26396\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__26385\,
            I => \N__26380\
        );

    \I__5933\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26370\
        );

    \I__5932\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26365\
        );

    \I__5931\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26365\
        );

    \I__5930\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26362\
        );

    \I__5929\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26359\
        );

    \I__5928\ : InMux
    port map (
            O => \N__26377\,
            I => \N__26353\
        );

    \I__5927\ : InMux
    port map (
            O => \N__26376\,
            I => \N__26349\
        );

    \I__5926\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26346\
        );

    \I__5925\ : InMux
    port map (
            O => \N__26374\,
            I => \N__26343\
        );

    \I__5924\ : InMux
    port map (
            O => \N__26373\,
            I => \N__26340\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__26370\,
            I => \N__26335\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__26365\,
            I => \N__26335\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__26362\,
            I => \N__26330\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__26359\,
            I => \N__26330\
        );

    \I__5919\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26325\
        );

    \I__5918\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26325\
        );

    \I__5917\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26322\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__26353\,
            I => \N__26319\
        );

    \I__5915\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26315\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__26349\,
            I => \N__26310\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26310\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__26343\,
            I => \N__26307\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__26340\,
            I => \N__26298\
        );

    \I__5910\ : Span4Mux_v
    port map (
            O => \N__26335\,
            I => \N__26298\
        );

    \I__5909\ : Span4Mux_h
    port map (
            O => \N__26330\,
            I => \N__26298\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__26325\,
            I => \N__26298\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__26322\,
            I => \N__26293\
        );

    \I__5906\ : Span4Mux_h
    port map (
            O => \N__26319\,
            I => \N__26293\
        );

    \I__5905\ : InMux
    port map (
            O => \N__26318\,
            I => \N__26287\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__26315\,
            I => \N__26284\
        );

    \I__5903\ : Span4Mux_h
    port map (
            O => \N__26310\,
            I => \N__26281\
        );

    \I__5902\ : Span4Mux_h
    port map (
            O => \N__26307\,
            I => \N__26276\
        );

    \I__5901\ : Span4Mux_h
    port map (
            O => \N__26298\,
            I => \N__26276\
        );

    \I__5900\ : Span4Mux_h
    port map (
            O => \N__26293\,
            I => \N__26273\
        );

    \I__5899\ : InMux
    port map (
            O => \N__26292\,
            I => \N__26268\
        );

    \I__5898\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26268\
        );

    \I__5897\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26265\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__26287\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5895\ : Odrv12
    port map (
            O => \N__26284\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5894\ : Odrv4
    port map (
            O => \N__26281\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__26276\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__26273\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__26268\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__26265\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5889\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26247\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__26247\,
            I => \N__26244\
        );

    \I__5887\ : Span4Mux_v
    port map (
            O => \N__26244\,
            I => \N__26241\
        );

    \I__5886\ : Odrv4
    port map (
            O => \N__26241\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1\
        );

    \I__5885\ : CascadeMux
    port map (
            O => \N__26238\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_1_cascade_\
        );

    \I__5884\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26232\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__26232\,
            I => \N__26229\
        );

    \I__5882\ : Span4Mux_h
    port map (
            O => \N__26229\,
            I => \N__26226\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__26226\,
            I => \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__26223\,
            I => \N__26219\
        );

    \I__5879\ : CascadeMux
    port map (
            O => \N__26222\,
            I => \N__26216\
        );

    \I__5878\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26211\
        );

    \I__5877\ : InMux
    port map (
            O => \N__26216\,
            I => \N__26208\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__26215\,
            I => \N__26205\
        );

    \I__5875\ : CascadeMux
    port map (
            O => \N__26214\,
            I => \N__26202\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__26211\,
            I => \N__26191\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__26208\,
            I => \N__26191\
        );

    \I__5872\ : InMux
    port map (
            O => \N__26205\,
            I => \N__26188\
        );

    \I__5871\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26185\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__26201\,
            I => \N__26182\
        );

    \I__5869\ : CascadeMux
    port map (
            O => \N__26200\,
            I => \N__26179\
        );

    \I__5868\ : CascadeMux
    port map (
            O => \N__26199\,
            I => \N__26173\
        );

    \I__5867\ : CascadeMux
    port map (
            O => \N__26198\,
            I => \N__26170\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__26197\,
            I => \N__26167\
        );

    \I__5865\ : CascadeMux
    port map (
            O => \N__26196\,
            I => \N__26164\
        );

    \I__5864\ : Span4Mux_v
    port map (
            O => \N__26191\,
            I => \N__26157\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__26188\,
            I => \N__26157\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__26185\,
            I => \N__26157\
        );

    \I__5861\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26154\
        );

    \I__5860\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26151\
        );

    \I__5859\ : CascadeMux
    port map (
            O => \N__26178\,
            I => \N__26148\
        );

    \I__5858\ : CascadeMux
    port map (
            O => \N__26177\,
            I => \N__26144\
        );

    \I__5857\ : CascadeMux
    port map (
            O => \N__26176\,
            I => \N__26141\
        );

    \I__5856\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26135\
        );

    \I__5855\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26132\
        );

    \I__5854\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26129\
        );

    \I__5853\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26126\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__26157\,
            I => \N__26119\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__26154\,
            I => \N__26119\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__26151\,
            I => \N__26119\
        );

    \I__5849\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26116\
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__26147\,
            I => \N__26113\
        );

    \I__5847\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26110\
        );

    \I__5846\ : InMux
    port map (
            O => \N__26141\,
            I => \N__26107\
        );

    \I__5845\ : CascadeMux
    port map (
            O => \N__26140\,
            I => \N__26104\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__26139\,
            I => \N__26101\
        );

    \I__5843\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26098\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__26135\,
            I => \N__26090\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__26132\,
            I => \N__26090\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__26129\,
            I => \N__26090\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__26126\,
            I => \N__26087\
        );

    \I__5838\ : Span4Mux_v
    port map (
            O => \N__26119\,
            I => \N__26082\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__26116\,
            I => \N__26082\
        );

    \I__5836\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26079\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__26110\,
            I => \N__26074\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__26074\
        );

    \I__5833\ : InMux
    port map (
            O => \N__26104\,
            I => \N__26071\
        );

    \I__5832\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26068\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__26098\,
            I => \N__26065\
        );

    \I__5830\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26062\
        );

    \I__5829\ : Span12Mux_v
    port map (
            O => \N__26090\,
            I => \N__26057\
        );

    \I__5828\ : Span12Mux_s9_v
    port map (
            O => \N__26087\,
            I => \N__26057\
        );

    \I__5827\ : Span4Mux_v
    port map (
            O => \N__26082\,
            I => \N__26052\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__26079\,
            I => \N__26052\
        );

    \I__5825\ : Span4Mux_v
    port map (
            O => \N__26074\,
            I => \N__26045\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__26071\,
            I => \N__26045\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__26068\,
            I => \N__26045\
        );

    \I__5822\ : Span4Mux_v
    port map (
            O => \N__26065\,
            I => \N__26039\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__26062\,
            I => \N__26039\
        );

    \I__5820\ : Span12Mux_h
    port map (
            O => \N__26057\,
            I => \N__26036\
        );

    \I__5819\ : Span4Mux_v
    port map (
            O => \N__26052\,
            I => \N__26031\
        );

    \I__5818\ : Span4Mux_v
    port map (
            O => \N__26045\,
            I => \N__26031\
        );

    \I__5817\ : InMux
    port map (
            O => \N__26044\,
            I => \N__26028\
        );

    \I__5816\ : Span4Mux_h
    port map (
            O => \N__26039\,
            I => \N__26025\
        );

    \I__5815\ : Odrv12
    port map (
            O => \N__26036\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5814\ : Odrv4
    port map (
            O => \N__26031\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__26028\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__26025\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5811\ : InMux
    port map (
            O => \N__26016\,
            I => \bfn_21_19_0_\
        );

    \I__5810\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26007\
        );

    \I__5809\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26000\
        );

    \I__5808\ : InMux
    port map (
            O => \N__26011\,
            I => \N__26000\
        );

    \I__5807\ : InMux
    port map (
            O => \N__26010\,
            I => \N__26000\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__26007\,
            I => \this_ppu.vscroll8\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__26000\,
            I => \this_ppu.vscroll8\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__25995\,
            I => \N__25991\
        );

    \I__5803\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25988\
        );

    \I__5802\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25985\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__25988\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__25985\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__5799\ : InMux
    port map (
            O => \N__25980\,
            I => \N__25977\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__25977\,
            I => \N__25974\
        );

    \I__5797\ : Span4Mux_v
    port map (
            O => \N__25974\,
            I => \N__25971\
        );

    \I__5796\ : Span4Mux_h
    port map (
            O => \N__25971\,
            I => \N__25968\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__25968\,
            I => \N_48_0\
        );

    \I__5794\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25962\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__25962\,
            I => \N__25959\
        );

    \I__5792\ : Span4Mux_h
    port map (
            O => \N__25959\,
            I => \N__25956\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__25956\,
            I => \M_this_oam_ram_write_data_28\
        );

    \I__5790\ : CascadeMux
    port map (
            O => \N__25953\,
            I => \N__25948\
        );

    \I__5789\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25944\
        );

    \I__5788\ : InMux
    port map (
            O => \N__25951\,
            I => \N__25937\
        );

    \I__5787\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25937\
        );

    \I__5786\ : InMux
    port map (
            O => \N__25947\,
            I => \N__25937\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__25944\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__25937\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__5783\ : CascadeMux
    port map (
            O => \N__25932\,
            I => \N__25927\
        );

    \I__5782\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25922\
        );

    \I__5781\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25918\
        );

    \I__5780\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25915\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__25926\,
            I => \N__25912\
        );

    \I__5778\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25907\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__25922\,
            I => \N__25904\
        );

    \I__5776\ : InMux
    port map (
            O => \N__25921\,
            I => \N__25901\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__25918\,
            I => \N__25896\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__25915\,
            I => \N__25896\
        );

    \I__5773\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25891\
        );

    \I__5772\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25891\
        );

    \I__5771\ : InMux
    port map (
            O => \N__25910\,
            I => \N__25888\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__25907\,
            I => \N__25885\
        );

    \I__5769\ : Span4Mux_v
    port map (
            O => \N__25904\,
            I => \N__25880\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__25901\,
            I => \N__25880\
        );

    \I__5767\ : Span4Mux_v
    port map (
            O => \N__25896\,
            I => \N__25877\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__25891\,
            I => \N__25874\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__25888\,
            I => \N__25871\
        );

    \I__5764\ : Span4Mux_h
    port map (
            O => \N__25885\,
            I => \N__25866\
        );

    \I__5763\ : Span4Mux_h
    port map (
            O => \N__25880\,
            I => \N__25866\
        );

    \I__5762\ : Odrv4
    port map (
            O => \N__25877\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__25874\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__5760\ : Odrv12
    port map (
            O => \N__25871\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__5759\ : Odrv4
    port map (
            O => \N__25866\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__5758\ : InMux
    port map (
            O => \N__25857\,
            I => \N__25853\
        );

    \I__5757\ : InMux
    port map (
            O => \N__25856\,
            I => \N__25850\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__25853\,
            I => \N__25847\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__25850\,
            I => \N__25843\
        );

    \I__5754\ : Span12Mux_h
    port map (
            O => \N__25847\,
            I => \N__25840\
        );

    \I__5753\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25837\
        );

    \I__5752\ : Odrv12
    port map (
            O => \N__25843\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_7\
        );

    \I__5751\ : Odrv12
    port map (
            O => \N__25840\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_7\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__25837\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_7\
        );

    \I__5749\ : InMux
    port map (
            O => \N__25830\,
            I => \N__25827\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__25827\,
            I => \this_ppu.N_148\
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__25824\,
            I => \N__25821\
        );

    \I__5746\ : InMux
    port map (
            O => \N__25821\,
            I => \N__25818\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__25818\,
            I => \N__25815\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__25815\,
            I => \M_this_data_tmp_qZ0Z_20\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__5742\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25804\
        );

    \I__5741\ : CascadeMux
    port map (
            O => \N__25808\,
            I => \N__25801\
        );

    \I__5740\ : CascadeMux
    port map (
            O => \N__25807\,
            I => \N__25795\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__25804\,
            I => \N__25791\
        );

    \I__5738\ : InMux
    port map (
            O => \N__25801\,
            I => \N__25788\
        );

    \I__5737\ : CascadeMux
    port map (
            O => \N__25800\,
            I => \N__25785\
        );

    \I__5736\ : CascadeMux
    port map (
            O => \N__25799\,
            I => \N__25781\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__25798\,
            I => \N__25777\
        );

    \I__5734\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25772\
        );

    \I__5733\ : CascadeMux
    port map (
            O => \N__25794\,
            I => \N__25769\
        );

    \I__5732\ : Span4Mux_s2_v
    port map (
            O => \N__25791\,
            I => \N__25764\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__25788\,
            I => \N__25764\
        );

    \I__5730\ : InMux
    port map (
            O => \N__25785\,
            I => \N__25761\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__25784\,
            I => \N__25758\
        );

    \I__5728\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25754\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__25780\,
            I => \N__25751\
        );

    \I__5726\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25748\
        );

    \I__5725\ : CascadeMux
    port map (
            O => \N__25776\,
            I => \N__25745\
        );

    \I__5724\ : CascadeMux
    port map (
            O => \N__25775\,
            I => \N__25742\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__25772\,
            I => \N__25737\
        );

    \I__5722\ : InMux
    port map (
            O => \N__25769\,
            I => \N__25734\
        );

    \I__5721\ : Span4Mux_v
    port map (
            O => \N__25764\,
            I => \N__25729\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__25761\,
            I => \N__25729\
        );

    \I__5719\ : InMux
    port map (
            O => \N__25758\,
            I => \N__25726\
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__25757\,
            I => \N__25723\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__25754\,
            I => \N__25719\
        );

    \I__5716\ : InMux
    port map (
            O => \N__25751\,
            I => \N__25716\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__25748\,
            I => \N__25712\
        );

    \I__5714\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25709\
        );

    \I__5713\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25706\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__25741\,
            I => \N__25703\
        );

    \I__5711\ : CascadeMux
    port map (
            O => \N__25740\,
            I => \N__25700\
        );

    \I__5710\ : Span4Mux_h
    port map (
            O => \N__25737\,
            I => \N__25697\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__25734\,
            I => \N__25694\
        );

    \I__5708\ : Span4Mux_h
    port map (
            O => \N__25729\,
            I => \N__25689\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__25726\,
            I => \N__25689\
        );

    \I__5706\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25686\
        );

    \I__5705\ : CascadeMux
    port map (
            O => \N__25722\,
            I => \N__25683\
        );

    \I__5704\ : Span4Mux_v
    port map (
            O => \N__25719\,
            I => \N__25678\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__25716\,
            I => \N__25678\
        );

    \I__5702\ : CascadeMux
    port map (
            O => \N__25715\,
            I => \N__25675\
        );

    \I__5701\ : Span4Mux_v
    port map (
            O => \N__25712\,
            I => \N__25670\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__25709\,
            I => \N__25670\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__25706\,
            I => \N__25667\
        );

    \I__5698\ : InMux
    port map (
            O => \N__25703\,
            I => \N__25664\
        );

    \I__5697\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25661\
        );

    \I__5696\ : Span4Mux_h
    port map (
            O => \N__25697\,
            I => \N__25658\
        );

    \I__5695\ : Span4Mux_h
    port map (
            O => \N__25694\,
            I => \N__25655\
        );

    \I__5694\ : Span4Mux_v
    port map (
            O => \N__25689\,
            I => \N__25650\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25650\
        );

    \I__5692\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25647\
        );

    \I__5691\ : Span4Mux_h
    port map (
            O => \N__25678\,
            I => \N__25644\
        );

    \I__5690\ : InMux
    port map (
            O => \N__25675\,
            I => \N__25641\
        );

    \I__5689\ : Span4Mux_v
    port map (
            O => \N__25670\,
            I => \N__25632\
        );

    \I__5688\ : Span4Mux_v
    port map (
            O => \N__25667\,
            I => \N__25632\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__25664\,
            I => \N__25632\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__25661\,
            I => \N__25632\
        );

    \I__5685\ : Span4Mux_v
    port map (
            O => \N__25658\,
            I => \N__25627\
        );

    \I__5684\ : Span4Mux_h
    port map (
            O => \N__25655\,
            I => \N__25627\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__25650\,
            I => \N__25622\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__25647\,
            I => \N__25622\
        );

    \I__5681\ : Span4Mux_v
    port map (
            O => \N__25644\,
            I => \N__25619\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__25641\,
            I => \N__25616\
        );

    \I__5679\ : Span4Mux_v
    port map (
            O => \N__25632\,
            I => \N__25613\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__25627\,
            I => \N__25608\
        );

    \I__5677\ : Span4Mux_h
    port map (
            O => \N__25622\,
            I => \N__25608\
        );

    \I__5676\ : Sp12to4
    port map (
            O => \N__25619\,
            I => \N__25605\
        );

    \I__5675\ : Span12Mux_s11_h
    port map (
            O => \N__25616\,
            I => \N__25602\
        );

    \I__5674\ : Span4Mux_h
    port map (
            O => \N__25613\,
            I => \N__25597\
        );

    \I__5673\ : Span4Mux_h
    port map (
            O => \N__25608\,
            I => \N__25597\
        );

    \I__5672\ : Odrv12
    port map (
            O => \N__25605\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__5671\ : Odrv12
    port map (
            O => \N__25602\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__5670\ : Odrv4
    port map (
            O => \N__25597\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__5669\ : CascadeMux
    port map (
            O => \N__25590\,
            I => \N__25587\
        );

    \I__5668\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25584\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__5666\ : Span12Mux_v
    port map (
            O => \N__25581\,
            I => \N__25577\
        );

    \I__5665\ : CascadeMux
    port map (
            O => \N__25580\,
            I => \N__25574\
        );

    \I__5664\ : Span12Mux_h
    port map (
            O => \N__25577\,
            I => \N__25564\
        );

    \I__5663\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25553\
        );

    \I__5662\ : InMux
    port map (
            O => \N__25573\,
            I => \N__25553\
        );

    \I__5661\ : InMux
    port map (
            O => \N__25572\,
            I => \N__25553\
        );

    \I__5660\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25553\
        );

    \I__5659\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25553\
        );

    \I__5658\ : InMux
    port map (
            O => \N__25569\,
            I => \N__25550\
        );

    \I__5657\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25547\
        );

    \I__5656\ : InMux
    port map (
            O => \N__25567\,
            I => \N__25544\
        );

    \I__5655\ : Odrv12
    port map (
            O => \N__25564\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__25553\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__25550\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__25547\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__25544\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__25533\,
            I => \N__25530\
        );

    \I__5649\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25527\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__25527\,
            I => \N__25524\
        );

    \I__5647\ : Span4Mux_h
    port map (
            O => \N__25524\,
            I => \N__25521\
        );

    \I__5646\ : Span4Mux_h
    port map (
            O => \N__25521\,
            I => \N__25514\
        );

    \I__5645\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25509\
        );

    \I__5644\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25509\
        );

    \I__5643\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25506\
        );

    \I__5642\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25503\
        );

    \I__5641\ : Span4Mux_h
    port map (
            O => \N__25514\,
            I => \N__25498\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__25509\,
            I => \N__25491\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__25506\,
            I => \N__25491\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__25503\,
            I => \N__25491\
        );

    \I__5637\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25488\
        );

    \I__5636\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25485\
        );

    \I__5635\ : Odrv4
    port map (
            O => \N__25498\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__5634\ : Odrv4
    port map (
            O => \N__25491\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__25488\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__25485\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__5631\ : CascadeMux
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__5630\ : InMux
    port map (
            O => \N__25473\,
            I => \N__25470\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__25470\,
            I => \N__25465\
        );

    \I__5628\ : InMux
    port map (
            O => \N__25469\,
            I => \N__25455\
        );

    \I__5627\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25455\
        );

    \I__5626\ : Span12Mux_h
    port map (
            O => \N__25465\,
            I => \N__25452\
        );

    \I__5625\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25449\
        );

    \I__5624\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25444\
        );

    \I__5623\ : InMux
    port map (
            O => \N__25462\,
            I => \N__25444\
        );

    \I__5622\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25441\
        );

    \I__5621\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25438\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__25455\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__5619\ : Odrv12
    port map (
            O => \N__25452\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__25449\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__25444\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__25441\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__25438\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__25425\,
            I => \N__25422\
        );

    \I__5613\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25419\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__25419\,
            I => \M_this_oam_ram_read_data_i_11\
        );

    \I__5611\ : CascadeMux
    port map (
            O => \N__25416\,
            I => \N__25413\
        );

    \I__5610\ : CascadeBuf
    port map (
            O => \N__25413\,
            I => \N__25409\
        );

    \I__5609\ : CascadeMux
    port map (
            O => \N__25412\,
            I => \N__25406\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__25409\,
            I => \N__25403\
        );

    \I__5607\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25400\
        );

    \I__5606\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25397\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__25400\,
            I => \N__25394\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__25397\,
            I => \N__25391\
        );

    \I__5603\ : Span4Mux_h
    port map (
            O => \N__25394\,
            I => \N__25388\
        );

    \I__5602\ : Span4Mux_h
    port map (
            O => \N__25391\,
            I => \N__25385\
        );

    \I__5601\ : Span4Mux_h
    port map (
            O => \N__25388\,
            I => \N__25378\
        );

    \I__5600\ : Sp12to4
    port map (
            O => \N__25385\,
            I => \N__25375\
        );

    \I__5599\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25370\
        );

    \I__5598\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25370\
        );

    \I__5597\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25367\
        );

    \I__5596\ : InMux
    port map (
            O => \N__25381\,
            I => \N__25364\
        );

    \I__5595\ : Span4Mux_h
    port map (
            O => \N__25378\,
            I => \N__25361\
        );

    \I__5594\ : Span12Mux_v
    port map (
            O => \N__25375\,
            I => \N__25358\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__25370\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__25367\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__25364\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__25361\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__5589\ : Odrv12
    port map (
            O => \N__25358\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__5588\ : CascadeMux
    port map (
            O => \N__25347\,
            I => \N__25344\
        );

    \I__5587\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25341\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__25341\,
            I => \N__25338\
        );

    \I__5585\ : Odrv4
    port map (
            O => \N__25338\,
            I => \this_ppu.un1_M_haddress_q_2_4\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__25335\,
            I => \N__25331\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__25334\,
            I => \N__25328\
        );

    \I__5582\ : CascadeBuf
    port map (
            O => \N__25331\,
            I => \N__25325\
        );

    \I__5581\ : InMux
    port map (
            O => \N__25328\,
            I => \N__25322\
        );

    \I__5580\ : CascadeMux
    port map (
            O => \N__25325\,
            I => \N__25319\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25316\
        );

    \I__5578\ : InMux
    port map (
            O => \N__25319\,
            I => \N__25313\
        );

    \I__5577\ : Sp12to4
    port map (
            O => \N__25316\,
            I => \N__25309\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__25313\,
            I => \N__25306\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__25312\,
            I => \N__25303\
        );

    \I__5574\ : Span12Mux_v
    port map (
            O => \N__25309\,
            I => \N__25298\
        );

    \I__5573\ : Span12Mux_s8_v
    port map (
            O => \N__25306\,
            I => \N__25295\
        );

    \I__5572\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25292\
        );

    \I__5571\ : InMux
    port map (
            O => \N__25302\,
            I => \N__25289\
        );

    \I__5570\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25286\
        );

    \I__5569\ : Span12Mux_h
    port map (
            O => \N__25298\,
            I => \N__25281\
        );

    \I__5568\ : Span12Mux_h
    port map (
            O => \N__25295\,
            I => \N__25281\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__25292\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__25289\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__25286\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__5564\ : Odrv12
    port map (
            O => \N__25281\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__5562\ : CascadeBuf
    port map (
            O => \N__25269\,
            I => \N__25265\
        );

    \I__5561\ : CascadeMux
    port map (
            O => \N__25268\,
            I => \N__25262\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__25265\,
            I => \N__25259\
        );

    \I__5559\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25253\
        );

    \I__5558\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25250\
        );

    \I__5557\ : CascadeMux
    port map (
            O => \N__25258\,
            I => \N__25247\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__25257\,
            I => \N__25244\
        );

    \I__5555\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25240\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__25253\,
            I => \N__25237\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__25250\,
            I => \N__25234\
        );

    \I__5552\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25227\
        );

    \I__5551\ : InMux
    port map (
            O => \N__25244\,
            I => \N__25227\
        );

    \I__5550\ : InMux
    port map (
            O => \N__25243\,
            I => \N__25227\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__25240\,
            I => \N__25222\
        );

    \I__5548\ : Span12Mux_h
    port map (
            O => \N__25237\,
            I => \N__25222\
        );

    \I__5547\ : Span12Mux_h
    port map (
            O => \N__25234\,
            I => \N__25219\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__25227\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__5545\ : Odrv12
    port map (
            O => \N__25222\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__5544\ : Odrv12
    port map (
            O => \N__25219\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__25212\,
            I => \N__25209\
        );

    \I__5542\ : CascadeBuf
    port map (
            O => \N__25209\,
            I => \N__25206\
        );

    \I__5541\ : CascadeMux
    port map (
            O => \N__25206\,
            I => \N__25203\
        );

    \I__5540\ : InMux
    port map (
            O => \N__25203\,
            I => \N__25199\
        );

    \I__5539\ : CascadeMux
    port map (
            O => \N__25202\,
            I => \N__25196\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__25199\,
            I => \N__25193\
        );

    \I__5537\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25189\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__25193\,
            I => \N__25186\
        );

    \I__5535\ : InMux
    port map (
            O => \N__25192\,
            I => \N__25181\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__25189\,
            I => \N__25178\
        );

    \I__5533\ : Sp12to4
    port map (
            O => \N__25186\,
            I => \N__25175\
        );

    \I__5532\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25170\
        );

    \I__5531\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25170\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__25181\,
            I => \N__25165\
        );

    \I__5529\ : Span12Mux_s11_h
    port map (
            O => \N__25178\,
            I => \N__25165\
        );

    \I__5528\ : Span12Mux_h
    port map (
            O => \N__25175\,
            I => \N__25162\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__25170\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__5526\ : Odrv12
    port map (
            O => \N__25165\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__5525\ : Odrv12
    port map (
            O => \N__25162\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__5524\ : CascadeMux
    port map (
            O => \N__25155\,
            I => \N__25152\
        );

    \I__5523\ : CascadeBuf
    port map (
            O => \N__25152\,
            I => \N__25149\
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__25149\,
            I => \N__25146\
        );

    \I__5521\ : InMux
    port map (
            O => \N__25146\,
            I => \N__25143\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__25143\,
            I => \N__25140\
        );

    \I__5519\ : Span4Mux_v
    port map (
            O => \N__25140\,
            I => \N__25136\
        );

    \I__5518\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25132\
        );

    \I__5517\ : Sp12to4
    port map (
            O => \N__25136\,
            I => \N__25129\
        );

    \I__5516\ : InMux
    port map (
            O => \N__25135\,
            I => \N__25126\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__25132\,
            I => \N__25123\
        );

    \I__5514\ : Span12Mux_h
    port map (
            O => \N__25129\,
            I => \N__25120\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__25126\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__25123\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__5511\ : Odrv12
    port map (
            O => \N__25120\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__25113\,
            I => \N__25110\
        );

    \I__5509\ : InMux
    port map (
            O => \N__25110\,
            I => \N__25107\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__25107\,
            I => \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\
        );

    \I__5507\ : InMux
    port map (
            O => \N__25104\,
            I => \this_ppu.un2_hscroll_cry_0\
        );

    \I__5506\ : InMux
    port map (
            O => \N__25101\,
            I => \this_ppu.un2_hscroll_cry_1\
        );

    \I__5505\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25095\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__25095\,
            I => \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0\
        );

    \I__5503\ : CEMux
    port map (
            O => \N__25092\,
            I => \N__25089\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__25089\,
            I => \N__25085\
        );

    \I__5501\ : CEMux
    port map (
            O => \N__25088\,
            I => \N__25082\
        );

    \I__5500\ : Span4Mux_h
    port map (
            O => \N__25085\,
            I => \N__25077\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__25082\,
            I => \N__25077\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__25077\,
            I => \N__25074\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__25074\,
            I => \N__25071\
        );

    \I__5496\ : Odrv4
    port map (
            O => \N__25071\,
            I => \this_sprites_ram.mem_WE_12\
        );

    \I__5495\ : InMux
    port map (
            O => \N__25068\,
            I => \N__25065\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__25065\,
            I => \N__25062\
        );

    \I__5493\ : Span4Mux_h
    port map (
            O => \N__25062\,
            I => \N__25059\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__25059\,
            I => \N__25056\
        );

    \I__5491\ : Span4Mux_v
    port map (
            O => \N__25056\,
            I => \N__25053\
        );

    \I__5490\ : Odrv4
    port map (
            O => \N__25053\,
            I => \this_sprites_ram.mem_out_bus6_2\
        );

    \I__5489\ : InMux
    port map (
            O => \N__25050\,
            I => \N__25047\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__25047\,
            I => \N__25044\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__25044\,
            I => \N__25041\
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__25041\,
            I => \this_sprites_ram.mem_out_bus2_2\
        );

    \I__5485\ : InMux
    port map (
            O => \N__25038\,
            I => \N__25035\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__25035\,
            I => \N__25032\
        );

    \I__5483\ : Odrv12
    port map (
            O => \N__25032\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\
        );

    \I__5482\ : CascadeMux
    port map (
            O => \N__25029\,
            I => \N__25026\
        );

    \I__5481\ : InMux
    port map (
            O => \N__25026\,
            I => \N__25023\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__25023\,
            I => \M_this_oam_ram_read_data_i_9\
        );

    \I__5479\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25017\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__25017\,
            I => \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0\
        );

    \I__5477\ : CascadeMux
    port map (
            O => \N__25014\,
            I => \N__25009\
        );

    \I__5476\ : CascadeMux
    port map (
            O => \N__25013\,
            I => \N__25006\
        );

    \I__5475\ : InMux
    port map (
            O => \N__25012\,
            I => \N__24999\
        );

    \I__5474\ : InMux
    port map (
            O => \N__25009\,
            I => \N__24990\
        );

    \I__5473\ : InMux
    port map (
            O => \N__25006\,
            I => \N__24990\
        );

    \I__5472\ : InMux
    port map (
            O => \N__25005\,
            I => \N__24987\
        );

    \I__5471\ : InMux
    port map (
            O => \N__25004\,
            I => \N__24979\
        );

    \I__5470\ : InMux
    port map (
            O => \N__25003\,
            I => \N__24979\
        );

    \I__5469\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24976\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__24999\,
            I => \N__24973\
        );

    \I__5467\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24966\
        );

    \I__5466\ : InMux
    port map (
            O => \N__24997\,
            I => \N__24966\
        );

    \I__5465\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24966\
        );

    \I__5464\ : CascadeMux
    port map (
            O => \N__24995\,
            I => \N__24962\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__24990\,
            I => \N__24957\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__24987\,
            I => \N__24954\
        );

    \I__5461\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24949\
        );

    \I__5460\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24949\
        );

    \I__5459\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24946\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__24979\,
            I => \N__24937\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__24976\,
            I => \N__24937\
        );

    \I__5456\ : Span4Mux_v
    port map (
            O => \N__24973\,
            I => \N__24937\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__24966\,
            I => \N__24937\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__24965\,
            I => \N__24934\
        );

    \I__5453\ : InMux
    port map (
            O => \N__24962\,
            I => \N__24930\
        );

    \I__5452\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24927\
        );

    \I__5451\ : InMux
    port map (
            O => \N__24960\,
            I => \N__24924\
        );

    \I__5450\ : Span4Mux_h
    port map (
            O => \N__24957\,
            I => \N__24919\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__24954\,
            I => \N__24919\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__24949\,
            I => \N__24916\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__24946\,
            I => \N__24911\
        );

    \I__5446\ : Span4Mux_h
    port map (
            O => \N__24937\,
            I => \N__24911\
        );

    \I__5445\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24908\
        );

    \I__5444\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24905\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__24930\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__24927\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__24924\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__24919\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5439\ : Odrv12
    port map (
            O => \N__24916\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5438\ : Odrv4
    port map (
            O => \N__24911\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__24908\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__24905\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__24888\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_10_cascade_\
        );

    \I__5434\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24882\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__24882\,
            I => \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0\
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__24879\,
            I => \N__24876\
        );

    \I__5431\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24871\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__24875\,
            I => \N__24868\
        );

    \I__5429\ : CascadeMux
    port map (
            O => \N__24874\,
            I => \N__24865\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__24871\,
            I => \N__24861\
        );

    \I__5427\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24858\
        );

    \I__5426\ : InMux
    port map (
            O => \N__24865\,
            I => \N__24855\
        );

    \I__5425\ : CascadeMux
    port map (
            O => \N__24864\,
            I => \N__24852\
        );

    \I__5424\ : Span4Mux_h
    port map (
            O => \N__24861\,
            I => \N__24844\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__24858\,
            I => \N__24844\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__24855\,
            I => \N__24841\
        );

    \I__5421\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24838\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__24851\,
            I => \N__24835\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__24850\,
            I => \N__24832\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__24849\,
            I => \N__24827\
        );

    \I__5417\ : Span4Mux_v
    port map (
            O => \N__24844\,
            I => \N__24818\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__24841\,
            I => \N__24818\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__24838\,
            I => \N__24818\
        );

    \I__5414\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24815\
        );

    \I__5413\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24812\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__24831\,
            I => \N__24808\
        );

    \I__5411\ : CascadeMux
    port map (
            O => \N__24830\,
            I => \N__24803\
        );

    \I__5410\ : InMux
    port map (
            O => \N__24827\,
            I => \N__24800\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__24826\,
            I => \N__24797\
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__24825\,
            I => \N__24794\
        );

    \I__5407\ : Span4Mux_v
    port map (
            O => \N__24818\,
            I => \N__24788\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24788\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__24812\,
            I => \N__24785\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__24811\,
            I => \N__24782\
        );

    \I__5403\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24779\
        );

    \I__5402\ : CascadeMux
    port map (
            O => \N__24807\,
            I => \N__24776\
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__24806\,
            I => \N__24773\
        );

    \I__5400\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24770\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__24800\,
            I => \N__24767\
        );

    \I__5398\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24764\
        );

    \I__5397\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24761\
        );

    \I__5396\ : CascadeMux
    port map (
            O => \N__24793\,
            I => \N__24758\
        );

    \I__5395\ : Span4Mux_v
    port map (
            O => \N__24788\,
            I => \N__24753\
        );

    \I__5394\ : Span4Mux_h
    port map (
            O => \N__24785\,
            I => \N__24753\
        );

    \I__5393\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24750\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24747\
        );

    \I__5391\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24744\
        );

    \I__5390\ : InMux
    port map (
            O => \N__24773\,
            I => \N__24741\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__24770\,
            I => \N__24737\
        );

    \I__5388\ : Span4Mux_h
    port map (
            O => \N__24767\,
            I => \N__24732\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__24764\,
            I => \N__24732\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__24761\,
            I => \N__24729\
        );

    \I__5385\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24726\
        );

    \I__5384\ : Span4Mux_v
    port map (
            O => \N__24753\,
            I => \N__24721\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__24750\,
            I => \N__24721\
        );

    \I__5382\ : Span4Mux_v
    port map (
            O => \N__24747\,
            I => \N__24714\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__24744\,
            I => \N__24714\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__24741\,
            I => \N__24714\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__24740\,
            I => \N__24711\
        );

    \I__5378\ : Sp12to4
    port map (
            O => \N__24737\,
            I => \N__24708\
        );

    \I__5377\ : Span4Mux_v
    port map (
            O => \N__24732\,
            I => \N__24705\
        );

    \I__5376\ : Span12Mux_h
    port map (
            O => \N__24729\,
            I => \N__24702\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__24726\,
            I => \N__24699\
        );

    \I__5374\ : Span4Mux_v
    port map (
            O => \N__24721\,
            I => \N__24694\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__24714\,
            I => \N__24694\
        );

    \I__5372\ : InMux
    port map (
            O => \N__24711\,
            I => \N__24691\
        );

    \I__5371\ : Span12Mux_v
    port map (
            O => \N__24708\,
            I => \N__24683\
        );

    \I__5370\ : Sp12to4
    port map (
            O => \N__24705\,
            I => \N__24683\
        );

    \I__5369\ : Span12Mux_v
    port map (
            O => \N__24702\,
            I => \N__24674\
        );

    \I__5368\ : Span12Mux_h
    port map (
            O => \N__24699\,
            I => \N__24674\
        );

    \I__5367\ : Sp12to4
    port map (
            O => \N__24694\,
            I => \N__24674\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__24691\,
            I => \N__24674\
        );

    \I__5365\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24671\
        );

    \I__5364\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24668\
        );

    \I__5363\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24665\
        );

    \I__5362\ : Odrv12
    port map (
            O => \N__24683\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5361\ : Odrv12
    port map (
            O => \N__24674\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__24671\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__24668\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__24665\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5357\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24651\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__24651\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10\
        );

    \I__5355\ : CascadeMux
    port map (
            O => \N__24648\,
            I => \N__24645\
        );

    \I__5354\ : InMux
    port map (
            O => \N__24645\,
            I => \N__24642\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__24642\,
            I => \N__24639\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__24639\,
            I => \M_this_substate_q_RNOZ0Z_3\
        );

    \I__5351\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24633\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__24633\,
            I => \N__24630\
        );

    \I__5349\ : Span12Mux_h
    port map (
            O => \N__24630\,
            I => \N__24627\
        );

    \I__5348\ : Span12Mux_v
    port map (
            O => \N__24627\,
            I => \N__24624\
        );

    \I__5347\ : Odrv12
    port map (
            O => \N__24624\,
            I => \this_sprites_ram.mem_out_bus0_1\
        );

    \I__5346\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24618\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__24618\,
            I => \N__24615\
        );

    \I__5344\ : Span4Mux_h
    port map (
            O => \N__24615\,
            I => \N__24612\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__24612\,
            I => \N__24609\
        );

    \I__5342\ : Span4Mux_h
    port map (
            O => \N__24609\,
            I => \N__24606\
        );

    \I__5341\ : Span4Mux_h
    port map (
            O => \N__24606\,
            I => \N__24603\
        );

    \I__5340\ : Odrv4
    port map (
            O => \N__24603\,
            I => \this_sprites_ram.mem_out_bus4_1\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__24600\,
            I => \N__24596\
        );

    \I__5338\ : CascadeMux
    port map (
            O => \N__24599\,
            I => \N__24590\
        );

    \I__5337\ : InMux
    port map (
            O => \N__24596\,
            I => \N__24582\
        );

    \I__5336\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24582\
        );

    \I__5335\ : InMux
    port map (
            O => \N__24594\,
            I => \N__24577\
        );

    \I__5334\ : InMux
    port map (
            O => \N__24593\,
            I => \N__24577\
        );

    \I__5333\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24574\
        );

    \I__5332\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24569\
        );

    \I__5331\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24569\
        );

    \I__5330\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24566\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__24582\,
            I => \N__24561\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__24577\,
            I => \N__24561\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__24574\,
            I => \N__24554\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__24569\,
            I => \N__24554\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__24566\,
            I => \N__24554\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__24561\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__24554\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__5322\ : CascadeMux
    port map (
            O => \N__24549\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_\
        );

    \I__5321\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24543\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__24543\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1\
        );

    \I__5319\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24537\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__24537\,
            I => \N__24534\
        );

    \I__5317\ : Span4Mux_h
    port map (
            O => \N__24534\,
            I => \N__24531\
        );

    \I__5316\ : Span4Mux_v
    port map (
            O => \N__24531\,
            I => \N__24528\
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__24528\,
            I => \this_sprites_ram.mem_out_bus6_1\
        );

    \I__5314\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24522\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__24522\,
            I => \N__24519\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__24519\,
            I => \N__24516\
        );

    \I__5311\ : Odrv4
    port map (
            O => \N__24516\,
            I => \this_sprites_ram.mem_out_bus2_1\
        );

    \I__5310\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24510\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__24510\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\
        );

    \I__5308\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24504\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__24504\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12\
        );

    \I__5306\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24498\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__24498\,
            I => \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\
        );

    \I__5304\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24492\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__24492\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0\
        );

    \I__5302\ : InMux
    port map (
            O => \N__24489\,
            I => \N__24486\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__24486\,
            I => \M_this_sprites_address_q_RNIQ61C7Z0Z_0\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__24483\,
            I => \N__24480\
        );

    \I__5299\ : InMux
    port map (
            O => \N__24480\,
            I => \N__24477\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__24477\,
            I => \N__24474\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__24474\,
            I => \N__24471\
        );

    \I__5296\ : Odrv4
    port map (
            O => \N__24471\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_0\
        );

    \I__5295\ : CascadeMux
    port map (
            O => \N__24468\,
            I => \N__24464\
        );

    \I__5294\ : CascadeMux
    port map (
            O => \N__24467\,
            I => \N__24461\
        );

    \I__5293\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24457\
        );

    \I__5292\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24454\
        );

    \I__5291\ : CascadeMux
    port map (
            O => \N__24460\,
            I => \N__24451\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__24457\,
            I => \N__24446\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__24454\,
            I => \N__24443\
        );

    \I__5288\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24440\
        );

    \I__5287\ : CascadeMux
    port map (
            O => \N__24450\,
            I => \N__24437\
        );

    \I__5286\ : CascadeMux
    port map (
            O => \N__24449\,
            I => \N__24434\
        );

    \I__5285\ : Span4Mux_v
    port map (
            O => \N__24446\,
            I => \N__24420\
        );

    \I__5284\ : Span4Mux_h
    port map (
            O => \N__24443\,
            I => \N__24420\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__24440\,
            I => \N__24420\
        );

    \I__5282\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24417\
        );

    \I__5281\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24414\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__24433\,
            I => \N__24411\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__24432\,
            I => \N__24408\
        );

    \I__5278\ : CascadeMux
    port map (
            O => \N__24431\,
            I => \N__24405\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__24430\,
            I => \N__24400\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__24429\,
            I => \N__24397\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__24428\,
            I => \N__24394\
        );

    \I__5274\ : CascadeMux
    port map (
            O => \N__24427\,
            I => \N__24391\
        );

    \I__5273\ : Span4Mux_v
    port map (
            O => \N__24420\,
            I => \N__24385\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__24417\,
            I => \N__24385\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__24414\,
            I => \N__24382\
        );

    \I__5270\ : InMux
    port map (
            O => \N__24411\,
            I => \N__24379\
        );

    \I__5269\ : InMux
    port map (
            O => \N__24408\,
            I => \N__24376\
        );

    \I__5268\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24373\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__24404\,
            I => \N__24370\
        );

    \I__5266\ : CascadeMux
    port map (
            O => \N__24403\,
            I => \N__24367\
        );

    \I__5265\ : InMux
    port map (
            O => \N__24400\,
            I => \N__24364\
        );

    \I__5264\ : InMux
    port map (
            O => \N__24397\,
            I => \N__24361\
        );

    \I__5263\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24358\
        );

    \I__5262\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24355\
        );

    \I__5261\ : CascadeMux
    port map (
            O => \N__24390\,
            I => \N__24352\
        );

    \I__5260\ : Span4Mux_v
    port map (
            O => \N__24385\,
            I => \N__24345\
        );

    \I__5259\ : Span4Mux_h
    port map (
            O => \N__24382\,
            I => \N__24345\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__24379\,
            I => \N__24345\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__24376\,
            I => \N__24340\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__24373\,
            I => \N__24340\
        );

    \I__5255\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24337\
        );

    \I__5254\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24334\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__24364\,
            I => \N__24325\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__24361\,
            I => \N__24325\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__24358\,
            I => \N__24325\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__24355\,
            I => \N__24322\
        );

    \I__5249\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24319\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__24345\,
            I => \N__24316\
        );

    \I__5247\ : Span4Mux_v
    port map (
            O => \N__24340\,
            I => \N__24309\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__24337\,
            I => \N__24309\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__24334\,
            I => \N__24309\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__24333\,
            I => \N__24306\
        );

    \I__5243\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24303\
        );

    \I__5242\ : Span12Mux_v
    port map (
            O => \N__24325\,
            I => \N__24300\
        );

    \I__5241\ : Span12Mux_h
    port map (
            O => \N__24322\,
            I => \N__24297\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__24319\,
            I => \N__24294\
        );

    \I__5239\ : Span4Mux_v
    port map (
            O => \N__24316\,
            I => \N__24289\
        );

    \I__5238\ : Span4Mux_v
    port map (
            O => \N__24309\,
            I => \N__24289\
        );

    \I__5237\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24286\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__24303\,
            I => \N__24283\
        );

    \I__5235\ : Span12Mux_h
    port map (
            O => \N__24300\,
            I => \N__24278\
        );

    \I__5234\ : Span12Mux_v
    port map (
            O => \N__24297\,
            I => \N__24269\
        );

    \I__5233\ : Span12Mux_h
    port map (
            O => \N__24294\,
            I => \N__24269\
        );

    \I__5232\ : Sp12to4
    port map (
            O => \N__24289\,
            I => \N__24269\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__24286\,
            I => \N__24269\
        );

    \I__5230\ : Span4Mux_h
    port map (
            O => \N__24283\,
            I => \N__24266\
        );

    \I__5229\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24263\
        );

    \I__5228\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24260\
        );

    \I__5227\ : Odrv12
    port map (
            O => \N__24278\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5226\ : Odrv12
    port map (
            O => \N__24269\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5225\ : Odrv4
    port map (
            O => \N__24266\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__24263\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__24260\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5222\ : CascadeMux
    port map (
            O => \N__24249\,
            I => \N__24246\
        );

    \I__5221\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24243\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__24243\,
            I => \N__24240\
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__24240\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_11\
        );

    \I__5218\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24234\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__24234\,
            I => \N__24231\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__24231\,
            I => \M_this_substate_q_RNOZ0Z_1\
        );

    \I__5215\ : InMux
    port map (
            O => \N__24228\,
            I => \N__24225\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__24225\,
            I => \N__24222\
        );

    \I__5213\ : Odrv12
    port map (
            O => \N__24222\,
            I => \M_this_substate_q_s_1\
        );

    \I__5212\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24215\
        );

    \I__5211\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24212\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__24215\,
            I => \N__24209\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__24212\,
            I => \this_vga_signals_M_this_state_d_2_sqmuxa_0\
        );

    \I__5208\ : Odrv4
    port map (
            O => \N__24209\,
            I => \this_vga_signals_M_this_state_d_2_sqmuxa_0\
        );

    \I__5207\ : InMux
    port map (
            O => \N__24204\,
            I => \N__24201\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__24201\,
            I => \N__24196\
        );

    \I__5205\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24193\
        );

    \I__5204\ : InMux
    port map (
            O => \N__24199\,
            I => \N__24190\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__24196\,
            I => \N_17_0\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__24193\,
            I => \N_17_0\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__24190\,
            I => \N_17_0\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__24183\,
            I => \N__24179\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__24182\,
            I => \N__24173\
        );

    \I__5198\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24170\
        );

    \I__5197\ : CascadeMux
    port map (
            O => \N__24178\,
            I => \N__24167\
        );

    \I__5196\ : CascadeMux
    port map (
            O => \N__24177\,
            I => \N__24160\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__24176\,
            I => \N__24156\
        );

    \I__5194\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24152\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__24170\,
            I => \N__24149\
        );

    \I__5192\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24146\
        );

    \I__5191\ : CascadeMux
    port map (
            O => \N__24166\,
            I => \N__24143\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__24165\,
            I => \N__24140\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__24164\,
            I => \N__24137\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__24163\,
            I => \N__24134\
        );

    \I__5187\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24127\
        );

    \I__5186\ : CascadeMux
    port map (
            O => \N__24159\,
            I => \N__24124\
        );

    \I__5185\ : InMux
    port map (
            O => \N__24156\,
            I => \N__24121\
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__24155\,
            I => \N__24118\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__24152\,
            I => \N__24111\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__24149\,
            I => \N__24111\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__24146\,
            I => \N__24111\
        );

    \I__5180\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24108\
        );

    \I__5179\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24105\
        );

    \I__5178\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24102\
        );

    \I__5177\ : InMux
    port map (
            O => \N__24134\,
            I => \N__24099\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__24133\,
            I => \N__24095\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__24132\,
            I => \N__24092\
        );

    \I__5174\ : CascadeMux
    port map (
            O => \N__24131\,
            I => \N__24089\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__24130\,
            I => \N__24086\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N__24083\
        );

    \I__5171\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24080\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__24121\,
            I => \N__24077\
        );

    \I__5169\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24074\
        );

    \I__5168\ : Span4Mux_v
    port map (
            O => \N__24111\,
            I => \N__24067\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24067\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__24105\,
            I => \N__24067\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__24102\,
            I => \N__24062\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__24099\,
            I => \N__24062\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__24098\,
            I => \N__24059\
        );

    \I__5162\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24056\
        );

    \I__5161\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24053\
        );

    \I__5160\ : InMux
    port map (
            O => \N__24089\,
            I => \N__24050\
        );

    \I__5159\ : InMux
    port map (
            O => \N__24086\,
            I => \N__24047\
        );

    \I__5158\ : Span4Mux_v
    port map (
            O => \N__24083\,
            I => \N__24042\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__24080\,
            I => \N__24042\
        );

    \I__5156\ : Span4Mux_h
    port map (
            O => \N__24077\,
            I => \N__24039\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24035\
        );

    \I__5154\ : Span4Mux_v
    port map (
            O => \N__24067\,
            I => \N__24030\
        );

    \I__5153\ : Span4Mux_v
    port map (
            O => \N__24062\,
            I => \N__24030\
        );

    \I__5152\ : InMux
    port map (
            O => \N__24059\,
            I => \N__24026\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__24056\,
            I => \N__24023\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__24053\,
            I => \N__24020\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__24050\,
            I => \N__24017\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__24047\,
            I => \N__24014\
        );

    \I__5147\ : Span4Mux_h
    port map (
            O => \N__24042\,
            I => \N__24009\
        );

    \I__5146\ : Span4Mux_v
    port map (
            O => \N__24039\,
            I => \N__24009\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__24038\,
            I => \N__24006\
        );

    \I__5144\ : Span4Mux_h
    port map (
            O => \N__24035\,
            I => \N__24003\
        );

    \I__5143\ : Sp12to4
    port map (
            O => \N__24030\,
            I => \N__24000\
        );

    \I__5142\ : InMux
    port map (
            O => \N__24029\,
            I => \N__23996\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__24026\,
            I => \N__23989\
        );

    \I__5140\ : Span4Mux_v
    port map (
            O => \N__24023\,
            I => \N__23989\
        );

    \I__5139\ : Span4Mux_v
    port map (
            O => \N__24020\,
            I => \N__23989\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__24017\,
            I => \N__23986\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__24014\,
            I => \N__23981\
        );

    \I__5136\ : Span4Mux_v
    port map (
            O => \N__24009\,
            I => \N__23981\
        );

    \I__5135\ : InMux
    port map (
            O => \N__24006\,
            I => \N__23978\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__24003\,
            I => \N__23975\
        );

    \I__5133\ : Span12Mux_h
    port map (
            O => \N__24000\,
            I => \N__23972\
        );

    \I__5132\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23969\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__23996\,
            I => \N__23962\
        );

    \I__5130\ : Span4Mux_h
    port map (
            O => \N__23989\,
            I => \N__23962\
        );

    \I__5129\ : Span4Mux_v
    port map (
            O => \N__23986\,
            I => \N__23962\
        );

    \I__5128\ : Span4Mux_h
    port map (
            O => \N__23981\,
            I => \N__23959\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__23978\,
            I => \N__23956\
        );

    \I__5126\ : Sp12to4
    port map (
            O => \N__23975\,
            I => \N__23951\
        );

    \I__5125\ : Span12Mux_v
    port map (
            O => \N__23972\,
            I => \N__23951\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__23969\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__23962\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__23959\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__23956\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5120\ : Odrv12
    port map (
            O => \N__23951\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5119\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23937\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__23937\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_3\
        );

    \I__5117\ : CascadeMux
    port map (
            O => \N__23934\,
            I => \N__23931\
        );

    \I__5116\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23928\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__23928\,
            I => \N__23925\
        );

    \I__5114\ : Odrv12
    port map (
            O => \N__23925\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_12\
        );

    \I__5113\ : CascadeMux
    port map (
            O => \N__23922\,
            I => \N__23919\
        );

    \I__5112\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23916\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__23916\,
            I => \N__23913\
        );

    \I__5110\ : Odrv12
    port map (
            O => \N__23913\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_13\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__23910\,
            I => \N__23907\
        );

    \I__5108\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23901\
        );

    \I__5107\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23898\
        );

    \I__5106\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23893\
        );

    \I__5105\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23893\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__23901\,
            I => \this_ppu.N_1046_0\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__23898\,
            I => \this_ppu.N_1046_0\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__23893\,
            I => \this_ppu.N_1046_0\
        );

    \I__5101\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23882\
        );

    \I__5100\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23879\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__23882\,
            I => \this_ppu.un1_M_oam_idx_q_1_c1\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__23879\,
            I => \this_ppu.un1_M_oam_idx_q_1_c1\
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__23874\,
            I => \N__23871\
        );

    \I__5096\ : CascadeBuf
    port map (
            O => \N__23871\,
            I => \N__23868\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__23868\,
            I => \N__23865\
        );

    \I__5094\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23858\
        );

    \I__5093\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23855\
        );

    \I__5092\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23848\
        );

    \I__5091\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23848\
        );

    \I__5090\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23848\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__23858\,
            I => \N__23845\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__23855\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__23848\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__5086\ : Odrv12
    port map (
            O => \N__23845\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__23838\,
            I => \N__23835\
        );

    \I__5084\ : CascadeBuf
    port map (
            O => \N__23835\,
            I => \N__23832\
        );

    \I__5083\ : CascadeMux
    port map (
            O => \N__23832\,
            I => \N__23829\
        );

    \I__5082\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23826\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__23826\,
            I => \N__23822\
        );

    \I__5080\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23816\
        );

    \I__5079\ : Span4Mux_h
    port map (
            O => \N__23822\,
            I => \N__23813\
        );

    \I__5078\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23810\
        );

    \I__5077\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23805\
        );

    \I__5076\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23805\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__23816\,
            I => \N__23802\
        );

    \I__5074\ : Span4Mux_h
    port map (
            O => \N__23813\,
            I => \N__23799\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__23810\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__23805\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__5071\ : Odrv4
    port map (
            O => \N__23802\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__23799\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__5069\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23787\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__23787\,
            I => \this_ppu.N_144_4\
        );

    \I__5067\ : CascadeMux
    port map (
            O => \N__23784\,
            I => \N__23781\
        );

    \I__5066\ : InMux
    port map (
            O => \N__23781\,
            I => \N__23778\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__23778\,
            I => \N__23775\
        );

    \I__5064\ : Span4Mux_h
    port map (
            O => \N__23775\,
            I => \N__23772\
        );

    \I__5063\ : Odrv4
    port map (
            O => \N__23772\,
            I => \this_ppu.N_144\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__23769\,
            I => \N__23764\
        );

    \I__5061\ : InMux
    port map (
            O => \N__23768\,
            I => \N__23760\
        );

    \I__5060\ : CascadeMux
    port map (
            O => \N__23767\,
            I => \N__23757\
        );

    \I__5059\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23754\
        );

    \I__5058\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23751\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__23760\,
            I => \N__23747\
        );

    \I__5056\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23744\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__23754\,
            I => \N__23741\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__23751\,
            I => \N__23738\
        );

    \I__5053\ : CascadeMux
    port map (
            O => \N__23750\,
            I => \N__23735\
        );

    \I__5052\ : Span4Mux_v
    port map (
            O => \N__23747\,
            I => \N__23730\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__23744\,
            I => \N__23730\
        );

    \I__5050\ : Span4Mux_v
    port map (
            O => \N__23741\,
            I => \N__23723\
        );

    \I__5049\ : Span4Mux_v
    port map (
            O => \N__23738\,
            I => \N__23723\
        );

    \I__5048\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23720\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__23730\,
            I => \N__23717\
        );

    \I__5046\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23712\
        );

    \I__5045\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23712\
        );

    \I__5044\ : Odrv4
    port map (
            O => \N__23723\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__23720\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__5042\ : Odrv4
    port map (
            O => \N__23717\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__23712\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__5040\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23698\
        );

    \I__5039\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23694\
        );

    \I__5038\ : InMux
    port map (
            O => \N__23701\,
            I => \N__23691\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__23698\,
            I => \N__23687\
        );

    \I__5036\ : InMux
    port map (
            O => \N__23697\,
            I => \N__23684\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__23694\,
            I => \N__23681\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23678\
        );

    \I__5033\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23674\
        );

    \I__5032\ : Span4Mux_v
    port map (
            O => \N__23687\,
            I => \N__23670\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__23684\,
            I => \N__23663\
        );

    \I__5030\ : Span4Mux_v
    port map (
            O => \N__23681\,
            I => \N__23663\
        );

    \I__5029\ : Span4Mux_v
    port map (
            O => \N__23678\,
            I => \N__23663\
        );

    \I__5028\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23660\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__23674\,
            I => \N__23657\
        );

    \I__5026\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23654\
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__23670\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__23663\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__23660\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__23657\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__23654\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__5020\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23638\
        );

    \I__5019\ : InMux
    port map (
            O => \N__23642\,
            I => \N__23633\
        );

    \I__5018\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23630\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__23638\,
            I => \N__23626\
        );

    \I__5016\ : InMux
    port map (
            O => \N__23637\,
            I => \N__23623\
        );

    \I__5015\ : InMux
    port map (
            O => \N__23636\,
            I => \N__23620\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__23633\,
            I => \N__23615\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__23630\,
            I => \N__23612\
        );

    \I__5012\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23609\
        );

    \I__5011\ : Span12Mux_s8_v
    port map (
            O => \N__23626\,
            I => \N__23602\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__23623\,
            I => \N__23602\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__23620\,
            I => \N__23602\
        );

    \I__5008\ : InMux
    port map (
            O => \N__23619\,
            I => \N__23599\
        );

    \I__5007\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23596\
        );

    \I__5006\ : Span12Mux_v
    port map (
            O => \N__23615\,
            I => \N__23591\
        );

    \I__5005\ : Span12Mux_v
    port map (
            O => \N__23612\,
            I => \N__23591\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__23609\,
            I => \N__23582\
        );

    \I__5003\ : Span12Mux_v
    port map (
            O => \N__23602\,
            I => \N__23582\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__23599\,
            I => \N__23582\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__23596\,
            I => \N__23582\
        );

    \I__5000\ : Span12Mux_h
    port map (
            O => \N__23591\,
            I => \N__23579\
        );

    \I__4999\ : Span12Mux_s11_v
    port map (
            O => \N__23582\,
            I => \N__23576\
        );

    \I__4998\ : Odrv12
    port map (
            O => \N__23579\,
            I => \M_this_sprites_ram_write_data_2\
        );

    \I__4997\ : Odrv12
    port map (
            O => \N__23576\,
            I => \M_this_sprites_ram_write_data_2\
        );

    \I__4996\ : CEMux
    port map (
            O => \N__23571\,
            I => \N__23567\
        );

    \I__4995\ : CEMux
    port map (
            O => \N__23570\,
            I => \N__23564\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__23567\,
            I => \N__23561\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__23564\,
            I => \N__23558\
        );

    \I__4992\ : Span4Mux_h
    port map (
            O => \N__23561\,
            I => \N__23555\
        );

    \I__4991\ : Span4Mux_h
    port map (
            O => \N__23558\,
            I => \N__23552\
        );

    \I__4990\ : Span4Mux_h
    port map (
            O => \N__23555\,
            I => \N__23549\
        );

    \I__4989\ : Span4Mux_h
    port map (
            O => \N__23552\,
            I => \N__23546\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__23549\,
            I => \N__23543\
        );

    \I__4987\ : Span4Mux_h
    port map (
            O => \N__23546\,
            I => \N__23540\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__23543\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__23540\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__4984\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23532\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__23532\,
            I => \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\
        );

    \I__4982\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23526\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__23526\,
            I => \N__23523\
        );

    \I__4980\ : Span4Mux_v
    port map (
            O => \N__23523\,
            I => \N__23520\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__23520\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13\
        );

    \I__4978\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23514\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__23514\,
            I => \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__23511\,
            I => \this_ppu.N_1046_0_cascade_\
        );

    \I__4975\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23501\
        );

    \I__4974\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23496\
        );

    \I__4973\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23496\
        );

    \I__4972\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23491\
        );

    \I__4971\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23491\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__23501\,
            I => \N__23484\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__23496\,
            I => \N__23484\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__23491\,
            I => \N__23484\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__23484\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__23481\,
            I => \this_ppu.un1_M_oam_idx_q_1_c1_cascade_\
        );

    \I__4965\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23472\
        );

    \I__4964\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23472\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__23472\,
            I => \this_ppu.un1_M_oam_idx_q_1_c3\
        );

    \I__4962\ : CascadeMux
    port map (
            O => \N__23469\,
            I => \N__23466\
        );

    \I__4961\ : CascadeBuf
    port map (
            O => \N__23466\,
            I => \N__23463\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__23463\,
            I => \N__23460\
        );

    \I__4959\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23457\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__23457\,
            I => \N__23453\
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__23456\,
            I => \N__23450\
        );

    \I__4956\ : Span4Mux_h
    port map (
            O => \N__23453\,
            I => \N__23445\
        );

    \I__4955\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23442\
        );

    \I__4954\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23437\
        );

    \I__4953\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23437\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__23445\,
            I => \N__23434\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__23442\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__23437\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__4949\ : Odrv4
    port map (
            O => \N__23434\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__4948\ : CascadeMux
    port map (
            O => \N__23427\,
            I => \N__23424\
        );

    \I__4947\ : CascadeBuf
    port map (
            O => \N__23424\,
            I => \N__23421\
        );

    \I__4946\ : CascadeMux
    port map (
            O => \N__23421\,
            I => \N__23417\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__23420\,
            I => \N__23414\
        );

    \I__4944\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23409\
        );

    \I__4943\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23402\
        );

    \I__4942\ : InMux
    port map (
            O => \N__23413\,
            I => \N__23402\
        );

    \I__4941\ : InMux
    port map (
            O => \N__23412\,
            I => \N__23402\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23399\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__23402\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__4938\ : Odrv12
    port map (
            O => \N__23399\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__23394\,
            I => \N__23390\
        );

    \I__4936\ : InMux
    port map (
            O => \N__23393\,
            I => \N__23387\
        );

    \I__4935\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23384\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__23387\,
            I => \this_ppu.M_oam_idx_qZ0Z_4\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__23384\,
            I => \this_ppu.M_oam_idx_qZ0Z_4\
        );

    \I__4932\ : CascadeMux
    port map (
            O => \N__23379\,
            I => \this_ppu.N_144_4_cascade_\
        );

    \I__4931\ : InMux
    port map (
            O => \N__23376\,
            I => \N__23373\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__23373\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__4929\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23367\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__23367\,
            I => \N__23362\
        );

    \I__4927\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23359\
        );

    \I__4926\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23356\
        );

    \I__4925\ : Odrv4
    port map (
            O => \N__23362\,
            I => \this_ppu.N_156\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__23359\,
            I => \this_ppu.N_156\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__23356\,
            I => \this_ppu.N_156\
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__23349\,
            I => \this_ppu.un2_hscroll_axb_0_cascade_\
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__23346\,
            I => \N__23340\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__23345\,
            I => \N__23335\
        );

    \I__4919\ : CascadeMux
    port map (
            O => \N__23344\,
            I => \N__23329\
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__23343\,
            I => \N__23326\
        );

    \I__4917\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23321\
        );

    \I__4916\ : CascadeMux
    port map (
            O => \N__23339\,
            I => \N__23318\
        );

    \I__4915\ : CascadeMux
    port map (
            O => \N__23338\,
            I => \N__23315\
        );

    \I__4914\ : InMux
    port map (
            O => \N__23335\,
            I => \N__23310\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__23334\,
            I => \N__23307\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__23333\,
            I => \N__23304\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__23332\,
            I => \N__23301\
        );

    \I__4910\ : InMux
    port map (
            O => \N__23329\,
            I => \N__23298\
        );

    \I__4909\ : InMux
    port map (
            O => \N__23326\,
            I => \N__23295\
        );

    \I__4908\ : CascadeMux
    port map (
            O => \N__23325\,
            I => \N__23292\
        );

    \I__4907\ : CascadeMux
    port map (
            O => \N__23324\,
            I => \N__23289\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23285\
        );

    \I__4905\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23282\
        );

    \I__4904\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23279\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__23314\,
            I => \N__23276\
        );

    \I__4902\ : CascadeMux
    port map (
            O => \N__23313\,
            I => \N__23273\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__23310\,
            I => \N__23268\
        );

    \I__4900\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23265\
        );

    \I__4899\ : InMux
    port map (
            O => \N__23304\,
            I => \N__23262\
        );

    \I__4898\ : InMux
    port map (
            O => \N__23301\,
            I => \N__23259\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__23298\,
            I => \N__23254\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__23295\,
            I => \N__23254\
        );

    \I__4895\ : InMux
    port map (
            O => \N__23292\,
            I => \N__23251\
        );

    \I__4894\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23248\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__23288\,
            I => \N__23245\
        );

    \I__4892\ : Span4Mux_s2_v
    port map (
            O => \N__23285\,
            I => \N__23240\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__23282\,
            I => \N__23240\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23237\
        );

    \I__4889\ : InMux
    port map (
            O => \N__23276\,
            I => \N__23234\
        );

    \I__4888\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23231\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__23272\,
            I => \N__23228\
        );

    \I__4886\ : CascadeMux
    port map (
            O => \N__23271\,
            I => \N__23225\
        );

    \I__4885\ : Span4Mux_v
    port map (
            O => \N__23268\,
            I => \N__23220\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__23265\,
            I => \N__23220\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__23262\,
            I => \N__23217\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__23259\,
            I => \N__23214\
        );

    \I__4881\ : Span4Mux_v
    port map (
            O => \N__23254\,
            I => \N__23207\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23207\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__23248\,
            I => \N__23207\
        );

    \I__4878\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23204\
        );

    \I__4877\ : Span4Mux_v
    port map (
            O => \N__23240\,
            I => \N__23197\
        );

    \I__4876\ : Span4Mux_h
    port map (
            O => \N__23237\,
            I => \N__23197\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__23234\,
            I => \N__23197\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__23231\,
            I => \N__23194\
        );

    \I__4873\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23191\
        );

    \I__4872\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23188\
        );

    \I__4871\ : Span4Mux_v
    port map (
            O => \N__23220\,
            I => \N__23181\
        );

    \I__4870\ : Span4Mux_v
    port map (
            O => \N__23217\,
            I => \N__23181\
        );

    \I__4869\ : Span4Mux_v
    port map (
            O => \N__23214\,
            I => \N__23181\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__23207\,
            I => \N__23176\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__23204\,
            I => \N__23176\
        );

    \I__4866\ : Span4Mux_v
    port map (
            O => \N__23197\,
            I => \N__23169\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__23194\,
            I => \N__23169\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__23191\,
            I => \N__23169\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__23188\,
            I => \N__23166\
        );

    \I__4862\ : Span4Mux_h
    port map (
            O => \N__23181\,
            I => \N__23163\
        );

    \I__4861\ : Span4Mux_h
    port map (
            O => \N__23176\,
            I => \N__23160\
        );

    \I__4860\ : Span4Mux_v
    port map (
            O => \N__23169\,
            I => \N__23155\
        );

    \I__4859\ : Span4Mux_h
    port map (
            O => \N__23166\,
            I => \N__23155\
        );

    \I__4858\ : Span4Mux_h
    port map (
            O => \N__23163\,
            I => \N__23152\
        );

    \I__4857\ : Span4Mux_v
    port map (
            O => \N__23160\,
            I => \N__23149\
        );

    \I__4856\ : Span4Mux_h
    port map (
            O => \N__23155\,
            I => \N__23146\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__23152\,
            I => \M_this_ppu_sprites_addr_0\
        );

    \I__4854\ : Odrv4
    port map (
            O => \N__23149\,
            I => \M_this_ppu_sprites_addr_0\
        );

    \I__4853\ : Odrv4
    port map (
            O => \N__23146\,
            I => \M_this_ppu_sprites_addr_0\
        );

    \I__4852\ : InMux
    port map (
            O => \N__23139\,
            I => \N__23133\
        );

    \I__4851\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23133\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__23133\,
            I => \this_ppu.un1_M_haddress_q_3_c2\
        );

    \I__4849\ : SRMux
    port map (
            O => \N__23130\,
            I => \N__23126\
        );

    \I__4848\ : SRMux
    port map (
            O => \N__23129\,
            I => \N__23123\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__23126\,
            I => \this_ppu.M_state_q_RNIGL6V4Z0Z_0\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__23123\,
            I => \this_ppu.M_state_q_RNIGL6V4Z0Z_0\
        );

    \I__4845\ : CEMux
    port map (
            O => \N__23118\,
            I => \N__23115\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__23115\,
            I => \N__23111\
        );

    \I__4843\ : CEMux
    port map (
            O => \N__23114\,
            I => \N__23108\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__23111\,
            I => \N__23105\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__23108\,
            I => \N__23102\
        );

    \I__4840\ : Span4Mux_h
    port map (
            O => \N__23105\,
            I => \N__23099\
        );

    \I__4839\ : Span4Mux_h
    port map (
            O => \N__23102\,
            I => \N__23096\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__23099\,
            I => \N__23093\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__23096\,
            I => \N__23090\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__23093\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__23090\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__4834\ : CEMux
    port map (
            O => \N__23085\,
            I => \N__23081\
        );

    \I__4833\ : CEMux
    port map (
            O => \N__23084\,
            I => \N__23078\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__23081\,
            I => \N__23073\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__23078\,
            I => \N__23073\
        );

    \I__4830\ : Span4Mux_v
    port map (
            O => \N__23073\,
            I => \N__23070\
        );

    \I__4829\ : Span4Mux_v
    port map (
            O => \N__23070\,
            I => \N__23067\
        );

    \I__4828\ : Span4Mux_h
    port map (
            O => \N__23067\,
            I => \N__23064\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__23064\,
            I => \this_sprites_ram.mem_WE_14\
        );

    \I__4826\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__23055\
        );

    \I__4824\ : Span12Mux_h
    port map (
            O => \N__23055\,
            I => \N__23052\
        );

    \I__4823\ : Span12Mux_v
    port map (
            O => \N__23052\,
            I => \N__23049\
        );

    \I__4822\ : Odrv12
    port map (
            O => \N__23049\,
            I => \this_sprites_ram.mem_out_bus7_1\
        );

    \I__4821\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23043\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__23043\,
            I => \N__23040\
        );

    \I__4819\ : Span4Mux_h
    port map (
            O => \N__23040\,
            I => \N__23037\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__23037\,
            I => \this_sprites_ram.mem_out_bus3_1\
        );

    \I__4817\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23031\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__23031\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\
        );

    \I__4815\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23025\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__23025\,
            I => \N__23022\
        );

    \I__4813\ : Span12Mux_v
    port map (
            O => \N__23022\,
            I => \N__23019\
        );

    \I__4812\ : Span12Mux_h
    port map (
            O => \N__23019\,
            I => \N__23016\
        );

    \I__4811\ : Odrv12
    port map (
            O => \N__23016\,
            I => \this_sprites_ram.mem_out_bus4_3\
        );

    \I__4810\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23010\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__23010\,
            I => \N__23007\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__23007\,
            I => \N__23004\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__23004\,
            I => \N__23001\
        );

    \I__4806\ : Span4Mux_v
    port map (
            O => \N__23001\,
            I => \N__22998\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__22998\,
            I => \this_sprites_ram.mem_out_bus0_3\
        );

    \I__4804\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22992\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__22992\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\
        );

    \I__4802\ : InMux
    port map (
            O => \N__22989\,
            I => \N__22985\
        );

    \I__4801\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22982\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__22985\,
            I => \N__22979\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__22982\,
            I => \N__22975\
        );

    \I__4798\ : Span4Mux_h
    port map (
            O => \N__22979\,
            I => \N__22972\
        );

    \I__4797\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22969\
        );

    \I__4796\ : Span4Mux_h
    port map (
            O => \N__22975\,
            I => \N__22966\
        );

    \I__4795\ : Span4Mux_v
    port map (
            O => \N__22972\,
            I => \N__22963\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__22969\,
            I => \N__22960\
        );

    \I__4793\ : Span4Mux_v
    port map (
            O => \N__22966\,
            I => \N__22957\
        );

    \I__4792\ : Sp12to4
    port map (
            O => \N__22963\,
            I => \N__22949\
        );

    \I__4791\ : Span12Mux_v
    port map (
            O => \N__22960\,
            I => \N__22949\
        );

    \I__4790\ : Sp12to4
    port map (
            O => \N__22957\,
            I => \N__22949\
        );

    \I__4789\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22946\
        );

    \I__4788\ : Odrv12
    port map (
            O => \N__22949\,
            I => this_vga_signals_vvisibility
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__22946\,
            I => this_vga_signals_vvisibility
        );

    \I__4786\ : IoInMux
    port map (
            O => \N__22941\,
            I => \N__22938\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__22938\,
            I => \N__22935\
        );

    \I__4784\ : Span4Mux_s2_h
    port map (
            O => \N__22935\,
            I => \N__22932\
        );

    \I__4783\ : Span4Mux_v
    port map (
            O => \N__22932\,
            I => \N__22927\
        );

    \I__4782\ : InMux
    port map (
            O => \N__22931\,
            I => \N__22924\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__22930\,
            I => \N__22920\
        );

    \I__4780\ : Sp12to4
    port map (
            O => \N__22927\,
            I => \N__22917\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__22924\,
            I => \N__22914\
        );

    \I__4778\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22911\
        );

    \I__4777\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22908\
        );

    \I__4776\ : Span12Mux_h
    port map (
            O => \N__22917\,
            I => \N__22905\
        );

    \I__4775\ : Span12Mux_v
    port map (
            O => \N__22914\,
            I => \N__22902\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__22911\,
            I => \N__22898\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__22908\,
            I => \N__22895\
        );

    \I__4772\ : Span12Mux_v
    port map (
            O => \N__22905\,
            I => \N__22890\
        );

    \I__4771\ : Span12Mux_h
    port map (
            O => \N__22902\,
            I => \N__22890\
        );

    \I__4770\ : InMux
    port map (
            O => \N__22901\,
            I => \N__22887\
        );

    \I__4769\ : Span12Mux_s7_h
    port map (
            O => \N__22898\,
            I => \N__22882\
        );

    \I__4768\ : Span12Mux_v
    port map (
            O => \N__22895\,
            I => \N__22882\
        );

    \I__4767\ : Odrv12
    port map (
            O => \N__22890\,
            I => dma_0
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__22887\,
            I => dma_0
        );

    \I__4765\ : Odrv12
    port map (
            O => \N__22882\,
            I => dma_0
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__22875\,
            I => \this_ppu.N_150_cascade_\
        );

    \I__4763\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22867\
        );

    \I__4762\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22864\
        );

    \I__4761\ : InMux
    port map (
            O => \N__22870\,
            I => \N__22855\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__22867\,
            I => \N__22850\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__22864\,
            I => \N__22850\
        );

    \I__4758\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22839\
        );

    \I__4757\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22839\
        );

    \I__4756\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22839\
        );

    \I__4755\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22839\
        );

    \I__4754\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22839\
        );

    \I__4753\ : IoInMux
    port map (
            O => \N__22858\,
            I => \N__22836\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__22855\,
            I => \N__22833\
        );

    \I__4751\ : Span4Mux_v
    port map (
            O => \N__22850\,
            I => \N__22830\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__22839\,
            I => \N__22827\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__22836\,
            I => \N__22823\
        );

    \I__4748\ : Span4Mux_h
    port map (
            O => \N__22833\,
            I => \N__22820\
        );

    \I__4747\ : Span4Mux_h
    port map (
            O => \N__22830\,
            I => \N__22815\
        );

    \I__4746\ : Span4Mux_h
    port map (
            O => \N__22827\,
            I => \N__22815\
        );

    \I__4745\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22812\
        );

    \I__4744\ : Span12Mux_s5_v
    port map (
            O => \N__22823\,
            I => \N__22809\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__22820\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__22815\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__22812\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4740\ : Odrv12
    port map (
            O => \N__22809\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__22800\,
            I => \N__22795\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__22799\,
            I => \N__22790\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__22798\,
            I => \N__22787\
        );

    \I__4736\ : InMux
    port map (
            O => \N__22795\,
            I => \N__22782\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__22794\,
            I => \N__22779\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__22793\,
            I => \N__22776\
        );

    \I__4733\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22767\
        );

    \I__4732\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22764\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__22786\,
            I => \N__22761\
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__22785\,
            I => \N__22758\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__22782\,
            I => \N__22754\
        );

    \I__4728\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22751\
        );

    \I__4727\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22748\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__22775\,
            I => \N__22745\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__22774\,
            I => \N__22742\
        );

    \I__4724\ : CascadeMux
    port map (
            O => \N__22773\,
            I => \N__22737\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__22772\,
            I => \N__22734\
        );

    \I__4722\ : CascadeMux
    port map (
            O => \N__22771\,
            I => \N__22731\
        );

    \I__4721\ : CascadeMux
    port map (
            O => \N__22770\,
            I => \N__22728\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__22767\,
            I => \N__22723\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__22764\,
            I => \N__22723\
        );

    \I__4718\ : InMux
    port map (
            O => \N__22761\,
            I => \N__22720\
        );

    \I__4717\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22717\
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__22757\,
            I => \N__22714\
        );

    \I__4715\ : Span4Mux_v
    port map (
            O => \N__22754\,
            I => \N__22707\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__22751\,
            I => \N__22707\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__22748\,
            I => \N__22707\
        );

    \I__4712\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22704\
        );

    \I__4711\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22701\
        );

    \I__4710\ : CascadeMux
    port map (
            O => \N__22741\,
            I => \N__22698\
        );

    \I__4709\ : CascadeMux
    port map (
            O => \N__22740\,
            I => \N__22695\
        );

    \I__4708\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22692\
        );

    \I__4707\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22689\
        );

    \I__4706\ : InMux
    port map (
            O => \N__22731\,
            I => \N__22686\
        );

    \I__4705\ : InMux
    port map (
            O => \N__22728\,
            I => \N__22683\
        );

    \I__4704\ : Span4Mux_v
    port map (
            O => \N__22723\,
            I => \N__22676\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__22720\,
            I => \N__22676\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__22717\,
            I => \N__22676\
        );

    \I__4701\ : InMux
    port map (
            O => \N__22714\,
            I => \N__22673\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__22707\,
            I => \N__22666\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22666\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__22701\,
            I => \N__22666\
        );

    \I__4697\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22663\
        );

    \I__4696\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22660\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__22692\,
            I => \N__22653\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__22689\,
            I => \N__22653\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__22686\,
            I => \N__22653\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22650\
        );

    \I__4691\ : Span4Mux_v
    port map (
            O => \N__22676\,
            I => \N__22645\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__22673\,
            I => \N__22645\
        );

    \I__4689\ : Span4Mux_v
    port map (
            O => \N__22666\,
            I => \N__22640\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__22663\,
            I => \N__22640\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__22660\,
            I => \N__22637\
        );

    \I__4686\ : Span12Mux_v
    port map (
            O => \N__22653\,
            I => \N__22632\
        );

    \I__4685\ : Span12Mux_v
    port map (
            O => \N__22650\,
            I => \N__22632\
        );

    \I__4684\ : Span4Mux_v
    port map (
            O => \N__22645\,
            I => \N__22627\
        );

    \I__4683\ : Span4Mux_v
    port map (
            O => \N__22640\,
            I => \N__22627\
        );

    \I__4682\ : Span12Mux_h
    port map (
            O => \N__22637\,
            I => \N__22622\
        );

    \I__4681\ : Span12Mux_h
    port map (
            O => \N__22632\,
            I => \N__22622\
        );

    \I__4680\ : Span4Mux_h
    port map (
            O => \N__22627\,
            I => \N__22619\
        );

    \I__4679\ : Odrv12
    port map (
            O => \N__22622\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__22619\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__4677\ : CEMux
    port map (
            O => \N__22614\,
            I => \N__22611\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__22611\,
            I => \N__22608\
        );

    \I__4675\ : Span12Mux_h
    port map (
            O => \N__22608\,
            I => \N__22602\
        );

    \I__4674\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22597\
        );

    \I__4673\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22597\
        );

    \I__4672\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22594\
        );

    \I__4671\ : Odrv12
    port map (
            O => \N__22602\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__22597\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__22594\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4668\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22584\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__22584\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__22581\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_9_cascade_\
        );

    \I__4665\ : InMux
    port map (
            O => \N__22578\,
            I => \N__22575\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__22575\,
            I => \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\
        );

    \I__4663\ : CascadeMux
    port map (
            O => \N__22572\,
            I => \N__22565\
        );

    \I__4662\ : CascadeMux
    port map (
            O => \N__22571\,
            I => \N__22562\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__22570\,
            I => \N__22555\
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__22569\,
            I => \N__22549\
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__22568\,
            I => \N__22545\
        );

    \I__4658\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22542\
        );

    \I__4657\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22539\
        );

    \I__4656\ : CascadeMux
    port map (
            O => \N__22561\,
            I => \N__22536\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__22560\,
            I => \N__22533\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__22559\,
            I => \N__22530\
        );

    \I__4653\ : CascadeMux
    port map (
            O => \N__22558\,
            I => \N__22527\
        );

    \I__4652\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22524\
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__22554\,
            I => \N__22521\
        );

    \I__4650\ : CascadeMux
    port map (
            O => \N__22553\,
            I => \N__22517\
        );

    \I__4649\ : CascadeMux
    port map (
            O => \N__22552\,
            I => \N__22514\
        );

    \I__4648\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22511\
        );

    \I__4647\ : CascadeMux
    port map (
            O => \N__22548\,
            I => \N__22508\
        );

    \I__4646\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22505\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__22542\,
            I => \N__22500\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__22539\,
            I => \N__22500\
        );

    \I__4643\ : InMux
    port map (
            O => \N__22536\,
            I => \N__22497\
        );

    \I__4642\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22494\
        );

    \I__4641\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22491\
        );

    \I__4640\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22488\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__22524\,
            I => \N__22485\
        );

    \I__4638\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22482\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__22520\,
            I => \N__22479\
        );

    \I__4636\ : InMux
    port map (
            O => \N__22517\,
            I => \N__22475\
        );

    \I__4635\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22472\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__22511\,
            I => \N__22469\
        );

    \I__4633\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22466\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__22505\,
            I => \N__22459\
        );

    \I__4631\ : Span4Mux_v
    port map (
            O => \N__22500\,
            I => \N__22459\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__22497\,
            I => \N__22459\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__22494\,
            I => \N__22454\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__22491\,
            I => \N__22454\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__22488\,
            I => \N__22451\
        );

    \I__4626\ : Span4Mux_v
    port map (
            O => \N__22485\,
            I => \N__22446\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__22482\,
            I => \N__22446\
        );

    \I__4624\ : InMux
    port map (
            O => \N__22479\,
            I => \N__22443\
        );

    \I__4623\ : CascadeMux
    port map (
            O => \N__22478\,
            I => \N__22439\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__22475\,
            I => \N__22436\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22433\
        );

    \I__4620\ : Span4Mux_h
    port map (
            O => \N__22469\,
            I => \N__22430\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__22466\,
            I => \N__22427\
        );

    \I__4618\ : Span4Mux_v
    port map (
            O => \N__22459\,
            I => \N__22422\
        );

    \I__4617\ : Span4Mux_v
    port map (
            O => \N__22454\,
            I => \N__22422\
        );

    \I__4616\ : Span4Mux_h
    port map (
            O => \N__22451\,
            I => \N__22419\
        );

    \I__4615\ : Span4Mux_v
    port map (
            O => \N__22446\,
            I => \N__22413\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__22443\,
            I => \N__22413\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__22442\,
            I => \N__22410\
        );

    \I__4612\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22407\
        );

    \I__4611\ : Span4Mux_h
    port map (
            O => \N__22436\,
            I => \N__22404\
        );

    \I__4610\ : Span4Mux_h
    port map (
            O => \N__22433\,
            I => \N__22399\
        );

    \I__4609\ : Span4Mux_v
    port map (
            O => \N__22430\,
            I => \N__22399\
        );

    \I__4608\ : Span4Mux_h
    port map (
            O => \N__22427\,
            I => \N__22396\
        );

    \I__4607\ : Sp12to4
    port map (
            O => \N__22422\,
            I => \N__22393\
        );

    \I__4606\ : Span4Mux_h
    port map (
            O => \N__22419\,
            I => \N__22390\
        );

    \I__4605\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22387\
        );

    \I__4604\ : Span4Mux_h
    port map (
            O => \N__22413\,
            I => \N__22384\
        );

    \I__4603\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22381\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__22407\,
            I => \N__22378\
        );

    \I__4601\ : Span4Mux_h
    port map (
            O => \N__22404\,
            I => \N__22374\
        );

    \I__4600\ : Span4Mux_h
    port map (
            O => \N__22399\,
            I => \N__22370\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__22396\,
            I => \N__22367\
        );

    \I__4598\ : Span12Mux_h
    port map (
            O => \N__22393\,
            I => \N__22364\
        );

    \I__4597\ : Sp12to4
    port map (
            O => \N__22390\,
            I => \N__22361\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__22387\,
            I => \N__22356\
        );

    \I__4595\ : Span4Mux_v
    port map (
            O => \N__22384\,
            I => \N__22356\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__22381\,
            I => \N__22351\
        );

    \I__4593\ : Span12Mux_h
    port map (
            O => \N__22378\,
            I => \N__22351\
        );

    \I__4592\ : InMux
    port map (
            O => \N__22377\,
            I => \N__22348\
        );

    \I__4591\ : Span4Mux_h
    port map (
            O => \N__22374\,
            I => \N__22345\
        );

    \I__4590\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22342\
        );

    \I__4589\ : Span4Mux_h
    port map (
            O => \N__22370\,
            I => \N__22339\
        );

    \I__4588\ : Sp12to4
    port map (
            O => \N__22367\,
            I => \N__22334\
        );

    \I__4587\ : Span12Mux_v
    port map (
            O => \N__22364\,
            I => \N__22334\
        );

    \I__4586\ : Span12Mux_v
    port map (
            O => \N__22361\,
            I => \N__22331\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__22356\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4584\ : Odrv12
    port map (
            O => \N__22351\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__22348\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__22345\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__22342\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__22339\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4579\ : Odrv12
    port map (
            O => \N__22334\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4578\ : Odrv12
    port map (
            O => \N__22331\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__4577\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22311\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__22311\,
            I => \N__22308\
        );

    \I__4575\ : Odrv12
    port map (
            O => \N__22308\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2\
        );

    \I__4574\ : CascadeMux
    port map (
            O => \N__22305\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_2_cascade_\
        );

    \I__4573\ : InMux
    port map (
            O => \N__22302\,
            I => \N__22299\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__22299\,
            I => \N__22296\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__22296\,
            I => \un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0\
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__4569\ : InMux
    port map (
            O => \N__22290\,
            I => \N__22286\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__22289\,
            I => \N__22283\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__22286\,
            I => \N__22278\
        );

    \I__4566\ : InMux
    port map (
            O => \N__22283\,
            I => \N__22275\
        );

    \I__4565\ : CascadeMux
    port map (
            O => \N__22282\,
            I => \N__22272\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__22281\,
            I => \N__22268\
        );

    \I__4563\ : Span4Mux_v
    port map (
            O => \N__22278\,
            I => \N__22260\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__22275\,
            I => \N__22260\
        );

    \I__4561\ : InMux
    port map (
            O => \N__22272\,
            I => \N__22257\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__22271\,
            I => \N__22254\
        );

    \I__4559\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22250\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__22267\,
            I => \N__22247\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__22266\,
            I => \N__22243\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__22265\,
            I => \N__22238\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__22260\,
            I => \N__22232\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__22257\,
            I => \N__22232\
        );

    \I__4553\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22229\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__22253\,
            I => \N__22224\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22221\
        );

    \I__4550\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22218\
        );

    \I__4549\ : CascadeMux
    port map (
            O => \N__22246\,
            I => \N__22215\
        );

    \I__4548\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22212\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__22242\,
            I => \N__22209\
        );

    \I__4546\ : CascadeMux
    port map (
            O => \N__22241\,
            I => \N__22206\
        );

    \I__4545\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22203\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__22237\,
            I => \N__22200\
        );

    \I__4543\ : Span4Mux_v
    port map (
            O => \N__22232\,
            I => \N__22195\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__22229\,
            I => \N__22195\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__22228\,
            I => \N__22192\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__22227\,
            I => \N__22189\
        );

    \I__4539\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22186\
        );

    \I__4538\ : Span4Mux_h
    port map (
            O => \N__22221\,
            I => \N__22180\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__22218\,
            I => \N__22180\
        );

    \I__4536\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22177\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__22212\,
            I => \N__22174\
        );

    \I__4534\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22171\
        );

    \I__4533\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22168\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__22203\,
            I => \N__22165\
        );

    \I__4531\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22162\
        );

    \I__4530\ : Span4Mux_v
    port map (
            O => \N__22195\,
            I => \N__22159\
        );

    \I__4529\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22156\
        );

    \I__4528\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22153\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__22186\,
            I => \N__22150\
        );

    \I__4526\ : CascadeMux
    port map (
            O => \N__22185\,
            I => \N__22147\
        );

    \I__4525\ : Span4Mux_v
    port map (
            O => \N__22180\,
            I => \N__22144\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__22177\,
            I => \N__22141\
        );

    \I__4523\ : Span4Mux_v
    port map (
            O => \N__22174\,
            I => \N__22134\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__22171\,
            I => \N__22134\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__22168\,
            I => \N__22134\
        );

    \I__4520\ : Span12Mux_h
    port map (
            O => \N__22165\,
            I => \N__22129\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__22162\,
            I => \N__22126\
        );

    \I__4518\ : Sp12to4
    port map (
            O => \N__22159\,
            I => \N__22121\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__22156\,
            I => \N__22121\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__22153\,
            I => \N__22118\
        );

    \I__4515\ : Span12Mux_h
    port map (
            O => \N__22150\,
            I => \N__22115\
        );

    \I__4514\ : InMux
    port map (
            O => \N__22147\,
            I => \N__22112\
        );

    \I__4513\ : Span4Mux_h
    port map (
            O => \N__22144\,
            I => \N__22108\
        );

    \I__4512\ : Span4Mux_v
    port map (
            O => \N__22141\,
            I => \N__22103\
        );

    \I__4511\ : Span4Mux_v
    port map (
            O => \N__22134\,
            I => \N__22103\
        );

    \I__4510\ : InMux
    port map (
            O => \N__22133\,
            I => \N__22100\
        );

    \I__4509\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22097\
        );

    \I__4508\ : Span12Mux_v
    port map (
            O => \N__22129\,
            I => \N__22090\
        );

    \I__4507\ : Span12Mux_h
    port map (
            O => \N__22126\,
            I => \N__22090\
        );

    \I__4506\ : Span12Mux_h
    port map (
            O => \N__22121\,
            I => \N__22090\
        );

    \I__4505\ : Span12Mux_s10_h
    port map (
            O => \N__22118\,
            I => \N__22087\
        );

    \I__4504\ : Span12Mux_v
    port map (
            O => \N__22115\,
            I => \N__22082\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__22112\,
            I => \N__22082\
        );

    \I__4502\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22079\
        );

    \I__4501\ : Span4Mux_h
    port map (
            O => \N__22108\,
            I => \N__22072\
        );

    \I__4500\ : Span4Mux_h
    port map (
            O => \N__22103\,
            I => \N__22072\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__22100\,
            I => \N__22072\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__22097\,
            I => \N__22069\
        );

    \I__4497\ : Odrv12
    port map (
            O => \N__22090\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4496\ : Odrv12
    port map (
            O => \N__22087\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4495\ : Odrv12
    port map (
            O => \N__22082\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__22079\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__22072\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__22069\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__22056\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3_cascade_\
        );

    \I__4490\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22050\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__22050\,
            I => \N__22047\
        );

    \I__4488\ : Odrv4
    port map (
            O => \N__22047\,
            I => \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\
        );

    \I__4487\ : CascadeMux
    port map (
            O => \N__22044\,
            I => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_\
        );

    \I__4486\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22038\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__22035\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__22035\,
            I => \un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0\
        );

    \I__4483\ : CascadeMux
    port map (
            O => \N__22032\,
            I => \N__22028\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__22031\,
            I => \N__22025\
        );

    \I__4481\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22018\
        );

    \I__4480\ : InMux
    port map (
            O => \N__22025\,
            I => \N__22015\
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__22024\,
            I => \N__22012\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__22023\,
            I => \N__22009\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__22022\,
            I => \N__22004\
        );

    \I__4476\ : CascadeMux
    port map (
            O => \N__22021\,
            I => \N__22001\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__22018\,
            I => \N__21995\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__22015\,
            I => \N__21995\
        );

    \I__4473\ : InMux
    port map (
            O => \N__22012\,
            I => \N__21992\
        );

    \I__4472\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21989\
        );

    \I__4471\ : CascadeMux
    port map (
            O => \N__22008\,
            I => \N__21986\
        );

    \I__4470\ : CascadeMux
    port map (
            O => \N__22007\,
            I => \N__21983\
        );

    \I__4469\ : InMux
    port map (
            O => \N__22004\,
            I => \N__21979\
        );

    \I__4468\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21976\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__22000\,
            I => \N__21973\
        );

    \I__4466\ : Span4Mux_v
    port map (
            O => \N__21995\,
            I => \N__21965\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__21992\,
            I => \N__21965\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__21989\,
            I => \N__21965\
        );

    \I__4463\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21962\
        );

    \I__4462\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21959\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__21982\,
            I => \N__21956\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__21979\,
            I => \N__21949\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__21976\,
            I => \N__21949\
        );

    \I__4458\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21946\
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__21972\,
            I => \N__21943\
        );

    \I__4456\ : Span4Mux_v
    port map (
            O => \N__21965\,
            I => \N__21936\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__21962\,
            I => \N__21936\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__21959\,
            I => \N__21936\
        );

    \I__4453\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21933\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__21955\,
            I => \N__21928\
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__21954\,
            I => \N__21924\
        );

    \I__4450\ : Span4Mux_v
    port map (
            O => \N__21949\,
            I => \N__21919\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__21946\,
            I => \N__21919\
        );

    \I__4448\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21916\
        );

    \I__4447\ : Span4Mux_v
    port map (
            O => \N__21936\,
            I => \N__21911\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__21933\,
            I => \N__21911\
        );

    \I__4445\ : CascadeMux
    port map (
            O => \N__21932\,
            I => \N__21908\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__21931\,
            I => \N__21905\
        );

    \I__4443\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21902\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__21927\,
            I => \N__21899\
        );

    \I__4441\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21896\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__21919\,
            I => \N__21891\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__21916\,
            I => \N__21891\
        );

    \I__4438\ : Span4Mux_v
    port map (
            O => \N__21911\,
            I => \N__21888\
        );

    \I__4437\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21885\
        );

    \I__4436\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21882\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__21902\,
            I => \N__21879\
        );

    \I__4434\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21876\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__21896\,
            I => \N__21873\
        );

    \I__4432\ : Span4Mux_v
    port map (
            O => \N__21891\,
            I => \N__21870\
        );

    \I__4431\ : Sp12to4
    port map (
            O => \N__21888\,
            I => \N__21867\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__21885\,
            I => \N__21864\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__21882\,
            I => \N__21861\
        );

    \I__4428\ : Span4Mux_v
    port map (
            O => \N__21879\,
            I => \N__21855\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21855\
        );

    \I__4426\ : Span4Mux_s3_v
    port map (
            O => \N__21873\,
            I => \N__21852\
        );

    \I__4425\ : Sp12to4
    port map (
            O => \N__21870\,
            I => \N__21849\
        );

    \I__4424\ : Span12Mux_h
    port map (
            O => \N__21867\,
            I => \N__21846\
        );

    \I__4423\ : Span4Mux_h
    port map (
            O => \N__21864\,
            I => \N__21843\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__21861\,
            I => \N__21840\
        );

    \I__4421\ : InMux
    port map (
            O => \N__21860\,
            I => \N__21835\
        );

    \I__4420\ : Span4Mux_v
    port map (
            O => \N__21855\,
            I => \N__21830\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__21852\,
            I => \N__21830\
        );

    \I__4418\ : Span12Mux_h
    port map (
            O => \N__21849\,
            I => \N__21825\
        );

    \I__4417\ : Span12Mux_v
    port map (
            O => \N__21846\,
            I => \N__21825\
        );

    \I__4416\ : Span4Mux_h
    port map (
            O => \N__21843\,
            I => \N__21820\
        );

    \I__4415\ : Span4Mux_h
    port map (
            O => \N__21840\,
            I => \N__21820\
        );

    \I__4414\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21815\
        );

    \I__4413\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21815\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__21835\,
            I => \N__21812\
        );

    \I__4411\ : Sp12to4
    port map (
            O => \N__21830\,
            I => \N__21807\
        );

    \I__4410\ : Span12Mux_v
    port map (
            O => \N__21825\,
            I => \N__21807\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__21820\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__21815\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__21812\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4406\ : Odrv12
    port map (
            O => \N__21807\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4405\ : InMux
    port map (
            O => \N__21798\,
            I => \N__21795\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__21795\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_7\
        );

    \I__4403\ : InMux
    port map (
            O => \N__21792\,
            I => \N__21789\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__21789\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\
        );

    \I__4401\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21783\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__21783\,
            I => \N__21780\
        );

    \I__4399\ : Span12Mux_v
    port map (
            O => \N__21780\,
            I => \N__21777\
        );

    \I__4398\ : Span12Mux_h
    port map (
            O => \N__21777\,
            I => \N__21773\
        );

    \I__4397\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21770\
        );

    \I__4396\ : Odrv12
    port map (
            O => \N__21773\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__21770\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__4394\ : InMux
    port map (
            O => \N__21765\,
            I => \un1_M_this_sprites_address_q_cry_6\
        );

    \I__4393\ : InMux
    port map (
            O => \N__21762\,
            I => \bfn_19_23_0_\
        );

    \I__4392\ : InMux
    port map (
            O => \N__21759\,
            I => \un1_M_this_sprites_address_q_cry_8\
        );

    \I__4391\ : InMux
    port map (
            O => \N__21756\,
            I => \un1_M_this_sprites_address_q_cry_9\
        );

    \I__4390\ : InMux
    port map (
            O => \N__21753\,
            I => \un1_M_this_sprites_address_q_cry_10\
        );

    \I__4389\ : InMux
    port map (
            O => \N__21750\,
            I => \un1_M_this_sprites_address_q_cry_11\
        );

    \I__4388\ : InMux
    port map (
            O => \N__21747\,
            I => \un1_M_this_sprites_address_q_cry_12\
        );

    \I__4387\ : InMux
    port map (
            O => \N__21744\,
            I => \N__21741\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__21741\,
            I => \N__21738\
        );

    \I__4385\ : Span4Mux_v
    port map (
            O => \N__21738\,
            I => \N__21735\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__21735\,
            I => \M_this_state_d25\
        );

    \I__4383\ : InMux
    port map (
            O => \N__21732\,
            I => \N__21729\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__21729\,
            I => \N__21724\
        );

    \I__4381\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21721\
        );

    \I__4380\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21718\
        );

    \I__4379\ : Span12Mux_h
    port map (
            O => \N__21724\,
            I => \N__21711\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__21721\,
            I => \N__21711\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__21718\,
            I => \N__21711\
        );

    \I__4376\ : Span12Mux_h
    port map (
            O => \N__21711\,
            I => \N__21707\
        );

    \I__4375\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21704\
        );

    \I__4374\ : Odrv12
    port map (
            O => \N__21707\,
            I => port_rw_in
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__21704\,
            I => port_rw_in
        );

    \I__4372\ : IoInMux
    port map (
            O => \N__21699\,
            I => \N__21696\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__21696\,
            I => \N__21693\
        );

    \I__4370\ : Span4Mux_s3_h
    port map (
            O => \N__21693\,
            I => \N__21690\
        );

    \I__4369\ : Sp12to4
    port map (
            O => \N__21690\,
            I => \N__21686\
        );

    \I__4368\ : InMux
    port map (
            O => \N__21689\,
            I => \N__21683\
        );

    \I__4367\ : Span12Mux_v
    port map (
            O => \N__21686\,
            I => \N__21680\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__21683\,
            I => \N__21675\
        );

    \I__4365\ : Span12Mux_h
    port map (
            O => \N__21680\,
            I => \N__21672\
        );

    \I__4364\ : InMux
    port map (
            O => \N__21679\,
            I => \N__21669\
        );

    \I__4363\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21666\
        );

    \I__4362\ : Span4Mux_h
    port map (
            O => \N__21675\,
            I => \N__21663\
        );

    \I__4361\ : Odrv12
    port map (
            O => \N__21672\,
            I => led_c_1
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__21669\,
            I => led_c_1
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__21666\,
            I => led_c_1
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__21663\,
            I => led_c_1
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__21654\,
            I => \N__21651\
        );

    \I__4356\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21643\
        );

    \I__4355\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21643\
        );

    \I__4354\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21640\
        );

    \I__4353\ : InMux
    port map (
            O => \N__21648\,
            I => \N__21636\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21629\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__21640\,
            I => \N__21629\
        );

    \I__4350\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21626\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__21636\,
            I => \N__21623\
        );

    \I__4348\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21618\
        );

    \I__4347\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21618\
        );

    \I__4346\ : Span4Mux_v
    port map (
            O => \N__21629\,
            I => \N__21613\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__21626\,
            I => \N__21613\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__21623\,
            I => \N_459_0\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__21618\,
            I => \N_459_0\
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__21613\,
            I => \N_459_0\
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__21606\,
            I => \N__21602\
        );

    \I__4340\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21599\
        );

    \I__4339\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21596\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__21599\,
            I => \un1_M_this_state_q_12_0\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__21596\,
            I => \un1_M_this_state_q_12_0\
        );

    \I__4336\ : InMux
    port map (
            O => \N__21591\,
            I => \un1_M_this_sprites_address_q_cry_0\
        );

    \I__4335\ : InMux
    port map (
            O => \N__21588\,
            I => \un1_M_this_sprites_address_q_cry_1\
        );

    \I__4334\ : InMux
    port map (
            O => \N__21585\,
            I => \un1_M_this_sprites_address_q_cry_2\
        );

    \I__4333\ : InMux
    port map (
            O => \N__21582\,
            I => \un1_M_this_sprites_address_q_cry_3\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__21579\,
            I => \N__21573\
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__21578\,
            I => \N__21567\
        );

    \I__4330\ : CascadeMux
    port map (
            O => \N__21577\,
            I => \N__21560\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__21576\,
            I => \N__21557\
        );

    \I__4328\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21554\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__21572\,
            I => \N__21551\
        );

    \I__4326\ : CascadeMux
    port map (
            O => \N__21571\,
            I => \N__21545\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__21570\,
            I => \N__21542\
        );

    \I__4324\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21539\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__21566\,
            I => \N__21534\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__21565\,
            I => \N__21531\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__21564\,
            I => \N__21528\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__21563\,
            I => \N__21525\
        );

    \I__4319\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21522\
        );

    \I__4318\ : InMux
    port map (
            O => \N__21557\,
            I => \N__21519\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__21554\,
            I => \N__21516\
        );

    \I__4316\ : InMux
    port map (
            O => \N__21551\,
            I => \N__21513\
        );

    \I__4315\ : CascadeMux
    port map (
            O => \N__21550\,
            I => \N__21510\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__21549\,
            I => \N__21507\
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__21548\,
            I => \N__21504\
        );

    \I__4312\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21501\
        );

    \I__4311\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21498\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__21539\,
            I => \N__21495\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__21538\,
            I => \N__21492\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__21537\,
            I => \N__21489\
        );

    \I__4307\ : InMux
    port map (
            O => \N__21534\,
            I => \N__21486\
        );

    \I__4306\ : InMux
    port map (
            O => \N__21531\,
            I => \N__21483\
        );

    \I__4305\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21480\
        );

    \I__4304\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21477\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__21522\,
            I => \N__21470\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__21519\,
            I => \N__21470\
        );

    \I__4301\ : Span4Mux_v
    port map (
            O => \N__21516\,
            I => \N__21470\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__21513\,
            I => \N__21467\
        );

    \I__4299\ : InMux
    port map (
            O => \N__21510\,
            I => \N__21464\
        );

    \I__4298\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21461\
        );

    \I__4297\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21458\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__21501\,
            I => \N__21453\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__21498\,
            I => \N__21453\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__21495\,
            I => \N__21450\
        );

    \I__4293\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21447\
        );

    \I__4292\ : InMux
    port map (
            O => \N__21489\,
            I => \N__21444\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__21486\,
            I => \N__21441\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__21483\,
            I => \N__21434\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__21480\,
            I => \N__21434\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__21477\,
            I => \N__21434\
        );

    \I__4287\ : Span4Mux_v
    port map (
            O => \N__21470\,
            I => \N__21429\
        );

    \I__4286\ : Span4Mux_v
    port map (
            O => \N__21467\,
            I => \N__21429\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__21464\,
            I => \N__21424\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__21461\,
            I => \N__21419\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__21458\,
            I => \N__21419\
        );

    \I__4282\ : Span4Mux_v
    port map (
            O => \N__21453\,
            I => \N__21414\
        );

    \I__4281\ : Span4Mux_v
    port map (
            O => \N__21450\,
            I => \N__21414\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__21447\,
            I => \N__21405\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__21444\,
            I => \N__21405\
        );

    \I__4278\ : Span12Mux_s7_h
    port map (
            O => \N__21441\,
            I => \N__21405\
        );

    \I__4277\ : Span12Mux_s9_v
    port map (
            O => \N__21434\,
            I => \N__21405\
        );

    \I__4276\ : Sp12to4
    port map (
            O => \N__21429\,
            I => \N__21402\
        );

    \I__4275\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21398\
        );

    \I__4274\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21395\
        );

    \I__4273\ : Span12Mux_s7_h
    port map (
            O => \N__21424\,
            I => \N__21386\
        );

    \I__4272\ : Span12Mux_s10_v
    port map (
            O => \N__21419\,
            I => \N__21386\
        );

    \I__4271\ : Sp12to4
    port map (
            O => \N__21414\,
            I => \N__21386\
        );

    \I__4270\ : Span12Mux_v
    port map (
            O => \N__21405\,
            I => \N__21386\
        );

    \I__4269\ : Span12Mux_h
    port map (
            O => \N__21402\,
            I => \N__21383\
        );

    \I__4268\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21380\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__21398\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__21395\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__4265\ : Odrv12
    port map (
            O => \N__21386\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__4264\ : Odrv12
    port map (
            O => \N__21383\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__21380\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__4262\ : InMux
    port map (
            O => \N__21369\,
            I => \N__21366\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__21366\,
            I => \un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0\
        );

    \I__4260\ : InMux
    port map (
            O => \N__21363\,
            I => \un1_M_this_sprites_address_q_cry_4\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__21360\,
            I => \N__21356\
        );

    \I__4258\ : CascadeMux
    port map (
            O => \N__21359\,
            I => \N__21353\
        );

    \I__4257\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21348\
        );

    \I__4256\ : InMux
    port map (
            O => \N__21353\,
            I => \N__21345\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__21352\,
            I => \N__21342\
        );

    \I__4254\ : CascadeMux
    port map (
            O => \N__21351\,
            I => \N__21339\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__21348\,
            I => \N__21334\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__21345\,
            I => \N__21331\
        );

    \I__4251\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21328\
        );

    \I__4250\ : InMux
    port map (
            O => \N__21339\,
            I => \N__21325\
        );

    \I__4249\ : CascadeMux
    port map (
            O => \N__21338\,
            I => \N__21322\
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__21337\,
            I => \N__21319\
        );

    \I__4247\ : Span4Mux_v
    port map (
            O => \N__21334\,
            I => \N__21310\
        );

    \I__4246\ : Span4Mux_h
    port map (
            O => \N__21331\,
            I => \N__21310\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21310\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__21325\,
            I => \N__21307\
        );

    \I__4243\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21304\
        );

    \I__4242\ : InMux
    port map (
            O => \N__21319\,
            I => \N__21301\
        );

    \I__4241\ : CascadeMux
    port map (
            O => \N__21318\,
            I => \N__21298\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__21317\,
            I => \N__21293\
        );

    \I__4239\ : Span4Mux_v
    port map (
            O => \N__21310\,
            I => \N__21284\
        );

    \I__4238\ : Span4Mux_h
    port map (
            O => \N__21307\,
            I => \N__21284\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__21304\,
            I => \N__21284\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__21301\,
            I => \N__21281\
        );

    \I__4235\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21278\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__21297\,
            I => \N__21275\
        );

    \I__4233\ : CascadeMux
    port map (
            O => \N__21296\,
            I => \N__21272\
        );

    \I__4232\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21267\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__21292\,
            I => \N__21264\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__21291\,
            I => \N__21261\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__21284\,
            I => \N__21253\
        );

    \I__4228\ : Span4Mux_h
    port map (
            O => \N__21281\,
            I => \N__21253\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__21278\,
            I => \N__21253\
        );

    \I__4226\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21250\
        );

    \I__4225\ : InMux
    port map (
            O => \N__21272\,
            I => \N__21247\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__21271\,
            I => \N__21244\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__21270\,
            I => \N__21241\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__21267\,
            I => \N__21238\
        );

    \I__4221\ : InMux
    port map (
            O => \N__21264\,
            I => \N__21235\
        );

    \I__4220\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21232\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__21260\,
            I => \N__21229\
        );

    \I__4218\ : Span4Mux_v
    port map (
            O => \N__21253\,
            I => \N__21226\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__21250\,
            I => \N__21221\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__21247\,
            I => \N__21221\
        );

    \I__4215\ : InMux
    port map (
            O => \N__21244\,
            I => \N__21218\
        );

    \I__4214\ : InMux
    port map (
            O => \N__21241\,
            I => \N__21215\
        );

    \I__4213\ : Span4Mux_v
    port map (
            O => \N__21238\,
            I => \N__21208\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__21235\,
            I => \N__21208\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21205\
        );

    \I__4210\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21202\
        );

    \I__4209\ : Span4Mux_v
    port map (
            O => \N__21226\,
            I => \N__21193\
        );

    \I__4208\ : Span4Mux_v
    port map (
            O => \N__21221\,
            I => \N__21193\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__21218\,
            I => \N__21193\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21193\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__21214\,
            I => \N__21190\
        );

    \I__4204\ : InMux
    port map (
            O => \N__21213\,
            I => \N__21187\
        );

    \I__4203\ : Span4Mux_v
    port map (
            O => \N__21208\,
            I => \N__21181\
        );

    \I__4202\ : Span4Mux_v
    port map (
            O => \N__21205\,
            I => \N__21181\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__21202\,
            I => \N__21178\
        );

    \I__4200\ : Span4Mux_v
    port map (
            O => \N__21193\,
            I => \N__21175\
        );

    \I__4199\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21172\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__21187\,
            I => \N__21169\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__21186\,
            I => \N__21165\
        );

    \I__4196\ : Sp12to4
    port map (
            O => \N__21181\,
            I => \N__21162\
        );

    \I__4195\ : Span12Mux_h
    port map (
            O => \N__21178\,
            I => \N__21155\
        );

    \I__4194\ : Sp12to4
    port map (
            O => \N__21175\,
            I => \N__21155\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__21172\,
            I => \N__21155\
        );

    \I__4192\ : Span4Mux_h
    port map (
            O => \N__21169\,
            I => \N__21152\
        );

    \I__4191\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21149\
        );

    \I__4190\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21146\
        );

    \I__4189\ : Odrv12
    port map (
            O => \N__21162\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__4188\ : Odrv12
    port map (
            O => \N__21155\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__4187\ : Odrv4
    port map (
            O => \N__21152\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__21149\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__21146\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__4184\ : InMux
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__21132\,
            I => \un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0\
        );

    \I__4182\ : InMux
    port map (
            O => \N__21129\,
            I => \un1_M_this_sprites_address_q_cry_5\
        );

    \I__4181\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21123\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__21123\,
            I => \N__21120\
        );

    \I__4179\ : Span4Mux_h
    port map (
            O => \N__21120\,
            I => \N__21117\
        );

    \I__4178\ : Span4Mux_v
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__21114\,
            I => \N__21111\
        );

    \I__4176\ : Odrv4
    port map (
            O => \N__21111\,
            I => \this_sprites_ram.mem_out_bus6_3\
        );

    \I__4175\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21105\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__21105\,
            I => \N__21102\
        );

    \I__4173\ : Span4Mux_h
    port map (
            O => \N__21102\,
            I => \N__21099\
        );

    \I__4172\ : Span4Mux_v
    port map (
            O => \N__21099\,
            I => \N__21096\
        );

    \I__4171\ : Odrv4
    port map (
            O => \N__21096\,
            I => \this_sprites_ram.mem_out_bus2_3\
        );

    \I__4170\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21090\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__21090\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\
        );

    \I__4168\ : InMux
    port map (
            O => \N__21087\,
            I => \N__21084\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__21084\,
            I => \N__21081\
        );

    \I__4166\ : Span4Mux_h
    port map (
            O => \N__21081\,
            I => \N__21078\
        );

    \I__4165\ : Span4Mux_v
    port map (
            O => \N__21078\,
            I => \N__21075\
        );

    \I__4164\ : Span4Mux_v
    port map (
            O => \N__21075\,
            I => \N__21072\
        );

    \I__4163\ : Span4Mux_h
    port map (
            O => \N__21072\,
            I => \N__21069\
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__21069\,
            I => \this_sprites_ram.mem_out_bus7_3\
        );

    \I__4161\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21063\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__21063\,
            I => \N__21060\
        );

    \I__4159\ : Span4Mux_h
    port map (
            O => \N__21060\,
            I => \N__21057\
        );

    \I__4158\ : Span4Mux_h
    port map (
            O => \N__21057\,
            I => \N__21054\
        );

    \I__4157\ : Span4Mux_h
    port map (
            O => \N__21054\,
            I => \N__21051\
        );

    \I__4156\ : Odrv4
    port map (
            O => \N__21051\,
            I => \this_sprites_ram.mem_out_bus3_3\
        );

    \I__4155\ : InMux
    port map (
            O => \N__21048\,
            I => \N__21045\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__21045\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\
        );

    \I__4153\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21039\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__21039\,
            I => \N__21036\
        );

    \I__4151\ : Span4Mux_h
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__21033\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__4149\ : InMux
    port map (
            O => \N__21030\,
            I => \N__21024\
        );

    \I__4148\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21024\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__21024\,
            I => \N__21018\
        );

    \I__4146\ : InMux
    port map (
            O => \N__21023\,
            I => \N__21015\
        );

    \I__4145\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21010\
        );

    \I__4144\ : InMux
    port map (
            O => \N__21021\,
            I => \N__21010\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__21018\,
            I => \N__21007\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__21015\,
            I => \N__21004\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__21010\,
            I => \N__21001\
        );

    \I__4140\ : Span4Mux_v
    port map (
            O => \N__21007\,
            I => \N__20998\
        );

    \I__4139\ : Span4Mux_v
    port map (
            O => \N__21004\,
            I => \N__20993\
        );

    \I__4138\ : Span4Mux_h
    port map (
            O => \N__21001\,
            I => \N__20993\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__20998\,
            I => \N__20985\
        );

    \I__4136\ : Span4Mux_v
    port map (
            O => \N__20993\,
            I => \N__20982\
        );

    \I__4135\ : InMux
    port map (
            O => \N__20992\,
            I => \N__20973\
        );

    \I__4134\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20973\
        );

    \I__4133\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20973\
        );

    \I__4132\ : InMux
    port map (
            O => \N__20989\,
            I => \N__20973\
        );

    \I__4131\ : InMux
    port map (
            O => \N__20988\,
            I => \N__20970\
        );

    \I__4130\ : Span4Mux_v
    port map (
            O => \N__20985\,
            I => \N__20967\
        );

    \I__4129\ : Span4Mux_v
    port map (
            O => \N__20982\,
            I => \N__20964\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__20973\,
            I => \N__20959\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__20970\,
            I => \N__20959\
        );

    \I__4126\ : IoSpan4Mux
    port map (
            O => \N__20967\,
            I => \N__20956\
        );

    \I__4125\ : Span4Mux_v
    port map (
            O => \N__20964\,
            I => \N__20953\
        );

    \I__4124\ : Span12Mux_v
    port map (
            O => \N__20959\,
            I => \N__20950\
        );

    \I__4123\ : Odrv4
    port map (
            O => \N__20956\,
            I => rst_n_c
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__20953\,
            I => rst_n_c
        );

    \I__4121\ : Odrv12
    port map (
            O => \N__20950\,
            I => rst_n_c
        );

    \I__4120\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20940\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__20940\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__20937\,
            I => \N__20931\
        );

    \I__4117\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20928\
        );

    \I__4116\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20925\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__20934\,
            I => \N__20921\
        );

    \I__4114\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20917\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__20928\,
            I => \N__20914\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__20925\,
            I => \N__20911\
        );

    \I__4111\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20904\
        );

    \I__4110\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20904\
        );

    \I__4109\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20904\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__20917\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__4107\ : Odrv4
    port map (
            O => \N__20914\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__20911\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__20904\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__20895\,
            I => \N__20890\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__20894\,
            I => \N__20887\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__20893\,
            I => \N__20882\
        );

    \I__4101\ : InMux
    port map (
            O => \N__20890\,
            I => \N__20878\
        );

    \I__4100\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20875\
        );

    \I__4099\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20866\
        );

    \I__4098\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20866\
        );

    \I__4097\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20866\
        );

    \I__4096\ : InMux
    port map (
            O => \N__20881\,
            I => \N__20866\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__20878\,
            I => \N__20862\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__20875\,
            I => \N__20859\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20856\
        );

    \I__4092\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20853\
        );

    \I__4091\ : Span4Mux_v
    port map (
            O => \N__20862\,
            I => \N__20850\
        );

    \I__4090\ : Span4Mux_v
    port map (
            O => \N__20859\,
            I => \N__20847\
        );

    \I__4089\ : Span4Mux_v
    port map (
            O => \N__20856\,
            I => \N__20842\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__20853\,
            I => \N__20842\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__20850\,
            I => \N__20837\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__20847\,
            I => \N__20837\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__20842\,
            I => \N__20834\
        );

    \I__4084\ : Span4Mux_v
    port map (
            O => \N__20837\,
            I => \N__20831\
        );

    \I__4083\ : Sp12to4
    port map (
            O => \N__20834\,
            I => \N__20828\
        );

    \I__4082\ : Sp12to4
    port map (
            O => \N__20831\,
            I => \N__20823\
        );

    \I__4081\ : Span12Mux_v
    port map (
            O => \N__20828\,
            I => \N__20823\
        );

    \I__4080\ : Span12Mux_h
    port map (
            O => \N__20823\,
            I => \N__20820\
        );

    \I__4079\ : Odrv12
    port map (
            O => \N__20820\,
            I => port_enb_c
        );

    \I__4078\ : InMux
    port map (
            O => \N__20817\,
            I => \N__20813\
        );

    \I__4077\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20810\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__20813\,
            I => \N__20806\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__20810\,
            I => \N__20803\
        );

    \I__4074\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20796\
        );

    \I__4073\ : Span4Mux_h
    port map (
            O => \N__20806\,
            I => \N__20791\
        );

    \I__4072\ : Span4Mux_v
    port map (
            O => \N__20803\,
            I => \N__20791\
        );

    \I__4071\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20782\
        );

    \I__4070\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20782\
        );

    \I__4069\ : InMux
    port map (
            O => \N__20800\,
            I => \N__20782\
        );

    \I__4068\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20782\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__20796\,
            I => \M_this_delay_clk_out_0\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__20791\,
            I => \M_this_delay_clk_out_0\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__20782\,
            I => \M_this_delay_clk_out_0\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__20775\,
            I => \N_156_0_cascade_\
        );

    \I__4063\ : InMux
    port map (
            O => \N__20772\,
            I => \N__20769\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__20769\,
            I => \N__20766\
        );

    \I__4061\ : Span12Mux_h
    port map (
            O => \N__20766\,
            I => \N__20763\
        );

    \I__4060\ : Odrv12
    port map (
            O => \N__20763\,
            I => \N_35_0\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__20760\,
            I => \N__20757\
        );

    \I__4058\ : InMux
    port map (
            O => \N__20757\,
            I => \N__20754\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__20754\,
            I => \N__20751\
        );

    \I__4056\ : Span4Mux_v
    port map (
            O => \N__20751\,
            I => \N__20748\
        );

    \I__4055\ : Sp12to4
    port map (
            O => \N__20748\,
            I => \N__20745\
        );

    \I__4054\ : Span12Mux_h
    port map (
            O => \N__20745\,
            I => \N__20742\
        );

    \I__4053\ : Odrv12
    port map (
            O => \N__20742\,
            I => \M_this_map_ram_read_data_5\
        );

    \I__4052\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20736\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__20736\,
            I => \N__20733\
        );

    \I__4050\ : Span4Mux_v
    port map (
            O => \N__20733\,
            I => \N__20730\
        );

    \I__4049\ : Sp12to4
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__4048\ : Span12Mux_h
    port map (
            O => \N__20727\,
            I => \N__20724\
        );

    \I__4047\ : Odrv12
    port map (
            O => \N__20724\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__4046\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20718\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__20718\,
            I => \N__20715\
        );

    \I__4044\ : Span4Mux_h
    port map (
            O => \N__20715\,
            I => \N__20712\
        );

    \I__4043\ : Span4Mux_h
    port map (
            O => \N__20712\,
            I => \N__20709\
        );

    \I__4042\ : Span4Mux_h
    port map (
            O => \N__20709\,
            I => \N__20705\
        );

    \I__4041\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20702\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__20705\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__20702\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__4038\ : CascadeMux
    port map (
            O => \N__20697\,
            I => \M_this_ppu_vram_data_3_cascade_\
        );

    \I__4037\ : InMux
    port map (
            O => \N__20694\,
            I => \N__20691\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__4035\ : Span12Mux_v
    port map (
            O => \N__20688\,
            I => \N__20684\
        );

    \I__4034\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20681\
        );

    \I__4033\ : Odrv12
    port map (
            O => \N__20684\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__20681\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__20676\,
            I => \this_ppu.N_156_cascade_\
        );

    \I__4030\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20670\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__20670\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3\
        );

    \I__4028\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20664\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__20664\,
            I => \N__20661\
        );

    \I__4026\ : Span4Mux_h
    port map (
            O => \N__20661\,
            I => \N__20658\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__20658\,
            I => \N__20655\
        );

    \I__4024\ : Span4Mux_h
    port map (
            O => \N__20655\,
            I => \N__20652\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__20652\,
            I => \this_sprites_ram.mem_out_bus5_2\
        );

    \I__4022\ : InMux
    port map (
            O => \N__20649\,
            I => \N__20646\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__20646\,
            I => \N__20643\
        );

    \I__4020\ : Span4Mux_h
    port map (
            O => \N__20643\,
            I => \N__20640\
        );

    \I__4019\ : Span4Mux_h
    port map (
            O => \N__20640\,
            I => \N__20637\
        );

    \I__4018\ : Span4Mux_v
    port map (
            O => \N__20637\,
            I => \N__20634\
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__20634\,
            I => \this_sprites_ram.mem_out_bus1_2\
        );

    \I__4016\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20628\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__20628\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__20625\,
            I => \this_ppu.un1_M_haddress_q_3_c2_cascade_\
        );

    \I__4013\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20613\
        );

    \I__4012\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20613\
        );

    \I__4011\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20613\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__20613\,
            I => \this_ppu.un1_M_haddress_q_3_c5\
        );

    \I__4009\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20604\
        );

    \I__4008\ : InMux
    port map (
            O => \N__20609\,
            I => \N__20601\
        );

    \I__4007\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20597\
        );

    \I__4006\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20594\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__20604\,
            I => \N__20591\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__20601\,
            I => \N__20588\
        );

    \I__4003\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20585\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__20597\,
            I => \N__20580\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__20594\,
            I => \N__20580\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__20591\,
            I => \N__20574\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__20588\,
            I => \N__20574\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__20585\,
            I => \N__20571\
        );

    \I__3997\ : Span4Mux_h
    port map (
            O => \N__20580\,
            I => \N__20568\
        );

    \I__3996\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20565\
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__20574\,
            I => \M_this_state_d55\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__20571\,
            I => \M_this_state_d55\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__20568\,
            I => \M_this_state_d55\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__20565\,
            I => \M_this_state_d55\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__20556\,
            I => \this_vga_signals_M_this_state_q_ns_i_o3_0_7_cascade_\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__20553\,
            I => \N__20548\
        );

    \I__3989\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20545\
        );

    \I__3988\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20542\
        );

    \I__3987\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20539\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__20545\,
            I => \N__20536\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20533\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__20539\,
            I => \N__20530\
        );

    \I__3983\ : Odrv12
    port map (
            O => \N__20536\,
            I => \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__20533\,
            I => \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0\
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__20530\,
            I => \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0\
        );

    \I__3980\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__20520\,
            I => \N__20516\
        );

    \I__3978\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20513\
        );

    \I__3977\ : Span4Mux_v
    port map (
            O => \N__20516\,
            I => \N__20509\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__20513\,
            I => \N__20506\
        );

    \I__3975\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20503\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__20509\,
            I => \this_vga_signals.N_279\
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__20506\,
            I => \this_vga_signals.N_279\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__20503\,
            I => \this_vga_signals.N_279\
        );

    \I__3971\ : CascadeMux
    port map (
            O => \N__20496\,
            I => \N__20493\
        );

    \I__3970\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20489\
        );

    \I__3969\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20484\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__20489\,
            I => \N__20481\
        );

    \I__3967\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20476\
        );

    \I__3966\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20476\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__20484\,
            I => \N__20473\
        );

    \I__3964\ : Span4Mux_h
    port map (
            O => \N__20481\,
            I => \N__20470\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__20476\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__20473\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__20470\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__3960\ : InMux
    port map (
            O => \N__20463\,
            I => \N__20460\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__20460\,
            I => \N__20455\
        );

    \I__3958\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20452\
        );

    \I__3957\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20449\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__20455\,
            I => \N__20446\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20441\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__20449\,
            I => \N__20441\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__20446\,
            I => \N_210\
        );

    \I__3952\ : Odrv12
    port map (
            O => \N__20441\,
            I => \N_210\
        );

    \I__3951\ : InMux
    port map (
            O => \N__20436\,
            I => \N__20430\
        );

    \I__3950\ : InMux
    port map (
            O => \N__20435\,
            I => \N__20426\
        );

    \I__3949\ : InMux
    port map (
            O => \N__20434\,
            I => \N__20421\
        );

    \I__3948\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20421\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__20430\,
            I => \N__20417\
        );

    \I__3946\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20411\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__20426\,
            I => \N__20404\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__20421\,
            I => \N__20404\
        );

    \I__3943\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20401\
        );

    \I__3942\ : Span4Mux_v
    port map (
            O => \N__20417\,
            I => \N__20398\
        );

    \I__3941\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20395\
        );

    \I__3940\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20392\
        );

    \I__3939\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20389\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__20411\,
            I => \N__20386\
        );

    \I__3937\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20383\
        );

    \I__3936\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20380\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__20404\,
            I => \N__20377\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__20401\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3933\ : Odrv4
    port map (
            O => \N__20398\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__20395\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__20392\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__20389\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__20386\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__20383\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__20380\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__20377\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3925\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20355\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__20355\,
            I => \N__20351\
        );

    \I__3923\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20348\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__20351\,
            I => \this_vga_signals.N_166\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__20348\,
            I => \this_vga_signals.N_166\
        );

    \I__3920\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20339\
        );

    \I__3919\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20336\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__20339\,
            I => \N__20330\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__20336\,
            I => \N__20327\
        );

    \I__3916\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20320\
        );

    \I__3915\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20320\
        );

    \I__3914\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20320\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__20330\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__20327\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__20320\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__3910\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20310\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__20310\,
            I => \N__20307\
        );

    \I__3908\ : Span4Mux_h
    port map (
            O => \N__20307\,
            I => \N__20304\
        );

    \I__3907\ : Span4Mux_v
    port map (
            O => \N__20304\,
            I => \N__20301\
        );

    \I__3906\ : Span4Mux_h
    port map (
            O => \N__20301\,
            I => \N__20298\
        );

    \I__3905\ : Span4Mux_h
    port map (
            O => \N__20298\,
            I => \N__20295\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__20295\,
            I => \this_sprites_ram.mem_out_bus5_1\
        );

    \I__3903\ : InMux
    port map (
            O => \N__20292\,
            I => \N__20289\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__20289\,
            I => \N__20286\
        );

    \I__3901\ : Span4Mux_h
    port map (
            O => \N__20286\,
            I => \N__20283\
        );

    \I__3900\ : Span4Mux_v
    port map (
            O => \N__20283\,
            I => \N__20280\
        );

    \I__3899\ : Span4Mux_v
    port map (
            O => \N__20280\,
            I => \N__20277\
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__20277\,
            I => \this_sprites_ram.mem_out_bus1_1\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__20274\,
            I => \N_210_cascade_\
        );

    \I__3896\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20267\
        );

    \I__3895\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20264\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__20267\,
            I => \this_vga_signals.N_159_0\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__20264\,
            I => \this_vga_signals.N_159_0\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__20259\,
            I => \this_vga_signals.N_167_0_cascade_\
        );

    \I__3891\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20253\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__20253\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__20250\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_5_cascade_\
        );

    \I__3888\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20244\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__20244\,
            I => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__20241\,
            I => \N__20238\
        );

    \I__3885\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20235\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__20235\,
            I => \N__20232\
        );

    \I__3883\ : Span4Mux_v
    port map (
            O => \N__20232\,
            I => \N__20229\
        );

    \I__3882\ : Span4Mux_v
    port map (
            O => \N__20229\,
            I => \N__20226\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__20226\,
            I => \this_vga_signals.M_this_sprites_address_q_mZ0Z_6\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__20223\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__20220\,
            I => \N__20217\
        );

    \I__3878\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20214\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__20214\,
            I => \N__20211\
        );

    \I__3876\ : Span4Mux_v
    port map (
            O => \N__20211\,
            I => \N__20208\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__20208\,
            I => \N__20205\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__20205\,
            I => \N__20202\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__20202\,
            I => \N__20199\
        );

    \I__3872\ : Span4Mux_h
    port map (
            O => \N__20199\,
            I => \N__20196\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__20196\,
            I => \M_this_map_ram_read_data_7\
        );

    \I__3870\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__20190\,
            I => \N__20187\
        );

    \I__3868\ : Span4Mux_v
    port map (
            O => \N__20187\,
            I => \N__20184\
        );

    \I__3867\ : Sp12to4
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__3866\ : Span12Mux_h
    port map (
            O => \N__20181\,
            I => \N__20178\
        );

    \I__3865\ : Span12Mux_v
    port map (
            O => \N__20178\,
            I => \N__20175\
        );

    \I__3864\ : Odrv12
    port map (
            O => \N__20175\,
            I => \this_sprites_ram.mem_out_bus7_2\
        );

    \I__3863\ : InMux
    port map (
            O => \N__20172\,
            I => \N__20169\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__20169\,
            I => \N__20166\
        );

    \I__3861\ : Span4Mux_v
    port map (
            O => \N__20166\,
            I => \N__20163\
        );

    \I__3860\ : Span4Mux_h
    port map (
            O => \N__20163\,
            I => \N__20160\
        );

    \I__3859\ : Span4Mux_h
    port map (
            O => \N__20160\,
            I => \N__20157\
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__20157\,
            I => \this_sprites_ram.mem_out_bus3_2\
        );

    \I__3857\ : InMux
    port map (
            O => \N__20154\,
            I => \N__20151\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__20151\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\
        );

    \I__3855\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20141\
        );

    \I__3854\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20141\
        );

    \I__3853\ : InMux
    port map (
            O => \N__20146\,
            I => \N__20138\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__20141\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__20138\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__3850\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20128\
        );

    \I__3849\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20125\
        );

    \I__3848\ : InMux
    port map (
            O => \N__20131\,
            I => \N__20122\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__20128\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__20125\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__20122\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__20115\,
            I => \N__20111\
        );

    \I__3843\ : CascadeMux
    port map (
            O => \N__20114\,
            I => \N__20105\
        );

    \I__3842\ : InMux
    port map (
            O => \N__20111\,
            I => \N__20099\
        );

    \I__3841\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20096\
        );

    \I__3840\ : InMux
    port map (
            O => \N__20109\,
            I => \N__20093\
        );

    \I__3839\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20087\
        );

    \I__3838\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20082\
        );

    \I__3837\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20082\
        );

    \I__3836\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20079\
        );

    \I__3835\ : InMux
    port map (
            O => \N__20102\,
            I => \N__20075\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__20099\,
            I => \N__20072\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__20096\,
            I => \N__20069\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__20093\,
            I => \N__20066\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__20092\,
            I => \N__20063\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__20091\,
            I => \N__20060\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__20090\,
            I => \N__20057\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__20087\,
            I => \N__20054\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__20082\,
            I => \N__20051\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__20079\,
            I => \N__20048\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__20078\,
            I => \N__20045\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__20075\,
            I => \N__20036\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__20072\,
            I => \N__20036\
        );

    \I__3822\ : Span4Mux_v
    port map (
            O => \N__20069\,
            I => \N__20036\
        );

    \I__3821\ : Span4Mux_h
    port map (
            O => \N__20066\,
            I => \N__20036\
        );

    \I__3820\ : InMux
    port map (
            O => \N__20063\,
            I => \N__20031\
        );

    \I__3819\ : InMux
    port map (
            O => \N__20060\,
            I => \N__20031\
        );

    \I__3818\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20028\
        );

    \I__3817\ : Span4Mux_v
    port map (
            O => \N__20054\,
            I => \N__20021\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__20051\,
            I => \N__20021\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__20048\,
            I => \N__20021\
        );

    \I__3814\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20018\
        );

    \I__3813\ : Span4Mux_h
    port map (
            O => \N__20036\,
            I => \N__20015\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__20031\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__20028\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__20021\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__20018\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__20015\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__20004\,
            I => \N__20001\
        );

    \I__3806\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19997\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__20000\,
            I => \N__19994\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__19997\,
            I => \N__19991\
        );

    \I__3803\ : InMux
    port map (
            O => \N__19994\,
            I => \N__19988\
        );

    \I__3802\ : Span4Mux_v
    port map (
            O => \N__19991\,
            I => \N__19983\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__19988\,
            I => \N__19983\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__19983\,
            I => \this_vga_signals.line_clk_1\
        );

    \I__3799\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19977\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__19977\,
            I => \N__19971\
        );

    \I__3797\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19968\
        );

    \I__3796\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19964\
        );

    \I__3795\ : InMux
    port map (
            O => \N__19974\,
            I => \N__19961\
        );

    \I__3794\ : Span4Mux_h
    port map (
            O => \N__19971\,
            I => \N__19958\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__19968\,
            I => \N__19955\
        );

    \I__3792\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19952\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__19964\,
            I => \N__19949\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__19961\,
            I => \N__19945\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__19958\,
            I => \N__19939\
        );

    \I__3788\ : Span4Mux_h
    port map (
            O => \N__19955\,
            I => \N__19939\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19935\
        );

    \I__3786\ : Span4Mux_v
    port map (
            O => \N__19949\,
            I => \N__19932\
        );

    \I__3785\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19929\
        );

    \I__3784\ : Span4Mux_h
    port map (
            O => \N__19945\,
            I => \N__19926\
        );

    \I__3783\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19923\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__19939\,
            I => \N__19920\
        );

    \I__3781\ : InMux
    port map (
            O => \N__19938\,
            I => \N__19917\
        );

    \I__3780\ : Span4Mux_h
    port map (
            O => \N__19935\,
            I => \N__19914\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__19932\,
            I => \N__19909\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__19929\,
            I => \N__19909\
        );

    \I__3777\ : Span4Mux_v
    port map (
            O => \N__19926\,
            I => \N__19906\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__19923\,
            I => \N__19903\
        );

    \I__3775\ : Sp12to4
    port map (
            O => \N__19920\,
            I => \N__19898\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__19917\,
            I => \N__19898\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__19914\,
            I => \N__19895\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__19909\,
            I => \N__19892\
        );

    \I__3771\ : Span4Mux_h
    port map (
            O => \N__19906\,
            I => \N__19889\
        );

    \I__3770\ : Span12Mux_h
    port map (
            O => \N__19903\,
            I => \N__19884\
        );

    \I__3769\ : Span12Mux_h
    port map (
            O => \N__19898\,
            I => \N__19884\
        );

    \I__3768\ : Span4Mux_h
    port map (
            O => \N__19895\,
            I => \N__19879\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__19892\,
            I => \N__19879\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__19889\,
            I => \M_this_sprites_ram_write_data_3\
        );

    \I__3765\ : Odrv12
    port map (
            O => \N__19884\,
            I => \M_this_sprites_ram_write_data_3\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__19879\,
            I => \M_this_sprites_ram_write_data_3\
        );

    \I__3763\ : InMux
    port map (
            O => \N__19872\,
            I => \N__19866\
        );

    \I__3762\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19866\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__19866\,
            I => \N__19863\
        );

    \I__3760\ : Span4Mux_h
    port map (
            O => \N__19863\,
            I => \N__19859\
        );

    \I__3759\ : InMux
    port map (
            O => \N__19862\,
            I => \N__19856\
        );

    \I__3758\ : Odrv4
    port map (
            O => \N__19859\,
            I => \this_vga_signals.N_169_0\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__19856\,
            I => \this_vga_signals.N_169_0\
        );

    \I__3756\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19848\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__19848\,
            I => \N__19845\
        );

    \I__3754\ : Span4Mux_v
    port map (
            O => \N__19845\,
            I => \N__19842\
        );

    \I__3753\ : Sp12to4
    port map (
            O => \N__19842\,
            I => \N__19839\
        );

    \I__3752\ : Span12Mux_h
    port map (
            O => \N__19839\,
            I => \N__19836\
        );

    \I__3751\ : Odrv12
    port map (
            O => \N__19836\,
            I => \this_sprites_ram.mem_out_bus5_0\
        );

    \I__3750\ : InMux
    port map (
            O => \N__19833\,
            I => \N__19830\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__3748\ : Span4Mux_h
    port map (
            O => \N__19827\,
            I => \N__19824\
        );

    \I__3747\ : Span4Mux_h
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__3746\ : Span4Mux_v
    port map (
            O => \N__19821\,
            I => \N__19818\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__19818\,
            I => \this_sprites_ram.mem_out_bus1_0\
        );

    \I__3744\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__19812\,
            I => \N__19809\
        );

    \I__3742\ : Span4Mux_v
    port map (
            O => \N__19809\,
            I => \N__19806\
        );

    \I__3741\ : Span4Mux_v
    port map (
            O => \N__19806\,
            I => \N__19803\
        );

    \I__3740\ : Sp12to4
    port map (
            O => \N__19803\,
            I => \N__19800\
        );

    \I__3739\ : Odrv12
    port map (
            O => \N__19800\,
            I => \this_sprites_ram.mem_out_bus4_0\
        );

    \I__3738\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19794\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__19794\,
            I => \N__19791\
        );

    \I__3736\ : Span4Mux_h
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__19788\,
            I => \N__19785\
        );

    \I__3734\ : Span4Mux_v
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__3733\ : Span4Mux_v
    port map (
            O => \N__19782\,
            I => \N__19779\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__19779\,
            I => \this_sprites_ram.mem_out_bus0_0\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__19776\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_\
        );

    \I__3730\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__19770\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\
        );

    \I__3728\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19764\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__19764\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__19761\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_\
        );

    \I__3725\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__19755\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\
        );

    \I__3723\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19749\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__19749\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__3721\ : InMux
    port map (
            O => \N__19746\,
            I => \N__19743\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__19743\,
            I => \this_reset_cond.M_stage_qZ0Z_3\
        );

    \I__3719\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19737\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__19737\,
            I => \this_reset_cond.M_stage_qZ0Z_4\
        );

    \I__3717\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19731\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__19731\,
            I => \N__19728\
        );

    \I__3715\ : Span4Mux_v
    port map (
            O => \N__19728\,
            I => \N__19725\
        );

    \I__3714\ : Span4Mux_v
    port map (
            O => \N__19725\,
            I => \N__19722\
        );

    \I__3713\ : Sp12to4
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__3712\ : Odrv12
    port map (
            O => \N__19719\,
            I => \this_sprites_ram.mem_out_bus4_2\
        );

    \I__3711\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19713\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__19713\,
            I => \N__19710\
        );

    \I__3709\ : Span4Mux_h
    port map (
            O => \N__19710\,
            I => \N__19707\
        );

    \I__3708\ : Span4Mux_h
    port map (
            O => \N__19707\,
            I => \N__19704\
        );

    \I__3707\ : Span4Mux_v
    port map (
            O => \N__19704\,
            I => \N__19701\
        );

    \I__3706\ : Span4Mux_v
    port map (
            O => \N__19701\,
            I => \N__19698\
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__19698\,
            I => \this_sprites_ram.mem_out_bus0_2\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__19695\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__19692\,
            I => \N__19686\
        );

    \I__3702\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19683\
        );

    \I__3701\ : InMux
    port map (
            O => \N__19690\,
            I => \N__19678\
        );

    \I__3700\ : InMux
    port map (
            O => \N__19689\,
            I => \N__19678\
        );

    \I__3699\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19675\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__19683\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__19678\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__19675\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__3695\ : InMux
    port map (
            O => \N__19668\,
            I => \N__19662\
        );

    \I__3694\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19662\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__19662\,
            I => \N_456_0_1\
        );

    \I__3692\ : InMux
    port map (
            O => \N__19659\,
            I => \N__19656\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__19656\,
            I => \N_500\
        );

    \I__3690\ : InMux
    port map (
            O => \N__19653\,
            I => \N__19648\
        );

    \I__3689\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19644\
        );

    \I__3688\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19637\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__19648\,
            I => \N__19634\
        );

    \I__3686\ : InMux
    port map (
            O => \N__19647\,
            I => \N__19631\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__19644\,
            I => \N__19628\
        );

    \I__3684\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19625\
        );

    \I__3683\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19622\
        );

    \I__3682\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19619\
        );

    \I__3681\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19616\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__19637\,
            I => \N__19613\
        );

    \I__3679\ : Span12Mux_h
    port map (
            O => \N__19634\,
            I => \N__19610\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__19631\,
            I => \N__19607\
        );

    \I__3677\ : Span12Mux_s11_v
    port map (
            O => \N__19628\,
            I => \N__19602\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__19625\,
            I => \N__19602\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__19622\,
            I => \N__19599\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__19619\,
            I => \N__19596\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__19616\,
            I => \N__19593\
        );

    \I__3672\ : Span12Mux_h
    port map (
            O => \N__19613\,
            I => \N__19590\
        );

    \I__3671\ : Span12Mux_v
    port map (
            O => \N__19610\,
            I => \N__19585\
        );

    \I__3670\ : Span12Mux_h
    port map (
            O => \N__19607\,
            I => \N__19585\
        );

    \I__3669\ : Span12Mux_v
    port map (
            O => \N__19602\,
            I => \N__19576\
        );

    \I__3668\ : Span12Mux_s8_v
    port map (
            O => \N__19599\,
            I => \N__19576\
        );

    \I__3667\ : Span12Mux_h
    port map (
            O => \N__19596\,
            I => \N__19576\
        );

    \I__3666\ : Span12Mux_s7_h
    port map (
            O => \N__19593\,
            I => \N__19576\
        );

    \I__3665\ : Odrv12
    port map (
            O => \N__19590\,
            I => \M_this_sprites_ram_write_data_0\
        );

    \I__3664\ : Odrv12
    port map (
            O => \N__19585\,
            I => \M_this_sprites_ram_write_data_0\
        );

    \I__3663\ : Odrv12
    port map (
            O => \N__19576\,
            I => \M_this_sprites_ram_write_data_0\
        );

    \I__3662\ : CascadeMux
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__3661\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19563\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__19563\,
            I => \N__19559\
        );

    \I__3659\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19556\
        );

    \I__3658\ : Span4Mux_v
    port map (
            O => \N__19559\,
            I => \N__19553\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__19556\,
            I => \N__19550\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__19553\,
            I => \M_this_state_d_2_sqmuxa\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__19550\,
            I => \M_this_state_d_2_sqmuxa\
        );

    \I__3654\ : InMux
    port map (
            O => \N__19545\,
            I => \N__19540\
        );

    \I__3653\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19537\
        );

    \I__3652\ : InMux
    port map (
            O => \N__19543\,
            I => \N__19534\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__19540\,
            I => \M_this_substate_qZ0\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__19537\,
            I => \M_this_substate_qZ0\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__19534\,
            I => \M_this_substate_qZ0\
        );

    \I__3648\ : CascadeMux
    port map (
            O => \N__19527\,
            I => \N__19523\
        );

    \I__3647\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19518\
        );

    \I__3646\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19518\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__19518\,
            I => \N__19515\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__19515\,
            I => \this_vga_signals_M_this_state_q_ns_0_a3_0_0_1\
        );

    \I__3643\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19509\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__19509\,
            I => \N__19506\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__19506\,
            I => \N__19503\
        );

    \I__3640\ : Sp12to4
    port map (
            O => \N__19503\,
            I => \N__19500\
        );

    \I__3639\ : Span12Mux_h
    port map (
            O => \N__19500\,
            I => \N__19497\
        );

    \I__3638\ : Span12Mux_v
    port map (
            O => \N__19497\,
            I => \N__19494\
        );

    \I__3637\ : Odrv12
    port map (
            O => \N__19494\,
            I => \this_sprites_ram.mem_out_bus7_0\
        );

    \I__3636\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19488\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__19488\,
            I => \N__19485\
        );

    \I__3634\ : Span4Mux_h
    port map (
            O => \N__19485\,
            I => \N__19482\
        );

    \I__3633\ : Span4Mux_h
    port map (
            O => \N__19482\,
            I => \N__19479\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__19479\,
            I => \this_sprites_ram.mem_out_bus3_0\
        );

    \I__3631\ : InMux
    port map (
            O => \N__19476\,
            I => \N__19473\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__19473\,
            I => \N__19470\
        );

    \I__3629\ : Span4Mux_h
    port map (
            O => \N__19470\,
            I => \N__19467\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__3627\ : Span4Mux_v
    port map (
            O => \N__19464\,
            I => \N__19461\
        );

    \I__3626\ : Span4Mux_h
    port map (
            O => \N__19461\,
            I => \N__19458\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__19458\,
            I => \this_sprites_ram.mem_out_bus6_0\
        );

    \I__3624\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19452\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__19452\,
            I => \N__19449\
        );

    \I__3622\ : Span4Mux_h
    port map (
            O => \N__19449\,
            I => \N__19446\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__19446\,
            I => \N__19443\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__19443\,
            I => \this_sprites_ram.mem_out_bus2_0\
        );

    \I__3619\ : InMux
    port map (
            O => \N__19440\,
            I => \N__19437\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__19437\,
            I => \N__19433\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__19436\,
            I => \N__19430\
        );

    \I__3616\ : Span4Mux_v
    port map (
            O => \N__19433\,
            I => \N__19427\
        );

    \I__3615\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19424\
        );

    \I__3614\ : Span4Mux_h
    port map (
            O => \N__19427\,
            I => \N__19421\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__19424\,
            I => \N__19418\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__19421\,
            I => \this_vga_signals_N_419_i_i_0_a3_1_0\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__19418\,
            I => \this_vga_signals_N_419_i_i_0_a3_1_0\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__19413\,
            I => \N_496_0_cascade_\
        );

    \I__3609\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19406\
        );

    \I__3608\ : InMux
    port map (
            O => \N__19409\,
            I => \N__19403\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__19406\,
            I => \N__19400\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__19403\,
            I => \N__19397\
        );

    \I__3605\ : Span4Mux_h
    port map (
            O => \N__19400\,
            I => \N__19390\
        );

    \I__3604\ : Span4Mux_h
    port map (
            O => \N__19397\,
            I => \N__19390\
        );

    \I__3603\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19385\
        );

    \I__3602\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19385\
        );

    \I__3601\ : Odrv4
    port map (
            O => \N__19390\,
            I => \N_278\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__19385\,
            I => \N_278\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__19380\,
            I => \M_this_state_qsr_0_cascade_\
        );

    \I__3598\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19374\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__19374\,
            I => \N_462_0\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__19371\,
            I => \M_this_state_qsr_2_cascade_\
        );

    \I__3595\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19365\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__19365\,
            I => \N__19362\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__19362\,
            I => \N__19357\
        );

    \I__3592\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19352\
        );

    \I__3591\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19352\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__19357\,
            I => \N_484_0\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__19352\,
            I => \N_484_0\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__19347\,
            I => \this_vga_signals.N_159_0_cascade_\
        );

    \I__3587\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19340\
        );

    \I__3586\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19335\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__19340\,
            I => \N__19332\
        );

    \I__3584\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19329\
        );

    \I__3583\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19326\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__19335\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__3581\ : Odrv4
    port map (
            O => \N__19332\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__19329\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__19326\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__3578\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19314\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__19314\,
            I => \N__19310\
        );

    \I__3576\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19307\
        );

    \I__3575\ : Span4Mux_v
    port map (
            O => \N__19310\,
            I => \N__19302\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__19307\,
            I => \N__19302\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__19302\,
            I => \N_168_0\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__19299\,
            I => \N_168_0_cascade_\
        );

    \I__3571\ : InMux
    port map (
            O => \N__19296\,
            I => \N__19293\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__19293\,
            I => \this_vga_signals.M_this_external_address_d_0_sqmuxa_1Z0Z_2\
        );

    \I__3569\ : CascadeMux
    port map (
            O => \N__19290\,
            I => \N__19285\
        );

    \I__3568\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19278\
        );

    \I__3567\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19278\
        );

    \I__3566\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19273\
        );

    \I__3565\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19273\
        );

    \I__3564\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19270\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__19278\,
            I => \this_ppu.un16_0\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__19273\,
            I => \this_ppu.un16_0\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__19270\,
            I => \this_ppu.un16_0\
        );

    \I__3560\ : InMux
    port map (
            O => \N__19263\,
            I => \N__19260\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__19260\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__19257\,
            I => \this_ppu.un16_0_cascade_\
        );

    \I__3557\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19240\
        );

    \I__3556\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19240\
        );

    \I__3555\ : InMux
    port map (
            O => \N__19252\,
            I => \N__19240\
        );

    \I__3554\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19240\
        );

    \I__3553\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19237\
        );

    \I__3552\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19234\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__19240\,
            I => \this_ppu.N_1157_0\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__19237\,
            I => \this_ppu.N_1157_0\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__19234\,
            I => \this_ppu.N_1157_0\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__19227\,
            I => \N__19224\
        );

    \I__3547\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19221\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__19221\,
            I => \N__19216\
        );

    \I__3545\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19213\
        );

    \I__3544\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19210\
        );

    \I__3543\ : Span4Mux_h
    port map (
            O => \N__19216\,
            I => \N__19207\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__19213\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__19210\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__19207\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__19200\,
            I => \N_459_0_cascade_\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__19197\,
            I => \N_458_0_cascade_\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__19194\,
            I => \this_ppu.N_132_0_cascade_\
        );

    \I__3536\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19186\
        );

    \I__3535\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19181\
        );

    \I__3534\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19181\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__19186\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__19181\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__3531\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19173\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__19173\,
            I => \N__19170\
        );

    \I__3529\ : Span4Mux_h
    port map (
            O => \N__19170\,
            I => \N__19167\
        );

    \I__3528\ : Odrv4
    port map (
            O => \N__19167\,
            I => \this_vga_signals.M_vcounter_d8\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__19164\,
            I => \this_vga_signals.un1_M_hcounter_d7_1_0_cascade_\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__19161\,
            I => \N__19158\
        );

    \I__3525\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19155\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__19155\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\
        );

    \I__3523\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19147\
        );

    \I__3522\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19144\
        );

    \I__3521\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19141\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__19147\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__19144\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__19141\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__3517\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19124\
        );

    \I__3516\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19124\
        );

    \I__3515\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19124\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__19131\,
            I => \N__19120\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19116\
        );

    \I__3512\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19109\
        );

    \I__3511\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19106\
        );

    \I__3510\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19103\
        );

    \I__3509\ : Span4Mux_v
    port map (
            O => \N__19116\,
            I => \N__19099\
        );

    \I__3508\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19090\
        );

    \I__3507\ : InMux
    port map (
            O => \N__19114\,
            I => \N__19090\
        );

    \I__3506\ : InMux
    port map (
            O => \N__19113\,
            I => \N__19090\
        );

    \I__3505\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19090\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__19109\,
            I => \N__19083\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__19106\,
            I => \N__19083\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__19103\,
            I => \N__19083\
        );

    \I__3501\ : InMux
    port map (
            O => \N__19102\,
            I => \N__19080\
        );

    \I__3500\ : Span4Mux_h
    port map (
            O => \N__19099\,
            I => \N__19075\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__19090\,
            I => \N__19075\
        );

    \I__3498\ : Span4Mux_h
    port map (
            O => \N__19083\,
            I => \N__19072\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__19080\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__19075\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__19072\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__3494\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19048\
        );

    \I__3493\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19048\
        );

    \I__3492\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19039\
        );

    \I__3491\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19039\
        );

    \I__3490\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19039\
        );

    \I__3489\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19039\
        );

    \I__3488\ : InMux
    port map (
            O => \N__19059\,
            I => \N__19032\
        );

    \I__3487\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19032\
        );

    \I__3486\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19032\
        );

    \I__3485\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19029\
        );

    \I__3484\ : InMux
    port map (
            O => \N__19055\,
            I => \N__19026\
        );

    \I__3483\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19020\
        );

    \I__3482\ : InMux
    port map (
            O => \N__19053\,
            I => \N__19020\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__19048\,
            I => \N__19013\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__19039\,
            I => \N__19013\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__19032\,
            I => \N__19013\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__19029\,
            I => \N__19010\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__19026\,
            I => \N__19004\
        );

    \I__3476\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19001\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__19020\,
            I => \N__18994\
        );

    \I__3474\ : Span4Mux_v
    port map (
            O => \N__19013\,
            I => \N__18991\
        );

    \I__3473\ : Span12Mux_s1_h
    port map (
            O => \N__19010\,
            I => \N__18988\
        );

    \I__3472\ : CEMux
    port map (
            O => \N__19009\,
            I => \N__18985\
        );

    \I__3471\ : InMux
    port map (
            O => \N__19008\,
            I => \N__18980\
        );

    \I__3470\ : InMux
    port map (
            O => \N__19007\,
            I => \N__18980\
        );

    \I__3469\ : Span4Mux_v
    port map (
            O => \N__19004\,
            I => \N__18975\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__19001\,
            I => \N__18975\
        );

    \I__3467\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18969\
        );

    \I__3466\ : InMux
    port map (
            O => \N__18999\,
            I => \N__18969\
        );

    \I__3465\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18964\
        );

    \I__3464\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18964\
        );

    \I__3463\ : Span4Mux_h
    port map (
            O => \N__18994\,
            I => \N__18961\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__18991\,
            I => \N__18958\
        );

    \I__3461\ : Span12Mux_h
    port map (
            O => \N__18988\,
            I => \N__18955\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__18985\,
            I => \N__18948\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__18980\,
            I => \N__18948\
        );

    \I__3458\ : Span4Mux_h
    port map (
            O => \N__18975\,
            I => \N__18948\
        );

    \I__3457\ : InMux
    port map (
            O => \N__18974\,
            I => \N__18945\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__18969\,
            I => \this_vga_signals.GZ0Z_330\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__18964\,
            I => \this_vga_signals.GZ0Z_330\
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__18961\,
            I => \this_vga_signals.GZ0Z_330\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__18958\,
            I => \this_vga_signals.GZ0Z_330\
        );

    \I__3452\ : Odrv12
    port map (
            O => \N__18955\,
            I => \this_vga_signals.GZ0Z_330\
        );

    \I__3451\ : Odrv4
    port map (
            O => \N__18948\,
            I => \this_vga_signals.GZ0Z_330\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__18945\,
            I => \this_vga_signals.GZ0Z_330\
        );

    \I__3449\ : InMux
    port map (
            O => \N__18930\,
            I => \N__18927\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__18927\,
            I => \this_vga_signals.un1_M_hcounter_d7_1_0\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__18924\,
            I => \this_vga_signals.CO0_cascade_\
        );

    \I__3446\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18914\
        );

    \I__3445\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18914\
        );

    \I__3444\ : InMux
    port map (
            O => \N__18919\,
            I => \N__18911\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__18914\,
            I => \this_ppu.N_1157_0_1\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__18911\,
            I => \this_ppu.N_1157_0_1\
        );

    \I__3441\ : InMux
    port map (
            O => \N__18906\,
            I => \N__18903\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__18903\,
            I => \this_vga_signals.M_this_state_d55Z0Z_9\
        );

    \I__3439\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18897\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__18897\,
            I => \this_vga_signals.M_this_state_d55Z0Z_8\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__18894\,
            I => \this_vga_signals.M_this_state_d55Z0Z_7_cascade_\
        );

    \I__3436\ : InMux
    port map (
            O => \N__18891\,
            I => \N__18888\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__18888\,
            I => \this_vga_signals.M_this_state_d55Z0Z_6\
        );

    \I__3434\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18880\
        );

    \I__3433\ : InMux
    port map (
            O => \N__18884\,
            I => \N__18875\
        );

    \I__3432\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18875\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__18880\,
            I => \N__18872\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__18875\,
            I => \N__18868\
        );

    \I__3429\ : Span4Mux_v
    port map (
            O => \N__18872\,
            I => \N__18865\
        );

    \I__3428\ : InMux
    port map (
            O => \N__18871\,
            I => \N__18862\
        );

    \I__3427\ : Span4Mux_v
    port map (
            O => \N__18868\,
            I => \N__18859\
        );

    \I__3426\ : Sp12to4
    port map (
            O => \N__18865\,
            I => \N__18853\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__18862\,
            I => \N__18853\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__18859\,
            I => \N__18850\
        );

    \I__3423\ : InMux
    port map (
            O => \N__18858\,
            I => \N__18847\
        );

    \I__3422\ : Odrv12
    port map (
            O => \N__18853\,
            I => \M_this_vram_read_data_2\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__18850\,
            I => \M_this_vram_read_data_2\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__18847\,
            I => \M_this_vram_read_data_2\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__18840\,
            I => \N__18836\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__18839\,
            I => \N__18833\
        );

    \I__3417\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18824\
        );

    \I__3416\ : InMux
    port map (
            O => \N__18833\,
            I => \N__18824\
        );

    \I__3415\ : InMux
    port map (
            O => \N__18832\,
            I => \N__18824\
        );

    \I__3414\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18821\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__18824\,
            I => \N__18817\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__18821\,
            I => \N__18814\
        );

    \I__3411\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18810\
        );

    \I__3410\ : Span4Mux_v
    port map (
            O => \N__18817\,
            I => \N__18807\
        );

    \I__3409\ : Span4Mux_v
    port map (
            O => \N__18814\,
            I => \N__18804\
        );

    \I__3408\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18801\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__18810\,
            I => \N__18794\
        );

    \I__3406\ : Sp12to4
    port map (
            O => \N__18807\,
            I => \N__18794\
        );

    \I__3405\ : Sp12to4
    port map (
            O => \N__18804\,
            I => \N__18794\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__18801\,
            I => \M_this_vram_read_data_1\
        );

    \I__3403\ : Odrv12
    port map (
            O => \N__18794\,
            I => \M_this_vram_read_data_1\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__18789\,
            I => \N__18786\
        );

    \I__3401\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18781\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__18785\,
            I => \N__18778\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__18784\,
            I => \N__18774\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__18781\,
            I => \N__18770\
        );

    \I__3397\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18767\
        );

    \I__3396\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18760\
        );

    \I__3395\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18760\
        );

    \I__3394\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18760\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__18770\,
            I => \N__18756\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__18767\,
            I => \N__18751\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__18760\,
            I => \N__18751\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__18759\,
            I => \N__18748\
        );

    \I__3389\ : Span4Mux_h
    port map (
            O => \N__18756\,
            I => \N__18743\
        );

    \I__3388\ : Span4Mux_v
    port map (
            O => \N__18751\,
            I => \N__18743\
        );

    \I__3387\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18740\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__18743\,
            I => \N__18737\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__18740\,
            I => \M_this_vram_read_data_3\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__18737\,
            I => \M_this_vram_read_data_3\
        );

    \I__3383\ : InMux
    port map (
            O => \N__18732\,
            I => \N__18726\
        );

    \I__3382\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18719\
        );

    \I__3381\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18719\
        );

    \I__3380\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18719\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18716\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__18719\,
            I => \N__18712\
        );

    \I__3377\ : Span4Mux_v
    port map (
            O => \N__18716\,
            I => \N__18709\
        );

    \I__3376\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18706\
        );

    \I__3375\ : Span4Mux_h
    port map (
            O => \N__18712\,
            I => \N__18703\
        );

    \I__3374\ : Sp12to4
    port map (
            O => \N__18709\,
            I => \N__18697\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18697\
        );

    \I__3372\ : Span4Mux_h
    port map (
            O => \N__18703\,
            I => \N__18694\
        );

    \I__3371\ : InMux
    port map (
            O => \N__18702\,
            I => \N__18691\
        );

    \I__3370\ : Odrv12
    port map (
            O => \N__18697\,
            I => \M_this_vram_read_data_0\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__18694\,
            I => \M_this_vram_read_data_0\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__18691\,
            I => \M_this_vram_read_data_0\
        );

    \I__3367\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18681\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__18681\,
            I => \N__18678\
        );

    \I__3365\ : Span4Mux_h
    port map (
            O => \N__18678\,
            I => \N__18675\
        );

    \I__3364\ : Odrv4
    port map (
            O => \N__18675\,
            I => \this_vga_ramdac.m16\
        );

    \I__3363\ : InMux
    port map (
            O => \N__18672\,
            I => \N__18669\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__18669\,
            I => \this_reset_cond.M_stage_qZ0Z_5\
        );

    \I__3361\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18663\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__18663\,
            I => \N__18660\
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__18660\,
            I => \this_reset_cond.M_stage_qZ0Z_8\
        );

    \I__3358\ : InMux
    port map (
            O => \N__18657\,
            I => \N__18654\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__18654\,
            I => \this_reset_cond.M_stage_qZ0Z_6\
        );

    \I__3356\ : InMux
    port map (
            O => \N__18651\,
            I => \N__18648\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__18648\,
            I => \this_reset_cond.M_stage_qZ0Z_7\
        );

    \I__3354\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18641\
        );

    \I__3353\ : InMux
    port map (
            O => \N__18644\,
            I => \N__18638\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__18641\,
            I => \this_ppu.M_count_qZ0Z_7\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__18638\,
            I => \this_ppu.M_count_qZ0Z_7\
        );

    \I__3350\ : InMux
    port map (
            O => \N__18633\,
            I => \N__18630\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__18630\,
            I => \this_ppu.M_count_d_1_sqmuxa_1_i_a2_3\
        );

    \I__3348\ : InMux
    port map (
            O => \N__18627\,
            I => \N__18624\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__18624\,
            I => \N__18621\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__18621\,
            I => \M_this_state_qc_3_1\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__18618\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_4_cascade_\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__18615\,
            I => \N__18612\
        );

    \I__3343\ : InMux
    port map (
            O => \N__18612\,
            I => \N__18606\
        );

    \I__3342\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18599\
        );

    \I__3341\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18599\
        );

    \I__3340\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18599\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18596\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__18599\,
            I => \N__18593\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__18596\,
            I => \N_465_0\
        );

    \I__3336\ : Odrv12
    port map (
            O => \N__18593\,
            I => \N_465_0\
        );

    \I__3335\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18580\
        );

    \I__3334\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18580\
        );

    \I__3333\ : InMux
    port map (
            O => \N__18586\,
            I => \N__18576\
        );

    \I__3332\ : InMux
    port map (
            O => \N__18585\,
            I => \N__18573\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__18580\,
            I => \N__18570\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__18579\,
            I => \N__18561\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__18576\,
            I => \N__18555\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18552\
        );

    \I__3327\ : Span4Mux_h
    port map (
            O => \N__18570\,
            I => \N__18549\
        );

    \I__3326\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18546\
        );

    \I__3325\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18539\
        );

    \I__3324\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18539\
        );

    \I__3323\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18539\
        );

    \I__3322\ : InMux
    port map (
            O => \N__18565\,
            I => \N__18534\
        );

    \I__3321\ : InMux
    port map (
            O => \N__18564\,
            I => \N__18534\
        );

    \I__3320\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18525\
        );

    \I__3319\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18525\
        );

    \I__3318\ : InMux
    port map (
            O => \N__18559\,
            I => \N__18525\
        );

    \I__3317\ : InMux
    port map (
            O => \N__18558\,
            I => \N__18525\
        );

    \I__3316\ : Odrv12
    port map (
            O => \N__18555\,
            I => \N_610_0_i\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__18552\,
            I => \N_610_0_i\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__18549\,
            I => \N_610_0_i\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__18546\,
            I => \N_610_0_i\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__18539\,
            I => \N_610_0_i\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__18534\,
            I => \N_610_0_i\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__18525\,
            I => \N_610_0_i\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__18510\,
            I => \N__18507\
        );

    \I__3308\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18504\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__18504\,
            I => \N__18501\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__18501\,
            I => \M_this_data_count_q_cry_0_THRU_CO\
        );

    \I__3305\ : CEMux
    port map (
            O => \N__18498\,
            I => \N__18495\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__18495\,
            I => \N__18492\
        );

    \I__3303\ : Span4Mux_v
    port map (
            O => \N__18492\,
            I => \N__18488\
        );

    \I__3302\ : CEMux
    port map (
            O => \N__18491\,
            I => \N__18485\
        );

    \I__3301\ : Span4Mux_v
    port map (
            O => \N__18488\,
            I => \N__18478\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__18485\,
            I => \N__18478\
        );

    \I__3299\ : CEMux
    port map (
            O => \N__18484\,
            I => \N__18473\
        );

    \I__3298\ : CEMux
    port map (
            O => \N__18483\,
            I => \N__18470\
        );

    \I__3297\ : Span4Mux_v
    port map (
            O => \N__18478\,
            I => \N__18467\
        );

    \I__3296\ : CEMux
    port map (
            O => \N__18477\,
            I => \N__18464\
        );

    \I__3295\ : CEMux
    port map (
            O => \N__18476\,
            I => \N__18461\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__18473\,
            I => \M_this_data_count_qe_0_i\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__18470\,
            I => \M_this_data_count_qe_0_i\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__18467\,
            I => \M_this_data_count_qe_0_i\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__18464\,
            I => \M_this_data_count_qe_0_i\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__18461\,
            I => \M_this_data_count_qe_0_i\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__18450\,
            I => \N__18446\
        );

    \I__3288\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18442\
        );

    \I__3287\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18439\
        );

    \I__3286\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18436\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__18442\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__18439\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__18436\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3282\ : InMux
    port map (
            O => \N__18429\,
            I => \N__18424\
        );

    \I__3281\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18421\
        );

    \I__3280\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18418\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__18424\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__18421\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__18418\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__18411\,
            I => \N__18408\
        );

    \I__3275\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18404\
        );

    \I__3274\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18400\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__18404\,
            I => \N__18397\
        );

    \I__3272\ : InMux
    port map (
            O => \N__18403\,
            I => \N__18394\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__18400\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__18397\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__18394\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3268\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18383\
        );

    \I__3267\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18380\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__18383\,
            I => \N__18377\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__18380\,
            I => \N__18374\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__18377\,
            I => \N__18371\
        );

    \I__3263\ : Odrv4
    port map (
            O => \N__18374\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__18371\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3261\ : InMux
    port map (
            O => \N__18366\,
            I => \N__18361\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__18365\,
            I => \N__18358\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__18364\,
            I => \N__18355\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__18361\,
            I => \N__18352\
        );

    \I__3257\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18349\
        );

    \I__3256\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18346\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__18352\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__18349\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__18346\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3252\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18335\
        );

    \I__3251\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18331\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__18335\,
            I => \N__18328\
        );

    \I__3249\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18325\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__18331\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__18328\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__18325\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3245\ : CascadeMux
    port map (
            O => \N__18318\,
            I => \this_vga_signals.N_322_cascade_\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__18315\,
            I => \N__18312\
        );

    \I__3243\ : InMux
    port map (
            O => \N__18312\,
            I => \N__18309\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__18309\,
            I => \this_vga_signals_M_this_state_q_ns_i_o3_0_10\
        );

    \I__3241\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18299\
        );

    \I__3240\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18294\
        );

    \I__3239\ : InMux
    port map (
            O => \N__18304\,
            I => \N__18294\
        );

    \I__3238\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18289\
        );

    \I__3237\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18289\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__18299\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__18294\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__18289\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__3233\ : InMux
    port map (
            O => \N__18282\,
            I => \N__18277\
        );

    \I__3232\ : InMux
    port map (
            O => \N__18281\,
            I => \N__18274\
        );

    \I__3231\ : InMux
    port map (
            O => \N__18280\,
            I => \N__18271\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__18277\,
            I => \N__18268\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__18274\,
            I => \N_212\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__18271\,
            I => \N_212\
        );

    \I__3227\ : Odrv12
    port map (
            O => \N__18268\,
            I => \N_212\
        );

    \I__3226\ : CEMux
    port map (
            O => \N__18261\,
            I => \N__18257\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__18260\,
            I => \N__18252\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__18257\,
            I => \N__18245\
        );

    \I__3223\ : InMux
    port map (
            O => \N__18256\,
            I => \N__18242\
        );

    \I__3222\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18234\
        );

    \I__3221\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18231\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__18251\,
            I => \N__18228\
        );

    \I__3219\ : CEMux
    port map (
            O => \N__18250\,
            I => \N__18225\
        );

    \I__3218\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18220\
        );

    \I__3217\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18220\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__18245\,
            I => \N__18217\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__18242\,
            I => \N__18214\
        );

    \I__3214\ : InMux
    port map (
            O => \N__18241\,
            I => \N__18209\
        );

    \I__3213\ : InMux
    port map (
            O => \N__18240\,
            I => \N__18209\
        );

    \I__3212\ : InMux
    port map (
            O => \N__18239\,
            I => \N__18206\
        );

    \I__3211\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18201\
        );

    \I__3210\ : InMux
    port map (
            O => \N__18237\,
            I => \N__18201\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__18234\,
            I => \N__18196\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__18231\,
            I => \N__18196\
        );

    \I__3207\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18193\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__18225\,
            I => \N__18188\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__18220\,
            I => \N__18188\
        );

    \I__3204\ : Span4Mux_v
    port map (
            O => \N__18217\,
            I => \N__18185\
        );

    \I__3203\ : Span4Mux_h
    port map (
            O => \N__18214\,
            I => \N__18178\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18178\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__18206\,
            I => \N__18178\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__18201\,
            I => \N__18175\
        );

    \I__3199\ : Span4Mux_h
    port map (
            O => \N__18196\,
            I => \N__18172\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__18193\,
            I => \N__18169\
        );

    \I__3197\ : Span12Mux_h
    port map (
            O => \N__18188\,
            I => \N__18166\
        );

    \I__3196\ : Span4Mux_h
    port map (
            O => \N__18185\,
            I => \N__18161\
        );

    \I__3195\ : Span4Mux_v
    port map (
            O => \N__18178\,
            I => \N__18161\
        );

    \I__3194\ : Span4Mux_v
    port map (
            O => \N__18175\,
            I => \N__18156\
        );

    \I__3193\ : Span4Mux_h
    port map (
            O => \N__18172\,
            I => \N__18156\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__18169\,
            I => \N_160_0\
        );

    \I__3191\ : Odrv12
    port map (
            O => \N__18166\,
            I => \N_160_0\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__18161\,
            I => \N_160_0\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__18156\,
            I => \N_160_0\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__18147\,
            I => \N__18144\
        );

    \I__3187\ : InMux
    port map (
            O => \N__18144\,
            I => \N__18141\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__18141\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__18138\,
            I => \N__18134\
        );

    \I__3184\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18130\
        );

    \I__3183\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18125\
        );

    \I__3182\ : InMux
    port map (
            O => \N__18133\,
            I => \N__18125\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__18130\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__18125\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__18120\,
            I => \N__18117\
        );

    \I__3178\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18112\
        );

    \I__3177\ : InMux
    port map (
            O => \N__18116\,
            I => \N__18107\
        );

    \I__3176\ : InMux
    port map (
            O => \N__18115\,
            I => \N__18107\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__18112\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__18107\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__18102\,
            I => \N__18099\
        );

    \I__3172\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18094\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__18098\,
            I => \N__18091\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__18097\,
            I => \N__18088\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__18094\,
            I => \N__18085\
        );

    \I__3168\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18080\
        );

    \I__3167\ : InMux
    port map (
            O => \N__18088\,
            I => \N__18080\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__18085\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__18080\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__18075\,
            I => \N__18072\
        );

    \I__3163\ : InMux
    port map (
            O => \N__18072\,
            I => \N__18067\
        );

    \I__3162\ : InMux
    port map (
            O => \N__18071\,
            I => \N__18062\
        );

    \I__3161\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18062\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__18067\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__18062\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__3158\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18054\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__18054\,
            I => \N__18051\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__18051\,
            I => \this_ppu.M_count_d_1_sqmuxa_1_i_a2_4\
        );

    \I__3155\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18045\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__18045\,
            I => \N__18042\
        );

    \I__3153\ : Span4Mux_h
    port map (
            O => \N__18042\,
            I => \N__18039\
        );

    \I__3152\ : Odrv4
    port map (
            O => \N__18039\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__3151\ : CascadeMux
    port map (
            O => \N__18036\,
            I => \this_vga_signals.un20_i_a2_sxZ0Z_3_cascade_\
        );

    \I__3150\ : InMux
    port map (
            O => \N__18033\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1\
        );

    \I__3149\ : InMux
    port map (
            O => \N__18030\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1\
        );

    \I__3148\ : InMux
    port map (
            O => \N__18027\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1\
        );

    \I__3147\ : InMux
    port map (
            O => \N__18024\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1\
        );

    \I__3146\ : SRMux
    port map (
            O => \N__18021\,
            I => \N__18016\
        );

    \I__3145\ : SRMux
    port map (
            O => \N__18020\,
            I => \N__18013\
        );

    \I__3144\ : SRMux
    port map (
            O => \N__18019\,
            I => \N__18007\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__18016\,
            I => \N__18001\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__18013\,
            I => \N__18001\
        );

    \I__3141\ : SRMux
    port map (
            O => \N__18012\,
            I => \N__17998\
        );

    \I__3140\ : IoInMux
    port map (
            O => \N__18011\,
            I => \N__17993\
        );

    \I__3139\ : SRMux
    port map (
            O => \N__18010\,
            I => \N__17986\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__18007\,
            I => \N__17983\
        );

    \I__3137\ : SRMux
    port map (
            O => \N__18006\,
            I => \N__17980\
        );

    \I__3136\ : Span4Mux_v
    port map (
            O => \N__18001\,
            I => \N__17975\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__17998\,
            I => \N__17975\
        );

    \I__3134\ : SRMux
    port map (
            O => \N__17997\,
            I => \N__17972\
        );

    \I__3133\ : SRMux
    port map (
            O => \N__17996\,
            I => \N__17969\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__17993\,
            I => \N__17965\
        );

    \I__3131\ : SRMux
    port map (
            O => \N__17992\,
            I => \N__17960\
        );

    \I__3130\ : SRMux
    port map (
            O => \N__17991\,
            I => \N__17953\
        );

    \I__3129\ : IoInMux
    port map (
            O => \N__17990\,
            I => \N__17949\
        );

    \I__3128\ : SRMux
    port map (
            O => \N__17989\,
            I => \N__17944\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__17986\,
            I => \N__17935\
        );

    \I__3126\ : Span4Mux_h
    port map (
            O => \N__17983\,
            I => \N__17935\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__17980\,
            I => \N__17935\
        );

    \I__3124\ : Span4Mux_h
    port map (
            O => \N__17975\,
            I => \N__17927\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__17972\,
            I => \N__17927\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__17969\,
            I => \N__17927\
        );

    \I__3121\ : SRMux
    port map (
            O => \N__17968\,
            I => \N__17924\
        );

    \I__3120\ : IoSpan4Mux
    port map (
            O => \N__17965\,
            I => \N__17919\
        );

    \I__3119\ : SRMux
    port map (
            O => \N__17964\,
            I => \N__17916\
        );

    \I__3118\ : SRMux
    port map (
            O => \N__17963\,
            I => \N__17913\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__17960\,
            I => \N__17910\
        );

    \I__3116\ : SRMux
    port map (
            O => \N__17959\,
            I => \N__17907\
        );

    \I__3115\ : SRMux
    port map (
            O => \N__17958\,
            I => \N__17902\
        );

    \I__3114\ : SRMux
    port map (
            O => \N__17957\,
            I => \N__17899\
        );

    \I__3113\ : SRMux
    port map (
            O => \N__17956\,
            I => \N__17891\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__17953\,
            I => \N__17888\
        );

    \I__3111\ : SRMux
    port map (
            O => \N__17952\,
            I => \N__17885\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__17949\,
            I => \N__17881\
        );

    \I__3109\ : SRMux
    port map (
            O => \N__17948\,
            I => \N__17878\
        );

    \I__3108\ : SRMux
    port map (
            O => \N__17947\,
            I => \N__17875\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__17944\,
            I => \N__17872\
        );

    \I__3106\ : SRMux
    port map (
            O => \N__17943\,
            I => \N__17869\
        );

    \I__3105\ : SRMux
    port map (
            O => \N__17942\,
            I => \N__17866\
        );

    \I__3104\ : Span4Mux_v
    port map (
            O => \N__17935\,
            I => \N__17861\
        );

    \I__3103\ : SRMux
    port map (
            O => \N__17934\,
            I => \N__17858\
        );

    \I__3102\ : Span4Mux_v
    port map (
            O => \N__17927\,
            I => \N__17853\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__17924\,
            I => \N__17853\
        );

    \I__3100\ : SRMux
    port map (
            O => \N__17923\,
            I => \N__17850\
        );

    \I__3099\ : SRMux
    port map (
            O => \N__17922\,
            I => \N__17846\
        );

    \I__3098\ : Span4Mux_s3_h
    port map (
            O => \N__17919\,
            I => \N__17843\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__17916\,
            I => \N__17838\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__17913\,
            I => \N__17838\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__17910\,
            I => \N__17833\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__17907\,
            I => \N__17833\
        );

    \I__3093\ : SRMux
    port map (
            O => \N__17906\,
            I => \N__17830\
        );

    \I__3092\ : SRMux
    port map (
            O => \N__17905\,
            I => \N__17827\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__17902\,
            I => \N__17824\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__17899\,
            I => \N__17821\
        );

    \I__3089\ : SRMux
    port map (
            O => \N__17898\,
            I => \N__17818\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__17897\,
            I => \N__17814\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__17896\,
            I => \N__17811\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__17895\,
            I => \N__17807\
        );

    \I__3085\ : SRMux
    port map (
            O => \N__17894\,
            I => \N__17800\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__17891\,
            I => \N__17793\
        );

    \I__3083\ : Span4Mux_h
    port map (
            O => \N__17888\,
            I => \N__17793\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__17885\,
            I => \N__17793\
        );

    \I__3081\ : SRMux
    port map (
            O => \N__17884\,
            I => \N__17790\
        );

    \I__3080\ : IoSpan4Mux
    port map (
            O => \N__17881\,
            I => \N__17787\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__17878\,
            I => \N__17782\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__17875\,
            I => \N__17782\
        );

    \I__3077\ : Span4Mux_v
    port map (
            O => \N__17872\,
            I => \N__17775\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__17869\,
            I => \N__17775\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__17866\,
            I => \N__17775\
        );

    \I__3074\ : SRMux
    port map (
            O => \N__17865\,
            I => \N__17772\
        );

    \I__3073\ : SRMux
    port map (
            O => \N__17864\,
            I => \N__17769\
        );

    \I__3072\ : Span4Mux_h
    port map (
            O => \N__17861\,
            I => \N__17756\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__17858\,
            I => \N__17756\
        );

    \I__3070\ : Span4Mux_v
    port map (
            O => \N__17853\,
            I => \N__17756\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__17850\,
            I => \N__17756\
        );

    \I__3068\ : SRMux
    port map (
            O => \N__17849\,
            I => \N__17753\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__17846\,
            I => \N__17749\
        );

    \I__3066\ : Span4Mux_h
    port map (
            O => \N__17843\,
            I => \N__17740\
        );

    \I__3065\ : Span4Mux_v
    port map (
            O => \N__17838\,
            I => \N__17740\
        );

    \I__3064\ : Span4Mux_v
    port map (
            O => \N__17833\,
            I => \N__17740\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__17830\,
            I => \N__17740\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__17827\,
            I => \N__17735\
        );

    \I__3061\ : Span4Mux_h
    port map (
            O => \N__17824\,
            I => \N__17732\
        );

    \I__3060\ : Span4Mux_h
    port map (
            O => \N__17821\,
            I => \N__17729\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__17818\,
            I => \N__17726\
        );

    \I__3058\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17715\
        );

    \I__3057\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17715\
        );

    \I__3056\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17715\
        );

    \I__3055\ : InMux
    port map (
            O => \N__17810\,
            I => \N__17715\
        );

    \I__3054\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17715\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__17806\,
            I => \N__17710\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__17805\,
            I => \N__17706\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__17804\,
            I => \N__17702\
        );

    \I__3050\ : SRMux
    port map (
            O => \N__17803\,
            I => \N__17699\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__17800\,
            I => \N__17692\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__17793\,
            I => \N__17692\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__17790\,
            I => \N__17692\
        );

    \I__3046\ : Span4Mux_s0_h
    port map (
            O => \N__17787\,
            I => \N__17689\
        );

    \I__3045\ : Span4Mux_v
    port map (
            O => \N__17782\,
            I => \N__17680\
        );

    \I__3044\ : Span4Mux_v
    port map (
            O => \N__17775\,
            I => \N__17680\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__17772\,
            I => \N__17680\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__17769\,
            I => \N__17680\
        );

    \I__3041\ : SRMux
    port map (
            O => \N__17768\,
            I => \N__17677\
        );

    \I__3040\ : SRMux
    port map (
            O => \N__17767\,
            I => \N__17674\
        );

    \I__3039\ : SRMux
    port map (
            O => \N__17766\,
            I => \N__17671\
        );

    \I__3038\ : SRMux
    port map (
            O => \N__17765\,
            I => \N__17668\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__17756\,
            I => \N__17665\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__17753\,
            I => \N__17662\
        );

    \I__3035\ : SRMux
    port map (
            O => \N__17752\,
            I => \N__17659\
        );

    \I__3034\ : Span4Mux_v
    port map (
            O => \N__17749\,
            I => \N__17654\
        );

    \I__3033\ : Span4Mux_v
    port map (
            O => \N__17740\,
            I => \N__17654\
        );

    \I__3032\ : SRMux
    port map (
            O => \N__17739\,
            I => \N__17651\
        );

    \I__3031\ : SRMux
    port map (
            O => \N__17738\,
            I => \N__17648\
        );

    \I__3030\ : Span4Mux_h
    port map (
            O => \N__17735\,
            I => \N__17645\
        );

    \I__3029\ : Span4Mux_h
    port map (
            O => \N__17732\,
            I => \N__17642\
        );

    \I__3028\ : Span4Mux_v
    port map (
            O => \N__17729\,
            I => \N__17639\
        );

    \I__3027\ : Span4Mux_h
    port map (
            O => \N__17726\,
            I => \N__17636\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__17715\,
            I => \N__17633\
        );

    \I__3025\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17618\
        );

    \I__3024\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17618\
        );

    \I__3023\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17618\
        );

    \I__3022\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17618\
        );

    \I__3021\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17618\
        );

    \I__3020\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17618\
        );

    \I__3019\ : InMux
    port map (
            O => \N__17702\,
            I => \N__17618\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__17699\,
            I => \N__17615\
        );

    \I__3017\ : Span4Mux_v
    port map (
            O => \N__17692\,
            I => \N__17612\
        );

    \I__3016\ : Span4Mux_h
    port map (
            O => \N__17689\,
            I => \N__17605\
        );

    \I__3015\ : Span4Mux_v
    port map (
            O => \N__17680\,
            I => \N__17605\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__17677\,
            I => \N__17605\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__17674\,
            I => \N__17595\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__17671\,
            I => \N__17595\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__17668\,
            I => \N__17595\
        );

    \I__3010\ : Sp12to4
    port map (
            O => \N__17665\,
            I => \N__17592\
        );

    \I__3009\ : Span12Mux_s6_v
    port map (
            O => \N__17662\,
            I => \N__17581\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__17659\,
            I => \N__17581\
        );

    \I__3007\ : Sp12to4
    port map (
            O => \N__17654\,
            I => \N__17581\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__17651\,
            I => \N__17581\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__17648\,
            I => \N__17581\
        );

    \I__3004\ : Span4Mux_h
    port map (
            O => \N__17645\,
            I => \N__17578\
        );

    \I__3003\ : Span4Mux_v
    port map (
            O => \N__17642\,
            I => \N__17571\
        );

    \I__3002\ : Span4Mux_h
    port map (
            O => \N__17639\,
            I => \N__17571\
        );

    \I__3001\ : Span4Mux_h
    port map (
            O => \N__17636\,
            I => \N__17571\
        );

    \I__3000\ : Span4Mux_v
    port map (
            O => \N__17633\,
            I => \N__17566\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__17618\,
            I => \N__17566\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__17615\,
            I => \N__17559\
        );

    \I__2997\ : Span4Mux_h
    port map (
            O => \N__17612\,
            I => \N__17559\
        );

    \I__2996\ : Span4Mux_h
    port map (
            O => \N__17605\,
            I => \N__17559\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__17604\,
            I => \N__17555\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__17603\,
            I => \N__17551\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__17602\,
            I => \N__17547\
        );

    \I__2992\ : Span12Mux_v
    port map (
            O => \N__17595\,
            I => \N__17540\
        );

    \I__2991\ : Span12Mux_s7_h
    port map (
            O => \N__17592\,
            I => \N__17540\
        );

    \I__2990\ : Span12Mux_v
    port map (
            O => \N__17581\,
            I => \N__17540\
        );

    \I__2989\ : Span4Mux_h
    port map (
            O => \N__17578\,
            I => \N__17537\
        );

    \I__2988\ : Span4Mux_h
    port map (
            O => \N__17571\,
            I => \N__17534\
        );

    \I__2987\ : Span4Mux_v
    port map (
            O => \N__17566\,
            I => \N__17531\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__17559\,
            I => \N__17528\
        );

    \I__2985\ : InMux
    port map (
            O => \N__17558\,
            I => \N__17515\
        );

    \I__2984\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17515\
        );

    \I__2983\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17515\
        );

    \I__2982\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17515\
        );

    \I__2981\ : InMux
    port map (
            O => \N__17550\,
            I => \N__17515\
        );

    \I__2980\ : InMux
    port map (
            O => \N__17547\,
            I => \N__17515\
        );

    \I__2979\ : Odrv12
    port map (
            O => \N__17540\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2978\ : Odrv4
    port map (
            O => \N__17537\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__17534\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__17531\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2975\ : Odrv4
    port map (
            O => \N__17528\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__17515\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2973\ : InMux
    port map (
            O => \N__17502\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1\
        );

    \I__2972\ : InMux
    port map (
            O => \N__17499\,
            I => \this_ppu.un1_M_count_q_1_cry_6_s1\
        );

    \I__2971\ : InMux
    port map (
            O => \N__17496\,
            I => \N__17493\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__17493\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_7\
        );

    \I__2969\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17487\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__17487\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\
        );

    \I__2967\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17481\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__17481\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\
        );

    \I__2965\ : InMux
    port map (
            O => \N__17478\,
            I => \N__17475\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__17475\,
            I => \N__17472\
        );

    \I__2963\ : Odrv12
    port map (
            O => \N__17472\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__17469\,
            I => \N__17466\
        );

    \I__2961\ : InMux
    port map (
            O => \N__17466\,
            I => \N__17463\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__17463\,
            I => \M_this_data_count_q_cry_1_THRU_CO\
        );

    \I__2959\ : InMux
    port map (
            O => \N__17460\,
            I => \N__17457\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__17457\,
            I => \M_this_data_count_q_cry_8_THRU_CO\
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__17454\,
            I => \N__17450\
        );

    \I__2956\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17446\
        );

    \I__2955\ : InMux
    port map (
            O => \N__17450\,
            I => \N__17443\
        );

    \I__2954\ : InMux
    port map (
            O => \N__17449\,
            I => \N__17440\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__17446\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__17443\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__17440\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__2950\ : InMux
    port map (
            O => \N__17433\,
            I => \N__17430\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__17430\,
            I => \N__17427\
        );

    \I__2948\ : Span4Mux_v
    port map (
            O => \N__17427\,
            I => \N__17424\
        );

    \I__2947\ : Span4Mux_v
    port map (
            O => \N__17424\,
            I => \N__17421\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__17421\,
            I => \N__17418\
        );

    \I__2945\ : Span4Mux_h
    port map (
            O => \N__17418\,
            I => \N__17415\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__17415\,
            I => \M_this_map_ram_read_data_1\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__17412\,
            I => \N__17408\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__17411\,
            I => \N__17402\
        );

    \I__2941\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17396\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__17407\,
            I => \N__17393\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__17406\,
            I => \N__17388\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__17405\,
            I => \N__17385\
        );

    \I__2937\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17381\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__17401\,
            I => \N__17377\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__17400\,
            I => \N__17374\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__17399\,
            I => \N__17371\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__17396\,
            I => \N__17368\
        );

    \I__2932\ : InMux
    port map (
            O => \N__17393\,
            I => \N__17365\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__17392\,
            I => \N__17362\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__17391\,
            I => \N__17359\
        );

    \I__2929\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17355\
        );

    \I__2928\ : InMux
    port map (
            O => \N__17385\,
            I => \N__17352\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__17384\,
            I => \N__17349\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__17381\,
            I => \N__17344\
        );

    \I__2925\ : CascadeMux
    port map (
            O => \N__17380\,
            I => \N__17341\
        );

    \I__2924\ : InMux
    port map (
            O => \N__17377\,
            I => \N__17338\
        );

    \I__2923\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17335\
        );

    \I__2922\ : InMux
    port map (
            O => \N__17371\,
            I => \N__17332\
        );

    \I__2921\ : Span4Mux_s2_v
    port map (
            O => \N__17368\,
            I => \N__17327\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__17365\,
            I => \N__17327\
        );

    \I__2919\ : InMux
    port map (
            O => \N__17362\,
            I => \N__17324\
        );

    \I__2918\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17321\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__17358\,
            I => \N__17318\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__17355\,
            I => \N__17313\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__17352\,
            I => \N__17313\
        );

    \I__2914\ : InMux
    port map (
            O => \N__17349\,
            I => \N__17310\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__17348\,
            I => \N__17307\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__17347\,
            I => \N__17304\
        );

    \I__2911\ : Span4Mux_v
    port map (
            O => \N__17344\,
            I => \N__17301\
        );

    \I__2910\ : InMux
    port map (
            O => \N__17341\,
            I => \N__17298\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__17338\,
            I => \N__17295\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__17335\,
            I => \N__17292\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__17332\,
            I => \N__17289\
        );

    \I__2906\ : Span4Mux_v
    port map (
            O => \N__17327\,
            I => \N__17284\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__17324\,
            I => \N__17284\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__17321\,
            I => \N__17281\
        );

    \I__2903\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17278\
        );

    \I__2902\ : Span4Mux_v
    port map (
            O => \N__17313\,
            I => \N__17272\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__17310\,
            I => \N__17272\
        );

    \I__2900\ : InMux
    port map (
            O => \N__17307\,
            I => \N__17269\
        );

    \I__2899\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17266\
        );

    \I__2898\ : Sp12to4
    port map (
            O => \N__17301\,
            I => \N__17261\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__17298\,
            I => \N__17261\
        );

    \I__2896\ : Span4Mux_h
    port map (
            O => \N__17295\,
            I => \N__17258\
        );

    \I__2895\ : Span4Mux_h
    port map (
            O => \N__17292\,
            I => \N__17255\
        );

    \I__2894\ : Span4Mux_h
    port map (
            O => \N__17289\,
            I => \N__17252\
        );

    \I__2893\ : Span4Mux_v
    port map (
            O => \N__17284\,
            I => \N__17245\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__17281\,
            I => \N__17245\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__17278\,
            I => \N__17245\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__17277\,
            I => \N__17242\
        );

    \I__2889\ : Span4Mux_v
    port map (
            O => \N__17272\,
            I => \N__17237\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__17269\,
            I => \N__17237\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__17266\,
            I => \N__17234\
        );

    \I__2886\ : Span12Mux_h
    port map (
            O => \N__17261\,
            I => \N__17231\
        );

    \I__2885\ : Sp12to4
    port map (
            O => \N__17258\,
            I => \N__17224\
        );

    \I__2884\ : Sp12to4
    port map (
            O => \N__17255\,
            I => \N__17224\
        );

    \I__2883\ : Sp12to4
    port map (
            O => \N__17252\,
            I => \N__17224\
        );

    \I__2882\ : Span4Mux_v
    port map (
            O => \N__17245\,
            I => \N__17221\
        );

    \I__2881\ : InMux
    port map (
            O => \N__17242\,
            I => \N__17218\
        );

    \I__2880\ : Span4Mux_h
    port map (
            O => \N__17237\,
            I => \N__17215\
        );

    \I__2879\ : Span12Mux_h
    port map (
            O => \N__17234\,
            I => \N__17212\
        );

    \I__2878\ : Span12Mux_v
    port map (
            O => \N__17231\,
            I => \N__17203\
        );

    \I__2877\ : Span12Mux_v
    port map (
            O => \N__17224\,
            I => \N__17203\
        );

    \I__2876\ : Sp12to4
    port map (
            O => \N__17221\,
            I => \N__17203\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__17218\,
            I => \N__17203\
        );

    \I__2874\ : Span4Mux_h
    port map (
            O => \N__17215\,
            I => \N__17200\
        );

    \I__2873\ : Odrv12
    port map (
            O => \N__17212\,
            I => \M_this_ppu_sprites_addr_7\
        );

    \I__2872\ : Odrv12
    port map (
            O => \N__17203\,
            I => \M_this_ppu_sprites_addr_7\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__17200\,
            I => \M_this_ppu_sprites_addr_7\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__17193\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_7_cascade_\
        );

    \I__2869\ : InMux
    port map (
            O => \N__17190\,
            I => \N__17186\
        );

    \I__2868\ : InMux
    port map (
            O => \N__17189\,
            I => \N__17183\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__17186\,
            I => \this_vga_signals.un4_lvisibility_1\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__17183\,
            I => \this_vga_signals.un4_lvisibility_1\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__17178\,
            I => \N__17173\
        );

    \I__2864\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17163\
        );

    \I__2863\ : InMux
    port map (
            O => \N__17176\,
            I => \N__17160\
        );

    \I__2862\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17157\
        );

    \I__2861\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17154\
        );

    \I__2860\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17151\
        );

    \I__2859\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17146\
        );

    \I__2858\ : InMux
    port map (
            O => \N__17169\,
            I => \N__17146\
        );

    \I__2857\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17143\
        );

    \I__2856\ : InMux
    port map (
            O => \N__17167\,
            I => \N__17140\
        );

    \I__2855\ : InMux
    port map (
            O => \N__17166\,
            I => \N__17137\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__17163\,
            I => \N__17129\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__17160\,
            I => \N__17129\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__17157\,
            I => \N__17129\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__17154\,
            I => \N__17126\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__17151\,
            I => \N__17123\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__17146\,
            I => \N__17111\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__17143\,
            I => \N__17111\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__17140\,
            I => \N__17111\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__17137\,
            I => \N__17111\
        );

    \I__2845\ : InMux
    port map (
            O => \N__17136\,
            I => \N__17108\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__17129\,
            I => \N__17105\
        );

    \I__2843\ : Span4Mux_v
    port map (
            O => \N__17126\,
            I => \N__17100\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__17123\,
            I => \N__17100\
        );

    \I__2841\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17095\
        );

    \I__2840\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17095\
        );

    \I__2839\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17092\
        );

    \I__2838\ : Span4Mux_v
    port map (
            O => \N__17111\,
            I => \N__17087\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__17108\,
            I => \N__17087\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__17105\,
            I => \N__17084\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__17100\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__17095\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__17092\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__17087\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__17084\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2830\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17069\
        );

    \I__2829\ : InMux
    port map (
            O => \N__17072\,
            I => \N__17063\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__17069\,
            I => \N__17060\
        );

    \I__2827\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17057\
        );

    \I__2826\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17052\
        );

    \I__2825\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17052\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__17063\,
            I => \N__17042\
        );

    \I__2823\ : Span4Mux_v
    port map (
            O => \N__17060\,
            I => \N__17042\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__17057\,
            I => \N__17039\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__17052\,
            I => \N__17036\
        );

    \I__2820\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17031\
        );

    \I__2819\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17031\
        );

    \I__2818\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17028\
        );

    \I__2817\ : InMux
    port map (
            O => \N__17048\,
            I => \N__17025\
        );

    \I__2816\ : InMux
    port map (
            O => \N__17047\,
            I => \N__17022\
        );

    \I__2815\ : Span4Mux_h
    port map (
            O => \N__17042\,
            I => \N__17011\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__17039\,
            I => \N__17011\
        );

    \I__2813\ : Sp12to4
    port map (
            O => \N__17036\,
            I => \N__17004\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__17031\,
            I => \N__17004\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__17028\,
            I => \N__17004\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__17025\,
            I => \N__16999\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__17022\,
            I => \N__16999\
        );

    \I__2808\ : InMux
    port map (
            O => \N__17021\,
            I => \N__16994\
        );

    \I__2807\ : InMux
    port map (
            O => \N__17020\,
            I => \N__16994\
        );

    \I__2806\ : InMux
    port map (
            O => \N__17019\,
            I => \N__16991\
        );

    \I__2805\ : InMux
    port map (
            O => \N__17018\,
            I => \N__16988\
        );

    \I__2804\ : InMux
    port map (
            O => \N__17017\,
            I => \N__16983\
        );

    \I__2803\ : InMux
    port map (
            O => \N__17016\,
            I => \N__16983\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__17011\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2801\ : Odrv12
    port map (
            O => \N__17004\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2800\ : Odrv12
    port map (
            O => \N__16999\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__16994\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__16991\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__16988\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__16983\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2795\ : InMux
    port map (
            O => \N__16968\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1\
        );

    \I__2794\ : InMux
    port map (
            O => \N__16965\,
            I => \N__16961\
        );

    \I__2793\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16958\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__16961\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__16958\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__2790\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16950\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__16950\,
            I => \M_this_data_count_q_cry_3_THRU_CO\
        );

    \I__2788\ : InMux
    port map (
            O => \N__16947\,
            I => \N__16942\
        );

    \I__2787\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16937\
        );

    \I__2786\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16937\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__16942\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__16937\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__2783\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16929\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__16929\,
            I => \N__16926\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__16926\,
            I => \M_this_data_count_q_cry_4_THRU_CO\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__16923\,
            I => \N__16920\
        );

    \I__2779\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16915\
        );

    \I__2778\ : InMux
    port map (
            O => \N__16919\,
            I => \N__16910\
        );

    \I__2777\ : InMux
    port map (
            O => \N__16918\,
            I => \N__16910\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__16915\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__16910\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__2774\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16902\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__16902\,
            I => \M_this_data_count_q_cry_6_THRU_CO\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__16899\,
            I => \N__16895\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__16898\,
            I => \N__16891\
        );

    \I__2770\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16888\
        );

    \I__2769\ : InMux
    port map (
            O => \N__16894\,
            I => \N__16883\
        );

    \I__2768\ : InMux
    port map (
            O => \N__16891\,
            I => \N__16883\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__16888\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__16883\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__2765\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16875\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__16875\,
            I => \M_this_data_count_q_cry_2_THRU_CO\
        );

    \I__2763\ : InMux
    port map (
            O => \N__16872\,
            I => \N__16869\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__16869\,
            I => \M_this_data_count_q_cry_10_THRU_CO\
        );

    \I__2761\ : InMux
    port map (
            O => \N__16866\,
            I => \N__16863\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__16863\,
            I => \M_this_data_count_q_cry_11_THRU_CO\
        );

    \I__2759\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16855\
        );

    \I__2758\ : InMux
    port map (
            O => \N__16859\,
            I => \N__16850\
        );

    \I__2757\ : InMux
    port map (
            O => \N__16858\,
            I => \N__16850\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__16855\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__16850\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__16845\,
            I => \N__16841\
        );

    \I__2753\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16838\
        );

    \I__2752\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16835\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__16838\,
            I => \N__16830\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__16835\,
            I => \N__16830\
        );

    \I__2749\ : Odrv4
    port map (
            O => \N__16830\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__2748\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16824\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__16824\,
            I => \M_this_data_count_q_cry_7_THRU_CO\
        );

    \I__2746\ : InMux
    port map (
            O => \N__16821\,
            I => \N__16816\
        );

    \I__2745\ : InMux
    port map (
            O => \N__16820\,
            I => \N__16811\
        );

    \I__2744\ : InMux
    port map (
            O => \N__16819\,
            I => \N__16811\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__16816\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__16811\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__2741\ : InMux
    port map (
            O => \N__16806\,
            I => \N__16803\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__16803\,
            I => \M_this_state_q_RNIOE1SZ0Z_11\
        );

    \I__2739\ : InMux
    port map (
            O => \N__16800\,
            I => \N__16797\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__16797\,
            I => un20_i_a2_x_3
        );

    \I__2737\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16791\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__16791\,
            I => \M_this_state_q_RNIG01LZ0Z_12\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__16788\,
            I => \this_vga_signals.N_419_i_i_0Z0Z_1_cascade_\
        );

    \I__2734\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16782\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__16782\,
            I => \M_this_data_count_q_s_6\
        );

    \I__2732\ : CascadeMux
    port map (
            O => \N__16779\,
            I => \N__16772\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__16778\,
            I => \N__16768\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__16777\,
            I => \N__16761\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__16776\,
            I => \N__16757\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__16775\,
            I => \N__16754\
        );

    \I__2727\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16744\
        );

    \I__2726\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16744\
        );

    \I__2725\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16744\
        );

    \I__2724\ : InMux
    port map (
            O => \N__16767\,
            I => \N__16744\
        );

    \I__2723\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16737\
        );

    \I__2722\ : InMux
    port map (
            O => \N__16765\,
            I => \N__16737\
        );

    \I__2721\ : InMux
    port map (
            O => \N__16764\,
            I => \N__16731\
        );

    \I__2720\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16731\
        );

    \I__2719\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16728\
        );

    \I__2718\ : InMux
    port map (
            O => \N__16757\,
            I => \N__16725\
        );

    \I__2717\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16722\
        );

    \I__2716\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16719\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__16744\,
            I => \N__16716\
        );

    \I__2714\ : InMux
    port map (
            O => \N__16743\,
            I => \N__16713\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__16742\,
            I => \N__16708\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__16737\,
            I => \N__16704\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__16736\,
            I => \N__16700\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__16731\,
            I => \N__16697\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__16728\,
            I => \N__16692\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__16725\,
            I => \N__16692\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__16722\,
            I => \N__16687\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__16719\,
            I => \N__16682\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__16716\,
            I => \N__16677\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__16713\,
            I => \N__16677\
        );

    \I__2703\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16668\
        );

    \I__2702\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16668\
        );

    \I__2701\ : InMux
    port map (
            O => \N__16708\,
            I => \N__16668\
        );

    \I__2700\ : InMux
    port map (
            O => \N__16707\,
            I => \N__16668\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__16704\,
            I => \N__16665\
        );

    \I__2698\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16662\
        );

    \I__2697\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16659\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__16697\,
            I => \N__16656\
        );

    \I__2695\ : Span4Mux_v
    port map (
            O => \N__16692\,
            I => \N__16653\
        );

    \I__2694\ : InMux
    port map (
            O => \N__16691\,
            I => \N__16648\
        );

    \I__2693\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16648\
        );

    \I__2692\ : Span4Mux_h
    port map (
            O => \N__16687\,
            I => \N__16645\
        );

    \I__2691\ : InMux
    port map (
            O => \N__16686\,
            I => \N__16640\
        );

    \I__2690\ : InMux
    port map (
            O => \N__16685\,
            I => \N__16640\
        );

    \I__2689\ : Span4Mux_v
    port map (
            O => \N__16682\,
            I => \N__16635\
        );

    \I__2688\ : Span4Mux_h
    port map (
            O => \N__16677\,
            I => \N__16635\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__16668\,
            I => \N__16630\
        );

    \I__2686\ : Span4Mux_h
    port map (
            O => \N__16665\,
            I => \N__16630\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__16662\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__16659\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2683\ : Odrv4
    port map (
            O => \N__16656\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__16653\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__16648\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__16645\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__16640\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__16635\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__16630\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2676\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16603\
        );

    \I__2675\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16603\
        );

    \I__2674\ : InMux
    port map (
            O => \N__16609\,
            I => \N__16593\
        );

    \I__2673\ : InMux
    port map (
            O => \N__16608\,
            I => \N__16590\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__16603\,
            I => \N__16587\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__16602\,
            I => \N__16584\
        );

    \I__2670\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16578\
        );

    \I__2669\ : InMux
    port map (
            O => \N__16600\,
            I => \N__16578\
        );

    \I__2668\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16571\
        );

    \I__2667\ : InMux
    port map (
            O => \N__16598\,
            I => \N__16571\
        );

    \I__2666\ : InMux
    port map (
            O => \N__16597\,
            I => \N__16571\
        );

    \I__2665\ : InMux
    port map (
            O => \N__16596\,
            I => \N__16568\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__16593\,
            I => \N__16565\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__16590\,
            I => \N__16560\
        );

    \I__2662\ : Span4Mux_h
    port map (
            O => \N__16587\,
            I => \N__16560\
        );

    \I__2661\ : InMux
    port map (
            O => \N__16584\,
            I => \N__16557\
        );

    \I__2660\ : InMux
    port map (
            O => \N__16583\,
            I => \N__16554\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__16578\,
            I => \N__16551\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__16571\,
            I => \N__16535\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__16568\,
            I => \N__16535\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__16565\,
            I => \N__16535\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__16560\,
            I => \N__16535\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__16557\,
            I => \N__16535\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__16554\,
            I => \N__16535\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__16551\,
            I => \N__16531\
        );

    \I__2651\ : InMux
    port map (
            O => \N__16550\,
            I => \N__16526\
        );

    \I__2650\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16526\
        );

    \I__2649\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16523\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__16535\,
            I => \N__16520\
        );

    \I__2647\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16517\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__16531\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__16526\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__16523\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__16520\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__16517\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__16506\,
            I => \N__16503\
        );

    \I__2640\ : InMux
    port map (
            O => \N__16503\,
            I => \N__16497\
        );

    \I__2639\ : InMux
    port map (
            O => \N__16502\,
            I => \N__16497\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__16497\,
            I => \this_vga_signals.M_vcounter_d7lt8_0\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__16494\,
            I => \this_vga_signals.M_vcounter_d7lto8_1_cascade_\
        );

    \I__2636\ : InMux
    port map (
            O => \N__16491\,
            I => \N__16485\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__16490\,
            I => \N__16470\
        );

    \I__2634\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16466\
        );

    \I__2633\ : InMux
    port map (
            O => \N__16488\,
            I => \N__16463\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__16485\,
            I => \N__16460\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__16484\,
            I => \N__16452\
        );

    \I__2630\ : InMux
    port map (
            O => \N__16483\,
            I => \N__16446\
        );

    \I__2629\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16446\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__16481\,
            I => \N__16443\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__16480\,
            I => \N__16440\
        );

    \I__2626\ : InMux
    port map (
            O => \N__16479\,
            I => \N__16437\
        );

    \I__2625\ : InMux
    port map (
            O => \N__16478\,
            I => \N__16434\
        );

    \I__2624\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16431\
        );

    \I__2623\ : InMux
    port map (
            O => \N__16476\,
            I => \N__16428\
        );

    \I__2622\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16415\
        );

    \I__2621\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16415\
        );

    \I__2620\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16415\
        );

    \I__2619\ : InMux
    port map (
            O => \N__16470\,
            I => \N__16415\
        );

    \I__2618\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16412\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__16466\,
            I => \N__16405\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__16463\,
            I => \N__16405\
        );

    \I__2615\ : Span4Mux_h
    port map (
            O => \N__16460\,
            I => \N__16405\
        );

    \I__2614\ : InMux
    port map (
            O => \N__16459\,
            I => \N__16400\
        );

    \I__2613\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16400\
        );

    \I__2612\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16395\
        );

    \I__2611\ : InMux
    port map (
            O => \N__16456\,
            I => \N__16395\
        );

    \I__2610\ : InMux
    port map (
            O => \N__16455\,
            I => \N__16389\
        );

    \I__2609\ : InMux
    port map (
            O => \N__16452\,
            I => \N__16389\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__16451\,
            I => \N__16386\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__16446\,
            I => \N__16382\
        );

    \I__2606\ : InMux
    port map (
            O => \N__16443\,
            I => \N__16377\
        );

    \I__2605\ : InMux
    port map (
            O => \N__16440\,
            I => \N__16377\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__16437\,
            I => \N__16370\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__16434\,
            I => \N__16370\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__16431\,
            I => \N__16370\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__16428\,
            I => \N__16367\
        );

    \I__2600\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16357\
        );

    \I__2599\ : InMux
    port map (
            O => \N__16426\,
            I => \N__16357\
        );

    \I__2598\ : InMux
    port map (
            O => \N__16425\,
            I => \N__16357\
        );

    \I__2597\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16357\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__16415\,
            I => \N__16354\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__16412\,
            I => \N__16347\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__16405\,
            I => \N__16347\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__16400\,
            I => \N__16347\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__16395\,
            I => \N__16344\
        );

    \I__2591\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16341\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__16389\,
            I => \N__16338\
        );

    \I__2589\ : InMux
    port map (
            O => \N__16386\,
            I => \N__16333\
        );

    \I__2588\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16333\
        );

    \I__2587\ : Span4Mux_h
    port map (
            O => \N__16382\,
            I => \N__16324\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__16377\,
            I => \N__16324\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__16370\,
            I => \N__16324\
        );

    \I__2584\ : Span4Mux_h
    port map (
            O => \N__16367\,
            I => \N__16324\
        );

    \I__2583\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16321\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__16357\,
            I => \N__16312\
        );

    \I__2581\ : Span4Mux_h
    port map (
            O => \N__16354\,
            I => \N__16312\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__16347\,
            I => \N__16312\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__16344\,
            I => \N__16312\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__16341\,
            I => \N__16307\
        );

    \I__2577\ : Span4Mux_h
    port map (
            O => \N__16338\,
            I => \N__16307\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__16333\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__16324\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__16321\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__16312\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2572\ : Odrv4
    port map (
            O => \N__16307\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__16296\,
            I => \this_vga_signals.M_vcounter_d8_cascade_\
        );

    \I__2570\ : IoInMux
    port map (
            O => \N__16293\,
            I => \N__16290\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__16290\,
            I => \N__16287\
        );

    \I__2568\ : Span12Mux_s7_h
    port map (
            O => \N__16287\,
            I => \N__16284\
        );

    \I__2567\ : Odrv12
    port map (
            O => \N__16284\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\
        );

    \I__2566\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16276\
        );

    \I__2565\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16271\
        );

    \I__2564\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16271\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__16276\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__16271\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__16266\,
            I => \N__16260\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__16265\,
            I => \N__16256\
        );

    \I__2559\ : InMux
    port map (
            O => \N__16264\,
            I => \N__16252\
        );

    \I__2558\ : InMux
    port map (
            O => \N__16263\,
            I => \N__16249\
        );

    \I__2557\ : InMux
    port map (
            O => \N__16260\,
            I => \N__16240\
        );

    \I__2556\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16240\
        );

    \I__2555\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16240\
        );

    \I__2554\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16240\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__16252\,
            I => \M_pcounter_q_ret_2_RNIH7PG8\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__16249\,
            I => \M_pcounter_q_ret_2_RNIH7PG8\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__16240\,
            I => \M_pcounter_q_ret_2_RNIH7PG8\
        );

    \I__2550\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16230\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__16230\,
            I => \N__16226\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__16229\,
            I => \N__16223\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__16226\,
            I => \N__16220\
        );

    \I__2546\ : InMux
    port map (
            O => \N__16223\,
            I => \N__16217\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__16220\,
            I => \this_vga_ramdac.N_2865_reto\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__16217\,
            I => \this_vga_ramdac.N_2865_reto\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__16212\,
            I => \dma_ac0_5_0_cascade_\
        );

    \I__2542\ : InMux
    port map (
            O => \N__16209\,
            I => \M_this_data_count_q_cry_8\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__16206\,
            I => \N__16203\
        );

    \I__2540\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16200\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__16200\,
            I => \N__16197\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__16197\,
            I => \M_this_data_count_q_s_10\
        );

    \I__2537\ : InMux
    port map (
            O => \N__16194\,
            I => \M_this_data_count_q_cry_9\
        );

    \I__2536\ : InMux
    port map (
            O => \N__16191\,
            I => \M_this_data_count_q_cry_10\
        );

    \I__2535\ : InMux
    port map (
            O => \N__16188\,
            I => \M_this_data_count_q_cry_11\
        );

    \I__2534\ : InMux
    port map (
            O => \N__16185\,
            I => \M_this_data_count_q_cry_12\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__16182\,
            I => \N__16179\
        );

    \I__2532\ : InMux
    port map (
            O => \N__16179\,
            I => \N__16176\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__16176\,
            I => \N__16173\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__16173\,
            I => \M_this_data_count_q_s_13\
        );

    \I__2529\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16167\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__16167\,
            I => \N__16164\
        );

    \I__2527\ : Span12Mux_h
    port map (
            O => \N__16164\,
            I => \N__16161\
        );

    \I__2526\ : Odrv12
    port map (
            O => \N__16161\,
            I => \N_87_0\
        );

    \I__2525\ : InMux
    port map (
            O => \N__16158\,
            I => \N__16155\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__16155\,
            I => \N__16152\
        );

    \I__2523\ : Odrv12
    port map (
            O => \N__16152\,
            I => \N_81_0\
        );

    \I__2522\ : InMux
    port map (
            O => \N__16149\,
            I => \M_this_data_count_q_cry_0\
        );

    \I__2521\ : InMux
    port map (
            O => \N__16146\,
            I => \M_this_data_count_q_cry_1\
        );

    \I__2520\ : InMux
    port map (
            O => \N__16143\,
            I => \M_this_data_count_q_cry_2\
        );

    \I__2519\ : InMux
    port map (
            O => \N__16140\,
            I => \M_this_data_count_q_cry_3\
        );

    \I__2518\ : InMux
    port map (
            O => \N__16137\,
            I => \M_this_data_count_q_cry_4\
        );

    \I__2517\ : InMux
    port map (
            O => \N__16134\,
            I => \M_this_data_count_q_cry_5\
        );

    \I__2516\ : InMux
    port map (
            O => \N__16131\,
            I => \M_this_data_count_q_cry_6\
        );

    \I__2515\ : InMux
    port map (
            O => \N__16128\,
            I => \bfn_14_26_0_\
        );

    \I__2514\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16122\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__16122\,
            I => \N__16119\
        );

    \I__2512\ : Span4Mux_h
    port map (
            O => \N__16119\,
            I => \N__16116\
        );

    \I__2511\ : Span4Mux_h
    port map (
            O => \N__16116\,
            I => \N__16113\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__16113\,
            I => \this_vga_ramdac.i2_mux\
        );

    \I__2509\ : InMux
    port map (
            O => \N__16110\,
            I => \N__16106\
        );

    \I__2508\ : InMux
    port map (
            O => \N__16109\,
            I => \N__16103\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__16106\,
            I => \this_vga_ramdac.N_2864_reto\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__16103\,
            I => \this_vga_ramdac.N_2864_reto\
        );

    \I__2505\ : IoInMux
    port map (
            O => \N__16098\,
            I => \N__16091\
        );

    \I__2504\ : IoInMux
    port map (
            O => \N__16097\,
            I => \N__16088\
        );

    \I__2503\ : IoInMux
    port map (
            O => \N__16096\,
            I => \N__16085\
        );

    \I__2502\ : IoInMux
    port map (
            O => \N__16095\,
            I => \N__16080\
        );

    \I__2501\ : IoInMux
    port map (
            O => \N__16094\,
            I => \N__16077\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__16091\,
            I => \N__16072\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__16088\,
            I => \N__16072\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__16085\,
            I => \N__16069\
        );

    \I__2497\ : IoInMux
    port map (
            O => \N__16084\,
            I => \N__16066\
        );

    \I__2496\ : IoInMux
    port map (
            O => \N__16083\,
            I => \N__16063\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__16080\,
            I => \N__16058\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__16077\,
            I => \N__16053\
        );

    \I__2493\ : IoSpan4Mux
    port map (
            O => \N__16072\,
            I => \N__16050\
        );

    \I__2492\ : IoSpan4Mux
    port map (
            O => \N__16069\,
            I => \N__16043\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__16066\,
            I => \N__16043\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__16063\,
            I => \N__16043\
        );

    \I__2489\ : IoInMux
    port map (
            O => \N__16062\,
            I => \N__16040\
        );

    \I__2488\ : IoInMux
    port map (
            O => \N__16061\,
            I => \N__16037\
        );

    \I__2487\ : IoSpan4Mux
    port map (
            O => \N__16058\,
            I => \N__16034\
        );

    \I__2486\ : IoInMux
    port map (
            O => \N__16057\,
            I => \N__16031\
        );

    \I__2485\ : IoInMux
    port map (
            O => \N__16056\,
            I => \N__16028\
        );

    \I__2484\ : IoSpan4Mux
    port map (
            O => \N__16053\,
            I => \N__16023\
        );

    \I__2483\ : Span4Mux_s1_h
    port map (
            O => \N__16050\,
            I => \N__16019\
        );

    \I__2482\ : IoSpan4Mux
    port map (
            O => \N__16043\,
            I => \N__16012\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__16040\,
            I => \N__16012\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__16037\,
            I => \N__16012\
        );

    \I__2479\ : IoSpan4Mux
    port map (
            O => \N__16034\,
            I => \N__16007\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__16031\,
            I => \N__16007\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__16028\,
            I => \N__16004\
        );

    \I__2476\ : IoInMux
    port map (
            O => \N__16027\,
            I => \N__16001\
        );

    \I__2475\ : IoInMux
    port map (
            O => \N__16026\,
            I => \N__15996\
        );

    \I__2474\ : Span4Mux_s3_h
    port map (
            O => \N__16023\,
            I => \N__15993\
        );

    \I__2473\ : IoInMux
    port map (
            O => \N__16022\,
            I => \N__15990\
        );

    \I__2472\ : Span4Mux_h
    port map (
            O => \N__16019\,
            I => \N__15984\
        );

    \I__2471\ : IoSpan4Mux
    port map (
            O => \N__16012\,
            I => \N__15984\
        );

    \I__2470\ : IoSpan4Mux
    port map (
            O => \N__16007\,
            I => \N__15977\
        );

    \I__2469\ : IoSpan4Mux
    port map (
            O => \N__16004\,
            I => \N__15977\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__16001\,
            I => \N__15977\
        );

    \I__2467\ : IoInMux
    port map (
            O => \N__16000\,
            I => \N__15974\
        );

    \I__2466\ : IoInMux
    port map (
            O => \N__15999\,
            I => \N__15971\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__15996\,
            I => \N__15968\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__15993\,
            I => \N__15965\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__15990\,
            I => \N__15962\
        );

    \I__2462\ : IoInMux
    port map (
            O => \N__15989\,
            I => \N__15959\
        );

    \I__2461\ : Span4Mux_s1_h
    port map (
            O => \N__15984\,
            I => \N__15956\
        );

    \I__2460\ : IoSpan4Mux
    port map (
            O => \N__15977\,
            I => \N__15949\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__15974\,
            I => \N__15949\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__15971\,
            I => \N__15949\
        );

    \I__2457\ : IoSpan4Mux
    port map (
            O => \N__15968\,
            I => \N__15946\
        );

    \I__2456\ : Sp12to4
    port map (
            O => \N__15965\,
            I => \N__15941\
        );

    \I__2455\ : Span12Mux_s6_h
    port map (
            O => \N__15962\,
            I => \N__15941\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__15959\,
            I => \N__15938\
        );

    \I__2453\ : Sp12to4
    port map (
            O => \N__15956\,
            I => \N__15935\
        );

    \I__2452\ : IoSpan4Mux
    port map (
            O => \N__15949\,
            I => \N__15932\
        );

    \I__2451\ : Span4Mux_s2_h
    port map (
            O => \N__15946\,
            I => \N__15929\
        );

    \I__2450\ : Span12Mux_h
    port map (
            O => \N__15941\,
            I => \N__15926\
        );

    \I__2449\ : Span12Mux_s2_v
    port map (
            O => \N__15938\,
            I => \N__15923\
        );

    \I__2448\ : Span12Mux_s6_h
    port map (
            O => \N__15935\,
            I => \N__15920\
        );

    \I__2447\ : Span4Mux_s2_v
    port map (
            O => \N__15932\,
            I => \N__15917\
        );

    \I__2446\ : Span4Mux_h
    port map (
            O => \N__15929\,
            I => \N__15914\
        );

    \I__2445\ : Span12Mux_v
    port map (
            O => \N__15926\,
            I => \N__15905\
        );

    \I__2444\ : Span12Mux_h
    port map (
            O => \N__15923\,
            I => \N__15905\
        );

    \I__2443\ : Span12Mux_h
    port map (
            O => \N__15920\,
            I => \N__15905\
        );

    \I__2442\ : Sp12to4
    port map (
            O => \N__15917\,
            I => \N__15905\
        );

    \I__2441\ : Span4Mux_h
    port map (
            O => \N__15914\,
            I => \N__15902\
        );

    \I__2440\ : Odrv12
    port map (
            O => \N__15905\,
            I => dma_0_i
        );

    \I__2439\ : Odrv4
    port map (
            O => \N__15902\,
            I => dma_0_i
        );

    \I__2438\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15892\
        );

    \I__2437\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15887\
        );

    \I__2436\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15887\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__15892\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__15887\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2433\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15879\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__15879\,
            I => \this_vga_signals.M_pcounter_q_3_0\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__15876\,
            I => \N__15871\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__15875\,
            I => \N__15868\
        );

    \I__2429\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15865\
        );

    \I__2428\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15860\
        );

    \I__2427\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15860\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__15865\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__15860\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__2424\ : InMux
    port map (
            O => \N__15855\,
            I => \N__15852\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__15852\,
            I => \this_vga_signals.M_pcounter_q_3_1\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__15849\,
            I => \N__15846\
        );

    \I__2421\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15840\
        );

    \I__2420\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15840\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__15840\,
            I => \this_vga_signals.N_3_0\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__15837\,
            I => \this_vga_signals.N_3_0_cascade_\
        );

    \I__2417\ : InMux
    port map (
            O => \N__15834\,
            I => \N__15822\
        );

    \I__2416\ : InMux
    port map (
            O => \N__15833\,
            I => \N__15822\
        );

    \I__2415\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15822\
        );

    \I__2414\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15822\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__15822\,
            I => \this_vga_signals.M_pcounter_q_i_3_1\
        );

    \I__2412\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15812\
        );

    \I__2411\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15812\
        );

    \I__2410\ : InMux
    port map (
            O => \N__15817\,
            I => \N__15809\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__15812\,
            I => \N__15806\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__15809\,
            I => \N__15801\
        );

    \I__2407\ : Span4Mux_h
    port map (
            O => \N__15806\,
            I => \N__15798\
        );

    \I__2406\ : InMux
    port map (
            O => \N__15805\,
            I => \N__15795\
        );

    \I__2405\ : InMux
    port map (
            O => \N__15804\,
            I => \N__15792\
        );

    \I__2404\ : Span4Mux_v
    port map (
            O => \N__15801\,
            I => \N__15787\
        );

    \I__2403\ : Span4Mux_h
    port map (
            O => \N__15798\,
            I => \N__15780\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__15795\,
            I => \N__15780\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__15792\,
            I => \N__15780\
        );

    \I__2400\ : InMux
    port map (
            O => \N__15791\,
            I => \N__15777\
        );

    \I__2399\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15774\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__15787\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__2397\ : Odrv4
    port map (
            O => \N__15780\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__15777\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__15774\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__2394\ : InMux
    port map (
            O => \N__15765\,
            I => \N__15762\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__15762\,
            I => \N__15758\
        );

    \I__2392\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15755\
        );

    \I__2391\ : Odrv12
    port map (
            O => \N__15758\,
            I => \this_vga_ramdac.N_2867_reto\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__15755\,
            I => \this_vga_ramdac.N_2867_reto\
        );

    \I__2389\ : IoInMux
    port map (
            O => \N__15750\,
            I => \N__15747\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__15747\,
            I => \N__15744\
        );

    \I__2387\ : Span4Mux_s3_h
    port map (
            O => \N__15744\,
            I => \N__15741\
        );

    \I__2386\ : Span4Mux_h
    port map (
            O => \N__15741\,
            I => \N__15738\
        );

    \I__2385\ : Sp12to4
    port map (
            O => \N__15738\,
            I => \N__15735\
        );

    \I__2384\ : Span12Mux_s11_v
    port map (
            O => \N__15735\,
            I => \N__15732\
        );

    \I__2383\ : Odrv12
    port map (
            O => \N__15732\,
            I => rgb_c_5
        );

    \I__2382\ : InMux
    port map (
            O => \N__15729\,
            I => \N__15724\
        );

    \I__2381\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15719\
        );

    \I__2380\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15719\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__15724\,
            I => \this_vga_signals.N_2_0\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__15719\,
            I => \this_vga_signals.N_2_0\
        );

    \I__2377\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15710\
        );

    \I__2376\ : InMux
    port map (
            O => \N__15713\,
            I => \N__15707\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__15710\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__15707\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__2373\ : InMux
    port map (
            O => \N__15702\,
            I => \N__15696\
        );

    \I__2372\ : InMux
    port map (
            O => \N__15701\,
            I => \N__15696\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__15696\,
            I => \this_pixel_clk_M_counter_q_i_1\
        );

    \I__2370\ : IoInMux
    port map (
            O => \N__15693\,
            I => \N__15690\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__15690\,
            I => \N__15687\
        );

    \I__2368\ : Span4Mux_s1_h
    port map (
            O => \N__15687\,
            I => \N__15684\
        );

    \I__2367\ : Span4Mux_h
    port map (
            O => \N__15684\,
            I => \N__15681\
        );

    \I__2366\ : Span4Mux_h
    port map (
            O => \N__15681\,
            I => \N__15678\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__15678\,
            I => \N__15675\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__15675\,
            I => rgb_c_2
        );

    \I__2363\ : InMux
    port map (
            O => \N__15672\,
            I => \N__15669\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__15669\,
            I => \N__15666\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__15666\,
            I => \this_vga_ramdac.m6\
        );

    \I__2360\ : InMux
    port map (
            O => \N__15663\,
            I => \N__15660\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__15660\,
            I => \N__15657\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__15657\,
            I => \N__15654\
        );

    \I__2357\ : Span4Mux_h
    port map (
            O => \N__15654\,
            I => \N__15650\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__15653\,
            I => \N__15647\
        );

    \I__2355\ : Span4Mux_h
    port map (
            O => \N__15650\,
            I => \N__15644\
        );

    \I__2354\ : InMux
    port map (
            O => \N__15647\,
            I => \N__15641\
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__15644\,
            I => \this_vga_ramdac.N_2863_reto\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__15641\,
            I => \this_vga_ramdac.N_2863_reto\
        );

    \I__2351\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15633\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__15633\,
            I => \N__15630\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__15630\,
            I => \this_vga_ramdac.i2_mux_0\
        );

    \I__2348\ : InMux
    port map (
            O => \N__15627\,
            I => \N__15624\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__15624\,
            I => \N__15621\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__15621\,
            I => \this_vga_ramdac.m19\
        );

    \I__2345\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15615\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__15615\,
            I => \N__15611\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__15614\,
            I => \N__15608\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__15611\,
            I => \N__15605\
        );

    \I__2341\ : InMux
    port map (
            O => \N__15608\,
            I => \N__15602\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__15605\,
            I => \this_vga_ramdac.N_2866_reto\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__15602\,
            I => \this_vga_ramdac.N_2866_reto\
        );

    \I__2338\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15594\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__15594\,
            I => \this_vga_signals.M_this_vga_signals_pixel_clk_0_0\
        );

    \I__2336\ : InMux
    port map (
            O => \N__15591\,
            I => \N__15584\
        );

    \I__2335\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15581\
        );

    \I__2334\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15578\
        );

    \I__2333\ : InMux
    port map (
            O => \N__15588\,
            I => \N__15573\
        );

    \I__2332\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15573\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__15584\,
            I => \N__15570\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__15581\,
            I => \N__15567\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__15578\,
            I => \N__15562\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__15573\,
            I => \N__15562\
        );

    \I__2327\ : Span4Mux_h
    port map (
            O => \N__15570\,
            I => \N__15555\
        );

    \I__2326\ : Span4Mux_h
    port map (
            O => \N__15567\,
            I => \N__15552\
        );

    \I__2325\ : Span4Mux_h
    port map (
            O => \N__15562\,
            I => \N__15549\
        );

    \I__2324\ : InMux
    port map (
            O => \N__15561\,
            I => \N__15546\
        );

    \I__2323\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15541\
        );

    \I__2322\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15541\
        );

    \I__2321\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15538\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__15555\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__15552\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__15549\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__15546\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__15541\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__15538\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__15525\,
            I => \M_pcounter_q_ret_2_RNIH7PG8_cascade_\
        );

    \I__2313\ : IoInMux
    port map (
            O => \N__15522\,
            I => \N__15519\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__15519\,
            I => \N__15516\
        );

    \I__2311\ : IoSpan4Mux
    port map (
            O => \N__15516\,
            I => \N__15513\
        );

    \I__2310\ : Span4Mux_s2_h
    port map (
            O => \N__15513\,
            I => \N__15510\
        );

    \I__2309\ : Span4Mux_h
    port map (
            O => \N__15510\,
            I => \N__15507\
        );

    \I__2308\ : Span4Mux_h
    port map (
            O => \N__15507\,
            I => \N__15504\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__15504\,
            I => rgb_c_3
        );

    \I__2306\ : InMux
    port map (
            O => \N__15501\,
            I => \N__15498\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__15498\,
            I => \N__15495\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__15495\,
            I => \N__15492\
        );

    \I__2303\ : Span4Mux_h
    port map (
            O => \N__15492\,
            I => \N__15489\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__15489\,
            I => \N_95_0\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__15486\,
            I => \N__15482\
        );

    \I__2300\ : InMux
    port map (
            O => \N__15485\,
            I => \N__15478\
        );

    \I__2299\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15475\
        );

    \I__2298\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15472\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__15478\,
            I => \N__15469\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__15475\,
            I => \N__15464\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__15472\,
            I => \N__15464\
        );

    \I__2294\ : Span4Mux_v
    port map (
            O => \N__15469\,
            I => \N__15458\
        );

    \I__2293\ : Span4Mux_v
    port map (
            O => \N__15464\,
            I => \N__15458\
        );

    \I__2292\ : InMux
    port map (
            O => \N__15463\,
            I => \N__15452\
        );

    \I__2291\ : Span4Mux_h
    port map (
            O => \N__15458\,
            I => \N__15449\
        );

    \I__2290\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15446\
        );

    \I__2289\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15443\
        );

    \I__2288\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15440\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__15452\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__15449\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__15446\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__15443\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__15440\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2282\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15426\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__15426\,
            I => \N__15422\
        );

    \I__2280\ : InMux
    port map (
            O => \N__15425\,
            I => \N__15418\
        );

    \I__2279\ : Span4Mux_h
    port map (
            O => \N__15422\,
            I => \N__15415\
        );

    \I__2278\ : InMux
    port map (
            O => \N__15421\,
            I => \N__15412\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__15418\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__15415\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__15412\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2274\ : InMux
    port map (
            O => \N__15405\,
            I => \N__15400\
        );

    \I__2273\ : InMux
    port map (
            O => \N__15404\,
            I => \N__15397\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__15403\,
            I => \N__15388\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__15400\,
            I => \N__15382\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__15397\,
            I => \N__15382\
        );

    \I__2269\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15379\
        );

    \I__2268\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15374\
        );

    \I__2267\ : InMux
    port map (
            O => \N__15394\,
            I => \N__15374\
        );

    \I__2266\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15371\
        );

    \I__2265\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15366\
        );

    \I__2264\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15366\
        );

    \I__2263\ : InMux
    port map (
            O => \N__15388\,
            I => \N__15362\
        );

    \I__2262\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15357\
        );

    \I__2261\ : Span4Mux_v
    port map (
            O => \N__15382\,
            I => \N__15352\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__15379\,
            I => \N__15352\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__15374\,
            I => \N__15347\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__15371\,
            I => \N__15347\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__15366\,
            I => \N__15344\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__15365\,
            I => \N__15341\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__15362\,
            I => \N__15338\
        );

    \I__2254\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15335\
        );

    \I__2253\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15332\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__15357\,
            I => \N__15325\
        );

    \I__2251\ : Span4Mux_h
    port map (
            O => \N__15352\,
            I => \N__15325\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__15347\,
            I => \N__15325\
        );

    \I__2249\ : Span12Mux_h
    port map (
            O => \N__15344\,
            I => \N__15322\
        );

    \I__2248\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15319\
        );

    \I__2247\ : Odrv12
    port map (
            O => \N__15338\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__15335\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__15332\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__15325\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2243\ : Odrv12
    port map (
            O => \N__15322\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__15319\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__15306\,
            I => \N__15303\
        );

    \I__2240\ : InMux
    port map (
            O => \N__15303\,
            I => \N__15299\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__15302\,
            I => \N__15292\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__15299\,
            I => \N__15288\
        );

    \I__2237\ : InMux
    port map (
            O => \N__15298\,
            I => \N__15283\
        );

    \I__2236\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15283\
        );

    \I__2235\ : InMux
    port map (
            O => \N__15296\,
            I => \N__15279\
        );

    \I__2234\ : InMux
    port map (
            O => \N__15295\,
            I => \N__15276\
        );

    \I__2233\ : InMux
    port map (
            O => \N__15292\,
            I => \N__15268\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__15291\,
            I => \N__15264\
        );

    \I__2231\ : Span4Mux_v
    port map (
            O => \N__15288\,
            I => \N__15258\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__15283\,
            I => \N__15258\
        );

    \I__2229\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15255\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__15279\,
            I => \N__15250\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__15276\,
            I => \N__15250\
        );

    \I__2226\ : InMux
    port map (
            O => \N__15275\,
            I => \N__15247\
        );

    \I__2225\ : InMux
    port map (
            O => \N__15274\,
            I => \N__15242\
        );

    \I__2224\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15242\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__15272\,
            I => \N__15237\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__15271\,
            I => \N__15231\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__15268\,
            I => \N__15227\
        );

    \I__2220\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15222\
        );

    \I__2219\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15217\
        );

    \I__2218\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15217\
        );

    \I__2217\ : Span4Mux_h
    port map (
            O => \N__15258\,
            I => \N__15214\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__15255\,
            I => \N__15205\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__15250\,
            I => \N__15205\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__15247\,
            I => \N__15205\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__15242\,
            I => \N__15205\
        );

    \I__2212\ : InMux
    port map (
            O => \N__15241\,
            I => \N__15198\
        );

    \I__2211\ : InMux
    port map (
            O => \N__15240\,
            I => \N__15198\
        );

    \I__2210\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15198\
        );

    \I__2209\ : InMux
    port map (
            O => \N__15236\,
            I => \N__15194\
        );

    \I__2208\ : InMux
    port map (
            O => \N__15235\,
            I => \N__15185\
        );

    \I__2207\ : InMux
    port map (
            O => \N__15234\,
            I => \N__15185\
        );

    \I__2206\ : InMux
    port map (
            O => \N__15231\,
            I => \N__15185\
        );

    \I__2205\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15185\
        );

    \I__2204\ : Span4Mux_v
    port map (
            O => \N__15227\,
            I => \N__15182\
        );

    \I__2203\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15177\
        );

    \I__2202\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15177\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__15222\,
            I => \N__15166\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__15217\,
            I => \N__15166\
        );

    \I__2199\ : Span4Mux_h
    port map (
            O => \N__15214\,
            I => \N__15166\
        );

    \I__2198\ : Span4Mux_h
    port map (
            O => \N__15205\,
            I => \N__15166\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__15198\,
            I => \N__15166\
        );

    \I__2196\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15163\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__15194\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__15185\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__15182\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__15177\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__15166\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__15163\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2189\ : InMux
    port map (
            O => \N__15150\,
            I => \N__15147\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__15147\,
            I => \N__15144\
        );

    \I__2187\ : Span4Mux_h
    port map (
            O => \N__15144\,
            I => \N__15141\
        );

    \I__2186\ : Span4Mux_v
    port map (
            O => \N__15141\,
            I => \N__15138\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__15138\,
            I => \N__15135\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__15135\,
            I => \M_this_map_ram_read_data_2\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__15132\,
            I => \N__15129\
        );

    \I__2182\ : InMux
    port map (
            O => \N__15129\,
            I => \N__15122\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__15128\,
            I => \N__15119\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__15127\,
            I => \N__15114\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__15126\,
            I => \N__15111\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__15125\,
            I => \N__15108\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__15122\,
            I => \N__15103\
        );

    \I__2176\ : InMux
    port map (
            O => \N__15119\,
            I => \N__15100\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__15118\,
            I => \N__15097\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__15117\,
            I => \N__15094\
        );

    \I__2173\ : InMux
    port map (
            O => \N__15114\,
            I => \N__15089\
        );

    \I__2172\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15085\
        );

    \I__2171\ : InMux
    port map (
            O => \N__15108\,
            I => \N__15082\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__15107\,
            I => \N__15079\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__15106\,
            I => \N__15076\
        );

    \I__2168\ : Span4Mux_h
    port map (
            O => \N__15103\,
            I => \N__15070\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__15100\,
            I => \N__15070\
        );

    \I__2166\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15067\
        );

    \I__2165\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15064\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__15093\,
            I => \N__15061\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__15092\,
            I => \N__15058\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__15089\,
            I => \N__15053\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__15088\,
            I => \N__15050\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__15085\,
            I => \N__15045\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__15082\,
            I => \N__15045\
        );

    \I__2158\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15042\
        );

    \I__2157\ : InMux
    port map (
            O => \N__15076\,
            I => \N__15039\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__15075\,
            I => \N__15035\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__15070\,
            I => \N__15030\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__15067\,
            I => \N__15030\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__15064\,
            I => \N__15027\
        );

    \I__2152\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15024\
        );

    \I__2151\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15021\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__15057\,
            I => \N__15018\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__15056\,
            I => \N__15015\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__15053\,
            I => \N__15012\
        );

    \I__2147\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15009\
        );

    \I__2146\ : Span4Mux_v
    port map (
            O => \N__15045\,
            I => \N__15002\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__15042\,
            I => \N__15002\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__15039\,
            I => \N__15002\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__15038\,
            I => \N__14999\
        );

    \I__2142\ : InMux
    port map (
            O => \N__15035\,
            I => \N__14996\
        );

    \I__2141\ : Span4Mux_h
    port map (
            O => \N__15030\,
            I => \N__14993\
        );

    \I__2140\ : Span4Mux_v
    port map (
            O => \N__15027\,
            I => \N__14988\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__15024\,
            I => \N__14988\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__15021\,
            I => \N__14985\
        );

    \I__2137\ : InMux
    port map (
            O => \N__15018\,
            I => \N__14982\
        );

    \I__2136\ : InMux
    port map (
            O => \N__15015\,
            I => \N__14979\
        );

    \I__2135\ : Sp12to4
    port map (
            O => \N__15012\,
            I => \N__14974\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__15009\,
            I => \N__14974\
        );

    \I__2133\ : Span4Mux_v
    port map (
            O => \N__15002\,
            I => \N__14971\
        );

    \I__2132\ : InMux
    port map (
            O => \N__14999\,
            I => \N__14968\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__14996\,
            I => \N__14965\
        );

    \I__2130\ : Span4Mux_v
    port map (
            O => \N__14993\,
            I => \N__14960\
        );

    \I__2129\ : Span4Mux_h
    port map (
            O => \N__14988\,
            I => \N__14960\
        );

    \I__2128\ : Span4Mux_h
    port map (
            O => \N__14985\,
            I => \N__14957\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__14982\,
            I => \N__14954\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__14979\,
            I => \N__14951\
        );

    \I__2125\ : Span12Mux_h
    port map (
            O => \N__14974\,
            I => \N__14948\
        );

    \I__2124\ : Sp12to4
    port map (
            O => \N__14971\,
            I => \N__14943\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__14968\,
            I => \N__14943\
        );

    \I__2122\ : Span4Mux_h
    port map (
            O => \N__14965\,
            I => \N__14940\
        );

    \I__2121\ : Span4Mux_h
    port map (
            O => \N__14960\,
            I => \N__14937\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__14957\,
            I => \N__14932\
        );

    \I__2119\ : Span4Mux_h
    port map (
            O => \N__14954\,
            I => \N__14932\
        );

    \I__2118\ : Span4Mux_h
    port map (
            O => \N__14951\,
            I => \N__14929\
        );

    \I__2117\ : Span12Mux_v
    port map (
            O => \N__14948\,
            I => \N__14926\
        );

    \I__2116\ : Span12Mux_h
    port map (
            O => \N__14943\,
            I => \N__14923\
        );

    \I__2115\ : Span4Mux_v
    port map (
            O => \N__14940\,
            I => \N__14920\
        );

    \I__2114\ : Span4Mux_h
    port map (
            O => \N__14937\,
            I => \N__14913\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__14932\,
            I => \N__14913\
        );

    \I__2112\ : Span4Mux_h
    port map (
            O => \N__14929\,
            I => \N__14913\
        );

    \I__2111\ : Odrv12
    port map (
            O => \N__14926\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__2110\ : Odrv12
    port map (
            O => \N__14923\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__14920\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__14913\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__2107\ : InMux
    port map (
            O => \N__14904\,
            I => \N__14901\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__14901\,
            I => \this_vga_ramdac.N_24_mux\
        );

    \I__2105\ : InMux
    port map (
            O => \N__14898\,
            I => \N__14895\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__14895\,
            I => \N__14892\
        );

    \I__2103\ : Span4Mux_h
    port map (
            O => \N__14892\,
            I => \N__14888\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__14891\,
            I => \N__14885\
        );

    \I__2101\ : Span4Mux_h
    port map (
            O => \N__14888\,
            I => \N__14882\
        );

    \I__2100\ : InMux
    port map (
            O => \N__14885\,
            I => \N__14879\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__14882\,
            I => \this_vga_ramdac.N_2862_reto\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__14879\,
            I => \this_vga_ramdac.N_2862_reto\
        );

    \I__2097\ : InMux
    port map (
            O => \N__14874\,
            I => \bfn_13_18_0_\
        );

    \I__2096\ : InMux
    port map (
            O => \N__14871\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__2095\ : InMux
    port map (
            O => \N__14868\,
            I => \N__14863\
        );

    \I__2094\ : InMux
    port map (
            O => \N__14867\,
            I => \N__14860\
        );

    \I__2093\ : InMux
    port map (
            O => \N__14866\,
            I => \N__14857\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__14863\,
            I => \N__14852\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__14860\,
            I => \N__14852\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__14857\,
            I => \N__14849\
        );

    \I__2089\ : Span4Mux_v
    port map (
            O => \N__14852\,
            I => \N__14846\
        );

    \I__2088\ : Span4Mux_h
    port map (
            O => \N__14849\,
            I => \N__14843\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__14846\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__14843\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__2085\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14834\
        );

    \I__2084\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14831\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__14834\,
            I => \N__14826\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__14831\,
            I => \N__14826\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__14826\,
            I => \N__14822\
        );

    \I__2080\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14819\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__14822\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__14819\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__14814\,
            I => \N__14810\
        );

    \I__2076\ : InMux
    port map (
            O => \N__14813\,
            I => \N__14807\
        );

    \I__2075\ : InMux
    port map (
            O => \N__14810\,
            I => \N__14804\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__14807\,
            I => \N__14799\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__14804\,
            I => \N__14799\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__14799\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__2071\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14792\
        );

    \I__2070\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14788\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__14792\,
            I => \N__14785\
        );

    \I__2068\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14782\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__14788\,
            I => \N__14779\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__14785\,
            I => \N__14774\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__14782\,
            I => \N__14774\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__14779\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__14774\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2062\ : CEMux
    port map (
            O => \N__14769\,
            I => \N__14742\
        );

    \I__2061\ : CEMux
    port map (
            O => \N__14768\,
            I => \N__14742\
        );

    \I__2060\ : CEMux
    port map (
            O => \N__14767\,
            I => \N__14742\
        );

    \I__2059\ : CEMux
    port map (
            O => \N__14766\,
            I => \N__14742\
        );

    \I__2058\ : CEMux
    port map (
            O => \N__14765\,
            I => \N__14742\
        );

    \I__2057\ : CEMux
    port map (
            O => \N__14764\,
            I => \N__14742\
        );

    \I__2056\ : CEMux
    port map (
            O => \N__14763\,
            I => \N__14742\
        );

    \I__2055\ : CEMux
    port map (
            O => \N__14762\,
            I => \N__14742\
        );

    \I__2054\ : CEMux
    port map (
            O => \N__14761\,
            I => \N__14742\
        );

    \I__2053\ : GlobalMux
    port map (
            O => \N__14742\,
            I => \N__14739\
        );

    \I__2052\ : gio2CtrlBuf
    port map (
            O => \N__14739\,
            I => \this_vga_signals.N_692_0_g\
        );

    \I__2051\ : InMux
    port map (
            O => \N__14736\,
            I => \N__14733\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__14733\,
            I => \N__14720\
        );

    \I__2049\ : SRMux
    port map (
            O => \N__14732\,
            I => \N__14697\
        );

    \I__2048\ : SRMux
    port map (
            O => \N__14731\,
            I => \N__14697\
        );

    \I__2047\ : SRMux
    port map (
            O => \N__14730\,
            I => \N__14697\
        );

    \I__2046\ : SRMux
    port map (
            O => \N__14729\,
            I => \N__14697\
        );

    \I__2045\ : SRMux
    port map (
            O => \N__14728\,
            I => \N__14697\
        );

    \I__2044\ : SRMux
    port map (
            O => \N__14727\,
            I => \N__14697\
        );

    \I__2043\ : SRMux
    port map (
            O => \N__14726\,
            I => \N__14697\
        );

    \I__2042\ : SRMux
    port map (
            O => \N__14725\,
            I => \N__14697\
        );

    \I__2041\ : SRMux
    port map (
            O => \N__14724\,
            I => \N__14697\
        );

    \I__2040\ : SRMux
    port map (
            O => \N__14723\,
            I => \N__14697\
        );

    \I__2039\ : Glb2LocalMux
    port map (
            O => \N__14720\,
            I => \N__14697\
        );

    \I__2038\ : GlobalMux
    port map (
            O => \N__14697\,
            I => \N__14694\
        );

    \I__2037\ : gio2CtrlBuf
    port map (
            O => \N__14694\,
            I => \this_vga_signals.N_988_g\
        );

    \I__2036\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14687\
        );

    \I__2035\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14684\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__14687\,
            I => \N__14681\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14675\
        );

    \I__2032\ : Span4Mux_h
    port map (
            O => \N__14681\,
            I => \N__14672\
        );

    \I__2031\ : InMux
    port map (
            O => \N__14680\,
            I => \N__14666\
        );

    \I__2030\ : InMux
    port map (
            O => \N__14679\,
            I => \N__14666\
        );

    \I__2029\ : InMux
    port map (
            O => \N__14678\,
            I => \N__14660\
        );

    \I__2028\ : Span4Mux_h
    port map (
            O => \N__14675\,
            I => \N__14655\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__14672\,
            I => \N__14655\
        );

    \I__2026\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14652\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__14666\,
            I => \N__14649\
        );

    \I__2024\ : InMux
    port map (
            O => \N__14665\,
            I => \N__14642\
        );

    \I__2023\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14642\
        );

    \I__2022\ : InMux
    port map (
            O => \N__14663\,
            I => \N__14642\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__14660\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__14655\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__14652\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__14649\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__14642\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2016\ : InMux
    port map (
            O => \N__14631\,
            I => \N__14628\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__14628\,
            I => \N__14625\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__14625\,
            I => \this_vga_signals.un4_hsynclt8_0\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__14622\,
            I => \N__14619\
        );

    \I__2012\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14616\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__14616\,
            I => \N__14613\
        );

    \I__2010\ : Span4Mux_h
    port map (
            O => \N__14613\,
            I => \N__14610\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__14610\,
            I => \this_vga_signals.un2_hsynclt8_0\
        );

    \I__2008\ : InMux
    port map (
            O => \N__14607\,
            I => \N__14603\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__14606\,
            I => \N__14598\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__14603\,
            I => \N__14593\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__14602\,
            I => \N__14588\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__14601\,
            I => \N__14584\
        );

    \I__2003\ : InMux
    port map (
            O => \N__14598\,
            I => \N__14581\
        );

    \I__2002\ : InMux
    port map (
            O => \N__14597\,
            I => \N__14578\
        );

    \I__2001\ : InMux
    port map (
            O => \N__14596\,
            I => \N__14575\
        );

    \I__2000\ : Span4Mux_v
    port map (
            O => \N__14593\,
            I => \N__14572\
        );

    \I__1999\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14569\
        );

    \I__1998\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14566\
        );

    \I__1997\ : InMux
    port map (
            O => \N__14588\,
            I => \N__14559\
        );

    \I__1996\ : InMux
    port map (
            O => \N__14587\,
            I => \N__14559\
        );

    \I__1995\ : InMux
    port map (
            O => \N__14584\,
            I => \N__14559\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__14581\,
            I => \N__14552\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__14578\,
            I => \N__14552\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__14575\,
            I => \N__14552\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__14572\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__14569\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__14566\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__14559\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__14552\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1986\ : IoInMux
    port map (
            O => \N__14541\,
            I => \N__14538\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__14538\,
            I => \N__14535\
        );

    \I__1984\ : Span4Mux_s3_v
    port map (
            O => \N__14535\,
            I => \N__14532\
        );

    \I__1983\ : Sp12to4
    port map (
            O => \N__14532\,
            I => \N__14529\
        );

    \I__1982\ : Span12Mux_h
    port map (
            O => \N__14529\,
            I => \N__14526\
        );

    \I__1981\ : Odrv12
    port map (
            O => \N__14526\,
            I => this_vga_signals_hsync_1_i
        );

    \I__1980\ : InMux
    port map (
            O => \N__14523\,
            I => \N__14520\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__14520\,
            I => \N__14517\
        );

    \I__1978\ : Span4Mux_h
    port map (
            O => \N__14517\,
            I => \N__14514\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__14514\,
            I => \N__14511\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__14511\,
            I => \N__14508\
        );

    \I__1975\ : Span4Mux_h
    port map (
            O => \N__14508\,
            I => \N__14505\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__14505\,
            I => \M_this_map_ram_read_data_0\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__14502\,
            I => \N__14497\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__14501\,
            I => \N__14491\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__14500\,
            I => \N__14484\
        );

    \I__1970\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14480\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__14496\,
            I => \N__14477\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__14495\,
            I => \N__14474\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__14494\,
            I => \N__14471\
        );

    \I__1966\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14466\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__14490\,
            I => \N__14461\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__14489\,
            I => \N__14457\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__14488\,
            I => \N__14454\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__14487\,
            I => \N__14451\
        );

    \I__1961\ : InMux
    port map (
            O => \N__14484\,
            I => \N__14448\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__14483\,
            I => \N__14445\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__14480\,
            I => \N__14442\
        );

    \I__1958\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14439\
        );

    \I__1957\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14436\
        );

    \I__1956\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14433\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__14470\,
            I => \N__14430\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__14469\,
            I => \N__14427\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__14466\,
            I => \N__14424\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__14465\,
            I => \N__14421\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__14464\,
            I => \N__14418\
        );

    \I__1950\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14415\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__14460\,
            I => \N__14412\
        );

    \I__1948\ : InMux
    port map (
            O => \N__14457\,
            I => \N__14409\
        );

    \I__1947\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14406\
        );

    \I__1946\ : InMux
    port map (
            O => \N__14451\,
            I => \N__14403\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__14448\,
            I => \N__14400\
        );

    \I__1944\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14397\
        );

    \I__1943\ : Span4Mux_h
    port map (
            O => \N__14442\,
            I => \N__14394\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__14439\,
            I => \N__14391\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__14436\,
            I => \N__14386\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__14433\,
            I => \N__14386\
        );

    \I__1939\ : InMux
    port map (
            O => \N__14430\,
            I => \N__14383\
        );

    \I__1938\ : InMux
    port map (
            O => \N__14427\,
            I => \N__14380\
        );

    \I__1937\ : Span4Mux_v
    port map (
            O => \N__14424\,
            I => \N__14377\
        );

    \I__1936\ : InMux
    port map (
            O => \N__14421\,
            I => \N__14374\
        );

    \I__1935\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14371\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__14415\,
            I => \N__14368\
        );

    \I__1933\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14365\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__14409\,
            I => \N__14362\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__14406\,
            I => \N__14359\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__14403\,
            I => \N__14356\
        );

    \I__1929\ : Span4Mux_v
    port map (
            O => \N__14400\,
            I => \N__14351\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__14397\,
            I => \N__14351\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__14394\,
            I => \N__14348\
        );

    \I__1926\ : Span4Mux_v
    port map (
            O => \N__14391\,
            I => \N__14341\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__14386\,
            I => \N__14341\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__14383\,
            I => \N__14341\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__14380\,
            I => \N__14338\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__14377\,
            I => \N__14335\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__14374\,
            I => \N__14328\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__14371\,
            I => \N__14328\
        );

    \I__1919\ : Sp12to4
    port map (
            O => \N__14368\,
            I => \N__14328\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__14365\,
            I => \N__14325\
        );

    \I__1917\ : Span12Mux_h
    port map (
            O => \N__14362\,
            I => \N__14322\
        );

    \I__1916\ : Span4Mux_v
    port map (
            O => \N__14359\,
            I => \N__14319\
        );

    \I__1915\ : Span4Mux_v
    port map (
            O => \N__14356\,
            I => \N__14314\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__14351\,
            I => \N__14314\
        );

    \I__1913\ : Sp12to4
    port map (
            O => \N__14348\,
            I => \N__14309\
        );

    \I__1912\ : Sp12to4
    port map (
            O => \N__14341\,
            I => \N__14309\
        );

    \I__1911\ : Sp12to4
    port map (
            O => \N__14338\,
            I => \N__14302\
        );

    \I__1910\ : Sp12to4
    port map (
            O => \N__14335\,
            I => \N__14302\
        );

    \I__1909\ : Span12Mux_s11_v
    port map (
            O => \N__14328\,
            I => \N__14302\
        );

    \I__1908\ : Span12Mux_s9_h
    port map (
            O => \N__14325\,
            I => \N__14299\
        );

    \I__1907\ : Span12Mux_v
    port map (
            O => \N__14322\,
            I => \N__14296\
        );

    \I__1906\ : Span4Mux_h
    port map (
            O => \N__14319\,
            I => \N__14291\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__14314\,
            I => \N__14291\
        );

    \I__1904\ : Span12Mux_h
    port map (
            O => \N__14309\,
            I => \N__14286\
        );

    \I__1903\ : Span12Mux_h
    port map (
            O => \N__14302\,
            I => \N__14286\
        );

    \I__1902\ : Odrv12
    port map (
            O => \N__14299\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__1901\ : Odrv12
    port map (
            O => \N__14296\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__14291\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__1899\ : Odrv12
    port map (
            O => \N__14286\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__1898\ : InMux
    port map (
            O => \N__14277\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__1897\ : InMux
    port map (
            O => \N__14274\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__1896\ : InMux
    port map (
            O => \N__14271\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__1895\ : InMux
    port map (
            O => \N__14268\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__1894\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14259\
        );

    \I__1893\ : InMux
    port map (
            O => \N__14264\,
            I => \N__14259\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__14259\,
            I => \N__14255\
        );

    \I__1891\ : InMux
    port map (
            O => \N__14258\,
            I => \N__14252\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__14255\,
            I => \N__14247\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__14252\,
            I => \N__14247\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__14247\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__1887\ : InMux
    port map (
            O => \N__14244\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__1886\ : InMux
    port map (
            O => \N__14241\,
            I => \N__14237\
        );

    \I__1885\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14234\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__14237\,
            I => \N__14230\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__14234\,
            I => \N__14227\
        );

    \I__1882\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14224\
        );

    \I__1881\ : Span4Mux_h
    port map (
            O => \N__14230\,
            I => \N__14221\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__14227\,
            I => \N__14218\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__14224\,
            I => \N__14215\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__14221\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__14218\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1876\ : Odrv12
    port map (
            O => \N__14215\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1875\ : InMux
    port map (
            O => \N__14208\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__1874\ : InMux
    port map (
            O => \N__14205\,
            I => \N__14202\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__14202\,
            I => \N__14198\
        );

    \I__1872\ : InMux
    port map (
            O => \N__14201\,
            I => \N__14195\
        );

    \I__1871\ : Span4Mux_h
    port map (
            O => \N__14198\,
            I => \N__14192\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__14195\,
            I => \N__14189\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__14192\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__1868\ : Odrv12
    port map (
            O => \N__14189\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__1867\ : InMux
    port map (
            O => \N__14184\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__14181\,
            I => \N__14178\
        );

    \I__1865\ : InMux
    port map (
            O => \N__14178\,
            I => \N__14175\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__14175\,
            I => \N__14168\
        );

    \I__1863\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14165\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__14173\,
            I => \N__14161\
        );

    \I__1861\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14155\
        );

    \I__1860\ : InMux
    port map (
            O => \N__14171\,
            I => \N__14152\
        );

    \I__1859\ : Span4Mux_h
    port map (
            O => \N__14168\,
            I => \N__14149\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__14165\,
            I => \N__14146\
        );

    \I__1857\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14139\
        );

    \I__1856\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14139\
        );

    \I__1855\ : InMux
    port map (
            O => \N__14160\,
            I => \N__14139\
        );

    \I__1854\ : InMux
    port map (
            O => \N__14159\,
            I => \N__14134\
        );

    \I__1853\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14134\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__14155\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__14152\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__14149\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__14146\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__14139\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__14134\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1846\ : InMux
    port map (
            O => \N__14121\,
            I => \N__14115\
        );

    \I__1845\ : InMux
    port map (
            O => \N__14120\,
            I => \N__14115\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__14115\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__14112\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_\
        );

    \I__1842\ : InMux
    port map (
            O => \N__14109\,
            I => \N__14106\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__14106\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0_0_0\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__14103\,
            I => \N__14097\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__14102\,
            I => \N__14094\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__14101\,
            I => \N__14090\
        );

    \I__1837\ : InMux
    port map (
            O => \N__14100\,
            I => \N__14084\
        );

    \I__1836\ : InMux
    port map (
            O => \N__14097\,
            I => \N__14079\
        );

    \I__1835\ : InMux
    port map (
            O => \N__14094\,
            I => \N__14079\
        );

    \I__1834\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14074\
        );

    \I__1833\ : InMux
    port map (
            O => \N__14090\,
            I => \N__14074\
        );

    \I__1832\ : InMux
    port map (
            O => \N__14089\,
            I => \N__14070\
        );

    \I__1831\ : InMux
    port map (
            O => \N__14088\,
            I => \N__14067\
        );

    \I__1830\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14064\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__14084\,
            I => \N__14057\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__14079\,
            I => \N__14057\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__14074\,
            I => \N__14057\
        );

    \I__1826\ : InMux
    port map (
            O => \N__14073\,
            I => \N__14054\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__14070\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__14067\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__14064\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__14057\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__14054\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1820\ : InMux
    port map (
            O => \N__14043\,
            I => \N__14033\
        );

    \I__1819\ : InMux
    port map (
            O => \N__14042\,
            I => \N__14033\
        );

    \I__1818\ : InMux
    port map (
            O => \N__14041\,
            I => \N__14028\
        );

    \I__1817\ : InMux
    port map (
            O => \N__14040\,
            I => \N__14028\
        );

    \I__1816\ : InMux
    port map (
            O => \N__14039\,
            I => \N__14024\
        );

    \I__1815\ : InMux
    port map (
            O => \N__14038\,
            I => \N__14021\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__14033\,
            I => \N__14018\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__14028\,
            I => \N__14015\
        );

    \I__1812\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14012\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__14024\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__14021\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__14018\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__14015\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__14012\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1806\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13995\
        );

    \I__1805\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13991\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__13999\,
            I => \N__13987\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__13998\,
            I => \N__13984\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__13995\,
            I => \N__13981\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__13994\,
            I => \N__13977\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__13991\,
            I => \N__13974\
        );

    \I__1799\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13971\
        );

    \I__1798\ : InMux
    port map (
            O => \N__13987\,
            I => \N__13966\
        );

    \I__1797\ : InMux
    port map (
            O => \N__13984\,
            I => \N__13966\
        );

    \I__1796\ : Span4Mux_v
    port map (
            O => \N__13981\,
            I => \N__13963\
        );

    \I__1795\ : InMux
    port map (
            O => \N__13980\,
            I => \N__13960\
        );

    \I__1794\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13957\
        );

    \I__1793\ : Span4Mux_h
    port map (
            O => \N__13974\,
            I => \N__13954\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__13971\,
            I => \N__13949\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__13966\,
            I => \N__13949\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__13963\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__13960\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__13957\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__13954\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__13949\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1785\ : InMux
    port map (
            O => \N__13938\,
            I => \N__13934\
        );

    \I__1784\ : InMux
    port map (
            O => \N__13937\,
            I => \N__13921\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__13934\,
            I => \N__13918\
        );

    \I__1782\ : InMux
    port map (
            O => \N__13933\,
            I => \N__13913\
        );

    \I__1781\ : InMux
    port map (
            O => \N__13932\,
            I => \N__13913\
        );

    \I__1780\ : InMux
    port map (
            O => \N__13931\,
            I => \N__13908\
        );

    \I__1779\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13908\
        );

    \I__1778\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13895\
        );

    \I__1777\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13895\
        );

    \I__1776\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13895\
        );

    \I__1775\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13895\
        );

    \I__1774\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13895\
        );

    \I__1773\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13895\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__13921\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__13918\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__13913\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__13908\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__13895\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__13884\,
            I => \N__13874\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__13883\,
            I => \N__13871\
        );

    \I__1765\ : InMux
    port map (
            O => \N__13882\,
            I => \N__13866\
        );

    \I__1764\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13861\
        );

    \I__1763\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13861\
        );

    \I__1762\ : InMux
    port map (
            O => \N__13879\,
            I => \N__13858\
        );

    \I__1761\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13849\
        );

    \I__1760\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13849\
        );

    \I__1759\ : InMux
    port map (
            O => \N__13874\,
            I => \N__13849\
        );

    \I__1758\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13849\
        );

    \I__1757\ : InMux
    port map (
            O => \N__13870\,
            I => \N__13844\
        );

    \I__1756\ : InMux
    port map (
            O => \N__13869\,
            I => \N__13844\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__13866\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__13861\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__13858\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__13849\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__13844\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__13833\,
            I => \this_vga_signals.un4_hsynclt4_0_cascade_\
        );

    \I__1749\ : InMux
    port map (
            O => \N__13830\,
            I => \N__13821\
        );

    \I__1748\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13816\
        );

    \I__1747\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13816\
        );

    \I__1746\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13811\
        );

    \I__1745\ : InMux
    port map (
            O => \N__13826\,
            I => \N__13811\
        );

    \I__1744\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13802\
        );

    \I__1743\ : InMux
    port map (
            O => \N__13824\,
            I => \N__13799\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__13821\,
            I => \N__13796\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__13816\,
            I => \N__13793\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__13811\,
            I => \N__13790\
        );

    \I__1739\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13783\
        );

    \I__1738\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13783\
        );

    \I__1737\ : InMux
    port map (
            O => \N__13808\,
            I => \N__13783\
        );

    \I__1736\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13776\
        );

    \I__1735\ : InMux
    port map (
            O => \N__13806\,
            I => \N__13776\
        );

    \I__1734\ : InMux
    port map (
            O => \N__13805\,
            I => \N__13776\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__13802\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__13799\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__13796\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1730\ : Odrv4
    port map (
            O => \N__13793\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__13790\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__13783\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__13776\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1726\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13758\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__13758\,
            I => \N__13755\
        );

    \I__1724\ : Odrv12
    port map (
            O => \N__13755\,
            I => \N_91_0\
        );

    \I__1723\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13749\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__13749\,
            I => \N__13746\
        );

    \I__1721\ : Span4Mux_h
    port map (
            O => \N__13746\,
            I => \N__13743\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__13743\,
            I => \N_93_0\
        );

    \I__1719\ : InMux
    port map (
            O => \N__13740\,
            I => \N__13737\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__13737\,
            I => \N__13734\
        );

    \I__1717\ : Sp12to4
    port map (
            O => \N__13734\,
            I => \N__13731\
        );

    \I__1716\ : Span12Mux_v
    port map (
            O => \N__13731\,
            I => \N__13728\
        );

    \I__1715\ : Odrv12
    port map (
            O => \N__13728\,
            I => \M_this_map_ram_read_data_3\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__13725\,
            I => \N__13721\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__13724\,
            I => \N__13718\
        );

    \I__1712\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13712\
        );

    \I__1711\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13708\
        );

    \I__1710\ : CascadeMux
    port map (
            O => \N__13717\,
            I => \N__13705\
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__13716\,
            I => \N__13701\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__13715\,
            I => \N__13697\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__13712\,
            I => \N__13692\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__13711\,
            I => \N__13689\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__13708\,
            I => \N__13685\
        );

    \I__1704\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13682\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__13704\,
            I => \N__13679\
        );

    \I__1702\ : InMux
    port map (
            O => \N__13701\,
            I => \N__13675\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__13700\,
            I => \N__13672\
        );

    \I__1700\ : InMux
    port map (
            O => \N__13697\,
            I => \N__13667\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__13696\,
            I => \N__13664\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__13695\,
            I => \N__13661\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__13692\,
            I => \N__13658\
        );

    \I__1696\ : InMux
    port map (
            O => \N__13689\,
            I => \N__13655\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__13688\,
            I => \N__13652\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__13685\,
            I => \N__13647\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__13682\,
            I => \N__13647\
        );

    \I__1692\ : InMux
    port map (
            O => \N__13679\,
            I => \N__13644\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__13678\,
            I => \N__13641\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__13675\,
            I => \N__13638\
        );

    \I__1689\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13635\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__13671\,
            I => \N__13632\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__13670\,
            I => \N__13628\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__13667\,
            I => \N__13625\
        );

    \I__1685\ : InMux
    port map (
            O => \N__13664\,
            I => \N__13622\
        );

    \I__1684\ : InMux
    port map (
            O => \N__13661\,
            I => \N__13619\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__13658\,
            I => \N__13616\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__13655\,
            I => \N__13613\
        );

    \I__1681\ : InMux
    port map (
            O => \N__13652\,
            I => \N__13610\
        );

    \I__1680\ : Span4Mux_h
    port map (
            O => \N__13647\,
            I => \N__13605\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__13644\,
            I => \N__13605\
        );

    \I__1678\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13602\
        );

    \I__1677\ : Span4Mux_h
    port map (
            O => \N__13638\,
            I => \N__13596\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__13635\,
            I => \N__13596\
        );

    \I__1675\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13593\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__13631\,
            I => \N__13590\
        );

    \I__1673\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13587\
        );

    \I__1672\ : Span4Mux_h
    port map (
            O => \N__13625\,
            I => \N__13584\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__13622\,
            I => \N__13581\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__13619\,
            I => \N__13578\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__13616\,
            I => \N__13571\
        );

    \I__1668\ : Span4Mux_v
    port map (
            O => \N__13613\,
            I => \N__13571\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__13610\,
            I => \N__13571\
        );

    \I__1666\ : Span4Mux_v
    port map (
            O => \N__13605\,
            I => \N__13566\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__13602\,
            I => \N__13566\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__13601\,
            I => \N__13563\
        );

    \I__1663\ : Span4Mux_v
    port map (
            O => \N__13596\,
            I => \N__13558\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__13593\,
            I => \N__13558\
        );

    \I__1661\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13555\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__13587\,
            I => \N__13552\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__13584\,
            I => \N__13547\
        );

    \I__1658\ : Span4Mux_h
    port map (
            O => \N__13581\,
            I => \N__13547\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__13578\,
            I => \N__13544\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__13571\,
            I => \N__13539\
        );

    \I__1655\ : Span4Mux_v
    port map (
            O => \N__13566\,
            I => \N__13539\
        );

    \I__1654\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13536\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__13558\,
            I => \N__13531\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__13555\,
            I => \N__13531\
        );

    \I__1651\ : Span12Mux_s9_h
    port map (
            O => \N__13552\,
            I => \N__13526\
        );

    \I__1650\ : Sp12to4
    port map (
            O => \N__13547\,
            I => \N__13526\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__13544\,
            I => \N__13521\
        );

    \I__1648\ : Span4Mux_h
    port map (
            O => \N__13539\,
            I => \N__13521\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__13536\,
            I => \N__13518\
        );

    \I__1646\ : Span4Mux_h
    port map (
            O => \N__13531\,
            I => \N__13515\
        );

    \I__1645\ : Span12Mux_v
    port map (
            O => \N__13526\,
            I => \N__13508\
        );

    \I__1644\ : Sp12to4
    port map (
            O => \N__13521\,
            I => \N__13508\
        );

    \I__1643\ : Span12Mux_s9_h
    port map (
            O => \N__13518\,
            I => \N__13508\
        );

    \I__1642\ : Span4Mux_h
    port map (
            O => \N__13515\,
            I => \N__13505\
        );

    \I__1641\ : Odrv12
    port map (
            O => \N__13508\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__13505\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__13500\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__13497\,
            I => \N__13494\
        );

    \I__1637\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13485\
        );

    \I__1636\ : InMux
    port map (
            O => \N__13493\,
            I => \N__13485\
        );

    \I__1635\ : InMux
    port map (
            O => \N__13492\,
            I => \N__13485\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__13485\,
            I => \this_vga_signals.mult1_un68_sum_axb2_1\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__13482\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1_cascade_\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__13479\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_\
        );

    \I__1631\ : InMux
    port map (
            O => \N__13476\,
            I => \N__13473\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__13473\,
            I => \N__13470\
        );

    \I__1629\ : Span4Mux_h
    port map (
            O => \N__13470\,
            I => \N__13467\
        );

    \I__1628\ : Span4Mux_v
    port map (
            O => \N__13467\,
            I => \N__13460\
        );

    \I__1627\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13455\
        );

    \I__1626\ : InMux
    port map (
            O => \N__13465\,
            I => \N__13455\
        );

    \I__1625\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13450\
        );

    \I__1624\ : InMux
    port map (
            O => \N__13463\,
            I => \N__13450\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__13460\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__13455\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__13450\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__13443\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_\
        );

    \I__1619\ : InMux
    port map (
            O => \N__13440\,
            I => \N__13437\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__13437\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_0\
        );

    \I__1617\ : InMux
    port map (
            O => \N__13434\,
            I => \N__13431\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__13431\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__13428\,
            I => \N__13425\
        );

    \I__1614\ : InMux
    port map (
            O => \N__13425\,
            I => \N__13422\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__13422\,
            I => \N__13419\
        );

    \I__1612\ : Span12Mux_s11_h
    port map (
            O => \N__13419\,
            I => \N__13416\
        );

    \I__1611\ : Odrv12
    port map (
            O => \N__13416\,
            I => \M_this_vga_signals_address_5\
        );

    \I__1610\ : InMux
    port map (
            O => \N__13413\,
            I => \N__13407\
        );

    \I__1609\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13407\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__13407\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__13404\,
            I => \this_vga_signals.SUM_3_cascade_\
        );

    \I__1606\ : InMux
    port map (
            O => \N__13401\,
            I => \N__13398\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__13398\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0\
        );

    \I__1604\ : InMux
    port map (
            O => \N__13395\,
            I => \N__13392\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__13392\,
            I => \this_vga_signals.N_6_1\
        );

    \I__1602\ : InMux
    port map (
            O => \N__13389\,
            I => \N__13378\
        );

    \I__1601\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13378\
        );

    \I__1600\ : InMux
    port map (
            O => \N__13387\,
            I => \N__13370\
        );

    \I__1599\ : InMux
    port map (
            O => \N__13386\,
            I => \N__13370\
        );

    \I__1598\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13370\
        );

    \I__1597\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13358\
        );

    \I__1596\ : InMux
    port map (
            O => \N__13383\,
            I => \N__13355\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__13378\,
            I => \N__13352\
        );

    \I__1594\ : InMux
    port map (
            O => \N__13377\,
            I => \N__13349\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__13370\,
            I => \N__13346\
        );

    \I__1592\ : InMux
    port map (
            O => \N__13369\,
            I => \N__13339\
        );

    \I__1591\ : InMux
    port map (
            O => \N__13368\,
            I => \N__13339\
        );

    \I__1590\ : InMux
    port map (
            O => \N__13367\,
            I => \N__13339\
        );

    \I__1589\ : InMux
    port map (
            O => \N__13366\,
            I => \N__13332\
        );

    \I__1588\ : InMux
    port map (
            O => \N__13365\,
            I => \N__13332\
        );

    \I__1587\ : InMux
    port map (
            O => \N__13364\,
            I => \N__13332\
        );

    \I__1586\ : InMux
    port map (
            O => \N__13363\,
            I => \N__13325\
        );

    \I__1585\ : InMux
    port map (
            O => \N__13362\,
            I => \N__13325\
        );

    \I__1584\ : InMux
    port map (
            O => \N__13361\,
            I => \N__13325\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__13358\,
            I => \this_vga_signals.mult1_un68_sum_axb1_571\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__13355\,
            I => \this_vga_signals.mult1_un68_sum_axb1_571\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__13352\,
            I => \this_vga_signals.mult1_un68_sum_axb1_571\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__13349\,
            I => \this_vga_signals.mult1_un68_sum_axb1_571\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__13346\,
            I => \this_vga_signals.mult1_un68_sum_axb1_571\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__13339\,
            I => \this_vga_signals.mult1_un68_sum_axb1_571\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__13332\,
            I => \this_vga_signals.mult1_un68_sum_axb1_571\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__13325\,
            I => \this_vga_signals.mult1_un68_sum_axb1_571\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__13308\,
            I => \N__13303\
        );

    \I__1574\ : InMux
    port map (
            O => \N__13307\,
            I => \N__13300\
        );

    \I__1573\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13290\
        );

    \I__1572\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13287\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__13300\,
            I => \N__13284\
        );

    \I__1570\ : InMux
    port map (
            O => \N__13299\,
            I => \N__13277\
        );

    \I__1569\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13277\
        );

    \I__1568\ : InMux
    port map (
            O => \N__13297\,
            I => \N__13277\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__13296\,
            I => \N__13271\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__13295\,
            I => \N__13265\
        );

    \I__1565\ : InMux
    port map (
            O => \N__13294\,
            I => \N__13261\
        );

    \I__1564\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13258\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__13290\,
            I => \N__13251\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__13287\,
            I => \N__13251\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__13284\,
            I => \N__13251\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__13277\,
            I => \N__13248\
        );

    \I__1559\ : InMux
    port map (
            O => \N__13276\,
            I => \N__13245\
        );

    \I__1558\ : InMux
    port map (
            O => \N__13275\,
            I => \N__13236\
        );

    \I__1557\ : InMux
    port map (
            O => \N__13274\,
            I => \N__13236\
        );

    \I__1556\ : InMux
    port map (
            O => \N__13271\,
            I => \N__13236\
        );

    \I__1555\ : InMux
    port map (
            O => \N__13270\,
            I => \N__13236\
        );

    \I__1554\ : InMux
    port map (
            O => \N__13269\,
            I => \N__13227\
        );

    \I__1553\ : InMux
    port map (
            O => \N__13268\,
            I => \N__13227\
        );

    \I__1552\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13227\
        );

    \I__1551\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13227\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__13261\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__13258\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__13251\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__13248\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__13245\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__13236\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__13227\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1543\ : InMux
    port map (
            O => \N__13212\,
            I => \N__13208\
        );

    \I__1542\ : InMux
    port map (
            O => \N__13211\,
            I => \N__13205\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__13208\,
            I => \N__13202\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__13205\,
            I => \this_vga_signals.N_4_0_0_1\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__13202\,
            I => \this_vga_signals.N_4_0_0_1\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__13197\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_cascade_\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__13194\,
            I => \N__13191\
        );

    \I__1536\ : InMux
    port map (
            O => \N__13191\,
            I => \N__13188\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__13188\,
            I => \N__13185\
        );

    \I__1534\ : Span4Mux_h
    port map (
            O => \N__13185\,
            I => \N__13182\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__13182\,
            I => \M_this_vga_signals_address_3\
        );

    \I__1532\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13176\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__13176\,
            I => \this_vga_signals.if_m2_0\
        );

    \I__1530\ : InMux
    port map (
            O => \N__13173\,
            I => \N__13167\
        );

    \I__1529\ : InMux
    port map (
            O => \N__13172\,
            I => \N__13167\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__13167\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1527\ : InMux
    port map (
            O => \N__13164\,
            I => \N__13161\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__13161\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__13158\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\
        );

    \I__1524\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13152\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__13152\,
            I => \this_vga_signals.mult1_un82_sum_c3_0\
        );

    \I__1522\ : InMux
    port map (
            O => \N__13149\,
            I => \N__13144\
        );

    \I__1521\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13139\
        );

    \I__1520\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13139\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__13144\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__13139\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__13134\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\
        );

    \I__1516\ : InMux
    port map (
            O => \N__13131\,
            I => \N__13128\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__13128\,
            I => \N__13125\
        );

    \I__1514\ : Span4Mux_h
    port map (
            O => \N__13125\,
            I => \N__13122\
        );

    \I__1513\ : Span4Mux_h
    port map (
            O => \N__13122\,
            I => \N__13117\
        );

    \I__1512\ : InMux
    port map (
            O => \N__13121\,
            I => \N__13114\
        );

    \I__1511\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13111\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__13117\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__13114\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__13111\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__13104\,
            I => \N__13101\
        );

    \I__1506\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13098\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__13098\,
            I => \N__13095\
        );

    \I__1504\ : Span4Mux_h
    port map (
            O => \N__13095\,
            I => \N__13092\
        );

    \I__1503\ : Odrv4
    port map (
            O => \N__13092\,
            I => \M_this_vga_signals_address_1\
        );

    \I__1502\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13082\
        );

    \I__1501\ : InMux
    port map (
            O => \N__13088\,
            I => \N__13082\
        );

    \I__1500\ : InMux
    port map (
            O => \N__13087\,
            I => \N__13079\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__13082\,
            I => \N__13076\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__13079\,
            I => \this_vga_signals.mult1_un75_sum_axb1\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__13076\,
            I => \this_vga_signals.mult1_un75_sum_axb1\
        );

    \I__1496\ : InMux
    port map (
            O => \N__13071\,
            I => \N__13067\
        );

    \I__1495\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13064\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__13067\,
            I => \this_vga_signals.mult1_un68_sum_ac0_2\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__13064\,
            I => \this_vga_signals.mult1_un68_sum_ac0_2\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__13059\,
            I => \this_vga_signals.g2_0_0_cascade_\
        );

    \I__1491\ : InMux
    port map (
            O => \N__13056\,
            I => \N__13053\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__13053\,
            I => \this_vga_signals.g0_0_0_a3_0\
        );

    \I__1489\ : InMux
    port map (
            O => \N__13050\,
            I => \N__13047\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__13047\,
            I => \N__13044\
        );

    \I__1487\ : Span4Mux_h
    port map (
            O => \N__13044\,
            I => \N__13040\
        );

    \I__1486\ : InMux
    port map (
            O => \N__13043\,
            I => \N__13037\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__13040\,
            I => \this_vga_signals.vaddress_c3_0\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__13037\,
            I => \this_vga_signals.vaddress_c3_0\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__13032\,
            I => \N__13029\
        );

    \I__1482\ : InMux
    port map (
            O => \N__13029\,
            I => \N__13026\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__13026\,
            I => \N__13022\
        );

    \I__1480\ : InMux
    port map (
            O => \N__13025\,
            I => \N__13019\
        );

    \I__1479\ : Span4Mux_h
    port map (
            O => \N__13022\,
            I => \N__13014\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__13019\,
            I => \N__13014\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__13014\,
            I => \this_vga_signals.SUM_2_i_1_1_3\
        );

    \I__1476\ : InMux
    port map (
            O => \N__13011\,
            I => \N__13008\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__13008\,
            I => \N__13005\
        );

    \I__1474\ : Span4Mux_h
    port map (
            O => \N__13005\,
            I => \N__13001\
        );

    \I__1473\ : InMux
    port map (
            O => \N__13004\,
            I => \N__12998\
        );

    \I__1472\ : Odrv4
    port map (
            O => \N__13001\,
            I => \this_vga_signals.SUM_2_i_1_2_3\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__12998\,
            I => \this_vga_signals.SUM_2_i_1_2_3\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__12993\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i_0_cascade_\
        );

    \I__1469\ : InMux
    port map (
            O => \N__12990\,
            I => \N__12987\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__12987\,
            I => \this_vga_signals.g0_i_x4_0\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__12984\,
            I => \this_vga_signals.g0_i_x4_4_1_cascade_\
        );

    \I__1466\ : InMux
    port map (
            O => \N__12981\,
            I => \N__12978\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__12978\,
            I => \N__12975\
        );

    \I__1464\ : Span4Mux_h
    port map (
            O => \N__12975\,
            I => \N__12972\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__12972\,
            I => \this_vga_signals.g0_i_x4_4\
        );

    \I__1462\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12958\
        );

    \I__1461\ : InMux
    port map (
            O => \N__12968\,
            I => \N__12958\
        );

    \I__1460\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12955\
        );

    \I__1459\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12950\
        );

    \I__1458\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12950\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__12964\,
            I => \N__12946\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__12963\,
            I => \N__12940\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__12958\,
            I => \N__12932\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__12955\,
            I => \N__12932\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__12950\,
            I => \N__12929\
        );

    \I__1452\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12926\
        );

    \I__1451\ : InMux
    port map (
            O => \N__12946\,
            I => \N__12921\
        );

    \I__1450\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12921\
        );

    \I__1449\ : InMux
    port map (
            O => \N__12944\,
            I => \N__12918\
        );

    \I__1448\ : InMux
    port map (
            O => \N__12943\,
            I => \N__12911\
        );

    \I__1447\ : InMux
    port map (
            O => \N__12940\,
            I => \N__12911\
        );

    \I__1446\ : InMux
    port map (
            O => \N__12939\,
            I => \N__12911\
        );

    \I__1445\ : InMux
    port map (
            O => \N__12938\,
            I => \N__12908\
        );

    \I__1444\ : InMux
    port map (
            O => \N__12937\,
            I => \N__12905\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__12932\,
            I => \N__12902\
        );

    \I__1442\ : Span4Mux_h
    port map (
            O => \N__12929\,
            I => \N__12891\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__12926\,
            I => \N__12891\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__12921\,
            I => \N__12891\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__12918\,
            I => \N__12891\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__12911\,
            I => \N__12891\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__12908\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__12905\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__12902\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__12891\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1433\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12876\
        );

    \I__1432\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12872\
        );

    \I__1431\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12869\
        );

    \I__1430\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12866\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__12876\,
            I => \N__12863\
        );

    \I__1428\ : InMux
    port map (
            O => \N__12875\,
            I => \N__12859\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__12872\,
            I => \N__12856\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__12869\,
            I => \N__12846\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__12866\,
            I => \N__12841\
        );

    \I__1424\ : Span4Mux_h
    port map (
            O => \N__12863\,
            I => \N__12841\
        );

    \I__1423\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12838\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__12859\,
            I => \N__12833\
        );

    \I__1421\ : Span4Mux_h
    port map (
            O => \N__12856\,
            I => \N__12833\
        );

    \I__1420\ : InMux
    port map (
            O => \N__12855\,
            I => \N__12826\
        );

    \I__1419\ : InMux
    port map (
            O => \N__12854\,
            I => \N__12826\
        );

    \I__1418\ : InMux
    port map (
            O => \N__12853\,
            I => \N__12826\
        );

    \I__1417\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12823\
        );

    \I__1416\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12816\
        );

    \I__1415\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12816\
        );

    \I__1414\ : InMux
    port map (
            O => \N__12849\,
            I => \N__12816\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__12846\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__12841\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__12838\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__12833\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__12826\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__12823\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__12816\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1406\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12798\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__12798\,
            I => \this_vga_signals.g2_0\
        );

    \I__1404\ : InMux
    port map (
            O => \N__12795\,
            I => \N__12792\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__12792\,
            I => \N__12789\
        );

    \I__1402\ : Span4Mux_v
    port map (
            O => \N__12789\,
            I => \N__12786\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__12786\,
            I => \this_vga_signals.g0_2_0_a2\
        );

    \I__1400\ : InMux
    port map (
            O => \N__12783\,
            I => \N__12777\
        );

    \I__1399\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12777\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__12777\,
            I => \N__12773\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__12776\,
            I => \N__12769\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__12773\,
            I => \N__12764\
        );

    \I__1395\ : InMux
    port map (
            O => \N__12772\,
            I => \N__12759\
        );

    \I__1394\ : InMux
    port map (
            O => \N__12769\,
            I => \N__12759\
        );

    \I__1393\ : InMux
    port map (
            O => \N__12768\,
            I => \N__12754\
        );

    \I__1392\ : InMux
    port map (
            O => \N__12767\,
            I => \N__12754\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__12764\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_ns\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__12759\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_ns\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__12754\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_ns\
        );

    \I__1388\ : InMux
    port map (
            O => \N__12747\,
            I => \N__12744\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__12744\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__12741\,
            I => \this_vga_signals.g0_13_x0_cascade_\
        );

    \I__1385\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12735\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__12735\,
            I => \this_vga_signals.mult1_un68_sum_axb1_1\
        );

    \I__1383\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12729\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__12729\,
            I => \this_vga_signals.mult1_un47_sum_c3_1\
        );

    \I__1381\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12721\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__12725\,
            I => \N__12718\
        );

    \I__1379\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12714\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__12721\,
            I => \N__12708\
        );

    \I__1377\ : InMux
    port map (
            O => \N__12718\,
            I => \N__12703\
        );

    \I__1376\ : InMux
    port map (
            O => \N__12717\,
            I => \N__12703\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__12714\,
            I => \N__12700\
        );

    \I__1374\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12697\
        );

    \I__1373\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12694\
        );

    \I__1372\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12691\
        );

    \I__1371\ : Odrv4
    port map (
            O => \N__12708\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__12703\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__12700\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__12697\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__12694\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__12691\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1365\ : InMux
    port map (
            O => \N__12678\,
            I => \N__12675\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__12675\,
            I => \N__12671\
        );

    \I__1363\ : InMux
    port map (
            O => \N__12674\,
            I => \N__12668\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__12671\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_2\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__12668\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_2\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__12663\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_2_cascade_\
        );

    \I__1359\ : InMux
    port map (
            O => \N__12660\,
            I => \N__12657\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__12657\,
            I => \this_vga_signals.g0_13_x1\
        );

    \I__1357\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12648\
        );

    \I__1356\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12642\
        );

    \I__1355\ : InMux
    port map (
            O => \N__12652\,
            I => \N__12637\
        );

    \I__1354\ : InMux
    port map (
            O => \N__12651\,
            I => \N__12637\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__12648\,
            I => \N__12634\
        );

    \I__1352\ : InMux
    port map (
            O => \N__12647\,
            I => \N__12631\
        );

    \I__1351\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12626\
        );

    \I__1350\ : InMux
    port map (
            O => \N__12645\,
            I => \N__12626\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__12642\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__12637\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__12634\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__12631\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__12626\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1344\ : InMux
    port map (
            O => \N__12615\,
            I => \N__12612\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__12612\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_x0\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__12609\,
            I => \this_vga_signals.mult1_un61_sum_c3_cascade_\
        );

    \I__1341\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12598\
        );

    \I__1340\ : InMux
    port map (
            O => \N__12605\,
            I => \N__12598\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__12604\,
            I => \N__12594\
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__12603\,
            I => \N__12590\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__12598\,
            I => \N__12586\
        );

    \I__1336\ : InMux
    port map (
            O => \N__12597\,
            I => \N__12583\
        );

    \I__1335\ : InMux
    port map (
            O => \N__12594\,
            I => \N__12572\
        );

    \I__1334\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12572\
        );

    \I__1333\ : InMux
    port map (
            O => \N__12590\,
            I => \N__12572\
        );

    \I__1332\ : InMux
    port map (
            O => \N__12589\,
            I => \N__12572\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__12586\,
            I => \N__12569\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__12583\,
            I => \N__12566\
        );

    \I__1329\ : InMux
    port map (
            O => \N__12582\,
            I => \N__12563\
        );

    \I__1328\ : InMux
    port map (
            O => \N__12581\,
            I => \N__12560\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__12572\,
            I => \N__12557\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__12569\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__12566\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__12563\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__12560\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__12557\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__1321\ : InMux
    port map (
            O => \N__12546\,
            I => \N__12543\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__12543\,
            I => \N__12534\
        );

    \I__1319\ : InMux
    port map (
            O => \N__12542\,
            I => \N__12529\
        );

    \I__1318\ : InMux
    port map (
            O => \N__12541\,
            I => \N__12529\
        );

    \I__1317\ : InMux
    port map (
            O => \N__12540\,
            I => \N__12524\
        );

    \I__1316\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12524\
        );

    \I__1315\ : InMux
    port map (
            O => \N__12538\,
            I => \N__12519\
        );

    \I__1314\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12519\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__12534\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__12529\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__12524\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__12519\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__12510\,
            I => \N__12507\
        );

    \I__1308\ : InMux
    port map (
            O => \N__12507\,
            I => \N__12504\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__12504\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_x1\
        );

    \I__1306\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12498\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__12498\,
            I => \this_vga_signals.g1_2_1_0\
        );

    \I__1304\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12492\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__12492\,
            I => \N__12489\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__12489\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_0\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__12486\,
            I => \this_vga_signals.M_vcounter_q_RNITVMCUZ0Z_3_cascade_\
        );

    \I__1300\ : InMux
    port map (
            O => \N__12483\,
            I => \N__12480\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__12480\,
            I => \this_vga_signals.M_vcounter_q_RNIANU4QZ0Z_3\
        );

    \I__1298\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12474\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__12474\,
            I => \N__12471\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__12471\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__12468\,
            I => \this_vga_signals.g1_0_1_cascade_\
        );

    \I__1294\ : InMux
    port map (
            O => \N__12465\,
            I => \N__12462\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__12462\,
            I => \this_vga_signals.g0_i_x4_0_0\
        );

    \I__1292\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12456\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__12456\,
            I => \N__12453\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__12453\,
            I => \this_vga_signals.g1\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__12450\,
            I => \N__12447\
        );

    \I__1288\ : InMux
    port map (
            O => \N__12447\,
            I => \N__12444\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__12444\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1\
        );

    \I__1286\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12438\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__12438\,
            I => \N__12435\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__12435\,
            I => \N__12432\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__12432\,
            I => \this_vga_signals.g0_1_0_0\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__12429\,
            I => \this_vga_signals.g1_2_1_cascade_\
        );

    \I__1281\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12423\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__12423\,
            I => \this_vga_signals.g0_0_0_0_0\
        );

    \I__1279\ : InMux
    port map (
            O => \N__12420\,
            I => \N__12417\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__12417\,
            I => \this_vga_signals.g0_2_0_a2_1\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__12414\,
            I => \this_vga_signals.g0_2_0_a2_1_cascade_\
        );

    \I__1276\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12408\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__12408\,
            I => \this_vga_signals.g0_3_x1\
        );

    \I__1274\ : InMux
    port map (
            O => \N__12405\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__1273\ : InMux
    port map (
            O => \N__12402\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__1272\ : InMux
    port map (
            O => \N__12399\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__1271\ : InMux
    port map (
            O => \N__12396\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__1270\ : InMux
    port map (
            O => \N__12393\,
            I => \bfn_11_24_0_\
        );

    \I__1269\ : CEMux
    port map (
            O => \N__12390\,
            I => \N__12387\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__12387\,
            I => \N__12384\
        );

    \I__1267\ : Span4Mux_h
    port map (
            O => \N__12384\,
            I => \N__12381\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__12381\,
            I => \this_vga_signals.N_692_1\
        );

    \I__1265\ : SRMux
    port map (
            O => \N__12378\,
            I => \N__12375\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__12375\,
            I => \N__12370\
        );

    \I__1263\ : SRMux
    port map (
            O => \N__12374\,
            I => \N__12367\
        );

    \I__1262\ : SRMux
    port map (
            O => \N__12373\,
            I => \N__12364\
        );

    \I__1261\ : Span4Mux_v
    port map (
            O => \N__12370\,
            I => \N__12358\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__12367\,
            I => \N__12358\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__12364\,
            I => \N__12355\
        );

    \I__1258\ : InMux
    port map (
            O => \N__12363\,
            I => \N__12352\
        );

    \I__1257\ : Span4Mux_h
    port map (
            O => \N__12358\,
            I => \N__12349\
        );

    \I__1256\ : Span4Mux_h
    port map (
            O => \N__12355\,
            I => \N__12344\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__12352\,
            I => \N__12344\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__12349\,
            I => \this_vga_signals.M_vcounter_q_379_0\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__12344\,
            I => \this_vga_signals.M_vcounter_q_379_0\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__12339\,
            I => \this_vga_signals.g0_3_x0_cascade_\
        );

    \I__1251\ : InMux
    port map (
            O => \N__12336\,
            I => \N__12333\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__12333\,
            I => \N__12330\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__12330\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0\
        );

    \I__1248\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12324\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__12324\,
            I => \this_vga_signals.M_hcounter_d7lto7_1\
        );

    \I__1246\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12318\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__12318\,
            I => \this_vga_signals.un2_hsynclto3_0\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__12315\,
            I => \this_vga_signals.un2_hsynclto3_0_cascade_\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__12312\,
            I => \this_vga_signals.un2_hsynclto6_0_cascade_\
        );

    \I__1242\ : IoInMux
    port map (
            O => \N__12309\,
            I => \N__12306\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__12306\,
            I => \N__12303\
        );

    \I__1240\ : Span4Mux_s3_h
    port map (
            O => \N__12303\,
            I => \N__12300\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__12300\,
            I => \N__12297\
        );

    \I__1238\ : Span4Mux_v
    port map (
            O => \N__12297\,
            I => \N__12294\
        );

    \I__1237\ : Span4Mux_v
    port map (
            O => \N__12294\,
            I => \N__12291\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__12291\,
            I => rgb_c_4
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__12288\,
            I => \N__12284\
        );

    \I__1234\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12277\
        );

    \I__1233\ : InMux
    port map (
            O => \N__12284\,
            I => \N__12272\
        );

    \I__1232\ : InMux
    port map (
            O => \N__12283\,
            I => \N__12272\
        );

    \I__1231\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12269\
        );

    \I__1230\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12264\
        );

    \I__1229\ : InMux
    port map (
            O => \N__12280\,
            I => \N__12264\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__12277\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__12272\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__12269\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__12264\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1224\ : InMux
    port map (
            O => \N__12255\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__1223\ : InMux
    port map (
            O => \N__12252\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__1222\ : InMux
    port map (
            O => \N__12249\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__12246\,
            I => \this_vga_signals.g3_0_0_0_cascade_\
        );

    \I__1220\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12240\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__12240\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0_0\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__12237\,
            I => \this_vga_signals.M_hcounter_d7lt7_0_cascade_\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__12234\,
            I => \this_vga_signals.if_m2_0_cascade_\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__12231\,
            I => \this_vga_signals.mult1_un89_sum_c3_0_1_cascade_\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__12228\,
            I => \this_vga_signals.haddress_1_0_cascade_\
        );

    \I__1214\ : CascadeMux
    port map (
            O => \N__12225\,
            I => \N__12222\
        );

    \I__1213\ : InMux
    port map (
            O => \N__12222\,
            I => \N__12219\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__12219\,
            I => \N__12216\
        );

    \I__1211\ : Span4Mux_h
    port map (
            O => \N__12216\,
            I => \N__12213\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__12213\,
            I => \N__12210\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__12210\,
            I => \M_this_vga_signals_address_0\
        );

    \I__1208\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12200\
        );

    \I__1207\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12197\
        );

    \I__1206\ : InMux
    port map (
            O => \N__12205\,
            I => \N__12192\
        );

    \I__1205\ : InMux
    port map (
            O => \N__12204\,
            I => \N__12192\
        );

    \I__1204\ : InMux
    port map (
            O => \N__12203\,
            I => \N__12189\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__12200\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__12197\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__12192\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__12189\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1199\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12169\
        );

    \I__1198\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12169\
        );

    \I__1197\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12169\
        );

    \I__1196\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12160\
        );

    \I__1195\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12160\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__12169\,
            I => \N__12157\
        );

    \I__1193\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12147\
        );

    \I__1192\ : InMux
    port map (
            O => \N__12167\,
            I => \N__12147\
        );

    \I__1191\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12147\
        );

    \I__1190\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12147\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__12160\,
            I => \N__12142\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__12157\,
            I => \N__12142\
        );

    \I__1187\ : InMux
    port map (
            O => \N__12156\,
            I => \N__12139\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__12147\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__12142\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__12139\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__12132\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_cascade_\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__12129\,
            I => \N__12126\
        );

    \I__1181\ : InMux
    port map (
            O => \N__12126\,
            I => \N__12123\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__12123\,
            I => \N__12120\
        );

    \I__1179\ : Span4Mux_h
    port map (
            O => \N__12120\,
            I => \N__12117\
        );

    \I__1178\ : Odrv4
    port map (
            O => \N__12117\,
            I => \this_vga_signals.if_m8_0_a3_1_1_6\
        );

    \I__1177\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12111\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__12111\,
            I => \N__12108\
        );

    \I__1175\ : Odrv4
    port map (
            O => \N__12108\,
            I => \this_vga_signals.N_5_i_0\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__12105\,
            I => \this_vga_signals.g1_2_1_0_0_cascade_\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__12102\,
            I => \this_vga_signals.g1_0_4_1_cascade_\
        );

    \I__1172\ : InMux
    port map (
            O => \N__12099\,
            I => \N__12096\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__12096\,
            I => \this_vga_signals.mult1_un47_sum_c3_2_0\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__12093\,
            I => \N__12090\
        );

    \I__1169\ : InMux
    port map (
            O => \N__12090\,
            I => \N__12087\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__12087\,
            I => \N__12084\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__12084\,
            I => \this_vga_signals.g1_0_4\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__12081\,
            I => \N__12078\
        );

    \I__1165\ : InMux
    port map (
            O => \N__12078\,
            I => \N__12075\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__12075\,
            I => \N__12072\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__12072\,
            I => \N__12069\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__12069\,
            I => \this_vga_signals.if_m8_0_a3_1_1_4\
        );

    \I__1161\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12063\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__12063\,
            I => \this_vga_signals.g1_0\
        );

    \I__1159\ : InMux
    port map (
            O => \N__12060\,
            I => \N__12057\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__12057\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__12054\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0_cascade_\
        );

    \I__1156\ : InMux
    port map (
            O => \N__12051\,
            I => \N__12048\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__12048\,
            I => \this_vga_signals.g0_1_0_0_0\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__12045\,
            I => \this_vga_signals.g2_1_0_1_cascade_\
        );

    \I__1153\ : InMux
    port map (
            O => \N__12042\,
            I => \N__12034\
        );

    \I__1152\ : InMux
    port map (
            O => \N__12041\,
            I => \N__12034\
        );

    \I__1151\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12029\
        );

    \I__1150\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12029\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__12034\,
            I => \N__12024\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__12029\,
            I => \N__12024\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__12024\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__12021\,
            I => \N__12016\
        );

    \I__1145\ : InMux
    port map (
            O => \N__12020\,
            I => \N__12012\
        );

    \I__1144\ : InMux
    port map (
            O => \N__12019\,
            I => \N__12009\
        );

    \I__1143\ : InMux
    port map (
            O => \N__12016\,
            I => \N__12004\
        );

    \I__1142\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12004\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__12012\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__12009\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__12004\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__11997\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\
        );

    \I__1137\ : InMux
    port map (
            O => \N__11994\,
            I => \N__11987\
        );

    \I__1136\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11987\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__11992\,
            I => \N__11984\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__11987\,
            I => \N__11979\
        );

    \I__1133\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11976\
        );

    \I__1132\ : InMux
    port map (
            O => \N__11983\,
            I => \N__11971\
        );

    \I__1131\ : InMux
    port map (
            O => \N__11982\,
            I => \N__11971\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__11979\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__11976\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__11971\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__1127\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11961\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__11961\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_0\
        );

    \I__1125\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11947\
        );

    \I__1124\ : InMux
    port map (
            O => \N__11957\,
            I => \N__11947\
        );

    \I__1123\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11944\
        );

    \I__1122\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11939\
        );

    \I__1121\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11939\
        );

    \I__1120\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11934\
        );

    \I__1119\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11934\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__11947\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__11944\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__11939\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__11934\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__11925\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\
        );

    \I__1113\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11919\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__11919\,
            I => \N__11914\
        );

    \I__1111\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11911\
        );

    \I__1110\ : InMux
    port map (
            O => \N__11917\,
            I => \N__11908\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__11914\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__11911\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__11908\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__11901\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\
        );

    \I__1105\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11895\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__11895\,
            I => \N__11892\
        );

    \I__1103\ : Span4Mux_h
    port map (
            O => \N__11892\,
            I => \N__11889\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__11889\,
            I => \this_vga_signals.g1_0_0_0\
        );

    \I__1101\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11883\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__11883\,
            I => \N__11880\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__11880\,
            I => \this_vga_signals.vaddress_2_5\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__11877\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_x0_cascade_\
        );

    \I__1097\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11867\
        );

    \I__1096\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11859\
        );

    \I__1095\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11859\
        );

    \I__1094\ : InMux
    port map (
            O => \N__11871\,
            I => \N__11859\
        );

    \I__1093\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11856\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__11867\,
            I => \N__11853\
        );

    \I__1091\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11850\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__11859\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__11856\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__11853\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__11850\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1086\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11837\
        );

    \I__1085\ : InMux
    port map (
            O => \N__11840\,
            I => \N__11834\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__11837\,
            I => \N__11831\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__11834\,
            I => \N__11828\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__11831\,
            I => \this_vga_signals.if_m8_0_a3_1_1_1\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__11828\,
            I => \this_vga_signals.if_m8_0_a3_1_1_1\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__11823\,
            I => \this_vga_signals.if_N_5_cascade_\
        );

    \I__1079\ : InMux
    port map (
            O => \N__11820\,
            I => \N__11817\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__11817\,
            I => \N__11814\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__11814\,
            I => \this_vga_signals.if_m8_0_a3_1_1_0\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__11811\,
            I => \this_vga_signals.N_5_i_0_cascade_\
        );

    \I__1075\ : InMux
    port map (
            O => \N__11808\,
            I => \N__11805\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__11805\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__1073\ : InMux
    port map (
            O => \N__11802\,
            I => \N__11797\
        );

    \I__1072\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11792\
        );

    \I__1071\ : InMux
    port map (
            O => \N__11800\,
            I => \N__11792\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__11797\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__11792\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1068\ : InMux
    port map (
            O => \N__11787\,
            I => \N__11782\
        );

    \I__1067\ : InMux
    port map (
            O => \N__11786\,
            I => \N__11777\
        );

    \I__1066\ : InMux
    port map (
            O => \N__11785\,
            I => \N__11777\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__11782\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__11777\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1063\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11769\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__11769\,
            I => \N__11766\
        );

    \I__1061\ : Span4Mux_h
    port map (
            O => \N__11766\,
            I => \N__11763\
        );

    \I__1060\ : Odrv4
    port map (
            O => \N__11763\,
            I => \this_vga_signals.SUM_3_1_tz\
        );

    \I__1059\ : IoInMux
    port map (
            O => \N__11760\,
            I => \N__11757\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__1057\ : IoSpan4Mux
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__1056\ : IoSpan4Mux
    port map (
            O => \N__11751\,
            I => \N__11748\
        );

    \I__1055\ : Span4Mux_s1_v
    port map (
            O => \N__11748\,
            I => \N__11745\
        );

    \I__1054\ : Span4Mux_v
    port map (
            O => \N__11745\,
            I => \N__11742\
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__11742\,
            I => this_vga_signals_hvisibility_i
        );

    \I__1052\ : SRMux
    port map (
            O => \N__11739\,
            I => \N__11736\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__11736\,
            I => \N__11732\
        );

    \I__1050\ : SRMux
    port map (
            O => \N__11735\,
            I => \N__11729\
        );

    \I__1049\ : Span4Mux_h
    port map (
            O => \N__11732\,
            I => \N__11726\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__11729\,
            I => \N__11723\
        );

    \I__1047\ : Odrv4
    port map (
            O => \N__11726\,
            I => \M_stage_q_RNIC68K4_9\
        );

    \I__1046\ : Odrv12
    port map (
            O => \N__11723\,
            I => \M_stage_q_RNIC68K4_9\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__11718\,
            I => \N__11715\
        );

    \I__1044\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11712\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__11712\,
            I => \N__11708\
        );

    \I__1042\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11705\
        );

    \I__1041\ : Span4Mux_h
    port map (
            O => \N__11708\,
            I => \N__11702\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__11705\,
            I => \this_vga_signals.vaddress_3_5\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__11702\,
            I => \this_vga_signals.vaddress_3_5\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__11697\,
            I => \this_vga_signals.if_m8_0_a3_1_1_5_cascade_\
        );

    \I__1037\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11691\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__11691\,
            I => \N__11688\
        );

    \I__1035\ : Span4Mux_v
    port map (
            O => \N__11688\,
            I => \N__11685\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__11685\,
            I => \this_vga_signals.g0_6_0_0\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__11682\,
            I => \this_vga_signals.un6_vvisibilitylt8_cascade_\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__11679\,
            I => \N__11676\
        );

    \I__1031\ : InMux
    port map (
            O => \N__11676\,
            I => \N__11673\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__11673\,
            I => \this_vga_signals.vvisibility_1\
        );

    \I__1029\ : InMux
    port map (
            O => \N__11670\,
            I => \N__11667\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__11667\,
            I => \this_vga_signals.vaddress_0_5\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__11664\,
            I => \this_vga_signals.if_m8_0_a3_1_1_3_cascade_\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__11661\,
            I => \this_vga_signals.g0_6_0_cascade_\
        );

    \I__1025\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11655\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__11655\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d\
        );

    \I__1023\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11649\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__11649\,
            I => \N__11646\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__11646\,
            I => \this_vga_signals.i6_mux_0\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__11643\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_\
        );

    \I__1019\ : InMux
    port map (
            O => \N__11640\,
            I => \N__11637\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__11637\,
            I => \this_vga_signals.g0_i_x4_0_a2_1\
        );

    \I__1017\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11631\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__11631\,
            I => \N__11628\
        );

    \I__1015\ : Span4Mux_v
    port map (
            O => \N__11628\,
            I => \N__11625\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__11625\,
            I => \this_vga_signals.if_m8_0_a3_1_1_2\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__11622\,
            I => \this_vga_signals.vaddress_1_0_5_cascade_\
        );

    \I__1012\ : CascadeMux
    port map (
            O => \N__11619\,
            I => \this_vga_signals.SUM_2_i_1_1_3_cascade_\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__11616\,
            I => \N__11613\
        );

    \I__1010\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11610\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__11610\,
            I => \this_vga_signals.SUM_2_i_1_1_1_3\
        );

    \I__1008\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11604\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__11604\,
            I => \N__11601\
        );

    \I__1006\ : Odrv4
    port map (
            O => \N__11601\,
            I => \this_vga_signals.N_1_3_1\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__11598\,
            I => \this_vga_signals.N_1_3_1_cascade_\
        );

    \I__1004\ : InMux
    port map (
            O => \N__11595\,
            I => \N__11592\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__11592\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__11589\,
            I => \N__11586\
        );

    \I__1001\ : CascadeBuf
    port map (
            O => \N__11586\,
            I => \N__11583\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__11583\,
            I => \N__11580\
        );

    \I__999\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11577\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__11577\,
            I => \N__11573\
        );

    \I__997\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11570\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__11573\,
            I => \N__11567\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__11570\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__11567\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__993\ : InMux
    port map (
            O => \N__11562\,
            I => \un1_M_this_map_address_q_cry_5\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__11559\,
            I => \N__11556\
        );

    \I__991\ : CascadeBuf
    port map (
            O => \N__11556\,
            I => \N__11553\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__11553\,
            I => \N__11550\
        );

    \I__989\ : InMux
    port map (
            O => \N__11550\,
            I => \N__11547\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__11547\,
            I => \N__11543\
        );

    \I__987\ : InMux
    port map (
            O => \N__11546\,
            I => \N__11540\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__11543\,
            I => \N__11537\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__11540\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__11537\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__983\ : InMux
    port map (
            O => \N__11532\,
            I => \un1_M_this_map_address_q_cry_6\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__11529\,
            I => \N__11526\
        );

    \I__981\ : CascadeBuf
    port map (
            O => \N__11526\,
            I => \N__11523\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__11523\,
            I => \N__11520\
        );

    \I__979\ : InMux
    port map (
            O => \N__11520\,
            I => \N__11517\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__11517\,
            I => \N__11513\
        );

    \I__977\ : InMux
    port map (
            O => \N__11516\,
            I => \N__11510\
        );

    \I__976\ : Span4Mux_v
    port map (
            O => \N__11513\,
            I => \N__11507\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__11510\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__974\ : Odrv4
    port map (
            O => \N__11507\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__973\ : InMux
    port map (
            O => \N__11502\,
            I => \bfn_9_24_0_\
        );

    \I__972\ : InMux
    port map (
            O => \N__11499\,
            I => \un1_M_this_map_address_q_cry_8\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__11496\,
            I => \N__11493\
        );

    \I__970\ : CascadeBuf
    port map (
            O => \N__11493\,
            I => \N__11490\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__11490\,
            I => \N__11487\
        );

    \I__968\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11484\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__11484\,
            I => \N__11480\
        );

    \I__966\ : InMux
    port map (
            O => \N__11483\,
            I => \N__11477\
        );

    \I__965\ : Span4Mux_v
    port map (
            O => \N__11480\,
            I => \N__11474\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__11477\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__963\ : Odrv4
    port map (
            O => \N__11474\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__962\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11466\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__11466\,
            I => \N_89_0\
        );

    \I__960\ : InMux
    port map (
            O => \N__11463\,
            I => \N__11460\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__11460\,
            I => \N_83_0\
        );

    \I__958\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11454\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__11454\,
            I => \N__11451\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__11451\,
            I => \N_85_0\
        );

    \I__955\ : CascadeMux
    port map (
            O => \N__11448\,
            I => \this_vga_signals.vaddress_3_0_5_cascade_\
        );

    \I__954\ : InMux
    port map (
            O => \N__11445\,
            I => \N__11442\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__11442\,
            I => \N__11439\
        );

    \I__952\ : Span4Mux_h
    port map (
            O => \N__11439\,
            I => \N__11436\
        );

    \I__951\ : Odrv4
    port map (
            O => \N__11436\,
            I => \this_vga_signals.g0_6_0_0_0\
        );

    \I__950\ : InMux
    port map (
            O => \N__11433\,
            I => \N__11430\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__11430\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__948\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11424\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__11424\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__946\ : InMux
    port map (
            O => \N__11421\,
            I => \N__11418\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__11418\,
            I => \this_vga_signals.g0_0_0\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__11415\,
            I => \N__11412\
        );

    \I__943\ : CascadeBuf
    port map (
            O => \N__11412\,
            I => \N__11409\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__11409\,
            I => \N__11406\
        );

    \I__941\ : InMux
    port map (
            O => \N__11406\,
            I => \N__11403\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__11403\,
            I => \N__11399\
        );

    \I__939\ : InMux
    port map (
            O => \N__11402\,
            I => \N__11396\
        );

    \I__938\ : Sp12to4
    port map (
            O => \N__11399\,
            I => \N__11393\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__11396\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__936\ : Odrv12
    port map (
            O => \N__11393\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__11388\,
            I => \N__11385\
        );

    \I__934\ : CascadeBuf
    port map (
            O => \N__11385\,
            I => \N__11382\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__11382\,
            I => \N__11379\
        );

    \I__932\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11376\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__11376\,
            I => \N__11372\
        );

    \I__930\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11369\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__11372\,
            I => \N__11366\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__11369\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__11366\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__926\ : InMux
    port map (
            O => \N__11361\,
            I => \un1_M_this_map_address_q_cry_0\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__11358\,
            I => \N__11355\
        );

    \I__924\ : CascadeBuf
    port map (
            O => \N__11355\,
            I => \N__11352\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__11352\,
            I => \N__11349\
        );

    \I__922\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11346\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__11346\,
            I => \N__11342\
        );

    \I__920\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11339\
        );

    \I__919\ : Span4Mux_v
    port map (
            O => \N__11342\,
            I => \N__11336\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__11339\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__917\ : Odrv4
    port map (
            O => \N__11336\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__916\ : InMux
    port map (
            O => \N__11331\,
            I => \un1_M_this_map_address_q_cry_1\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__11328\,
            I => \N__11325\
        );

    \I__914\ : CascadeBuf
    port map (
            O => \N__11325\,
            I => \N__11322\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__11322\,
            I => \N__11319\
        );

    \I__912\ : InMux
    port map (
            O => \N__11319\,
            I => \N__11316\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__11316\,
            I => \N__11312\
        );

    \I__910\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11309\
        );

    \I__909\ : Span4Mux_v
    port map (
            O => \N__11312\,
            I => \N__11306\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__11309\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__11306\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__906\ : InMux
    port map (
            O => \N__11301\,
            I => \un1_M_this_map_address_q_cry_2\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__11298\,
            I => \N__11295\
        );

    \I__904\ : CascadeBuf
    port map (
            O => \N__11295\,
            I => \N__11292\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__11292\,
            I => \N__11289\
        );

    \I__902\ : InMux
    port map (
            O => \N__11289\,
            I => \N__11286\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__11286\,
            I => \N__11282\
        );

    \I__900\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11279\
        );

    \I__899\ : Span4Mux_v
    port map (
            O => \N__11282\,
            I => \N__11276\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__11279\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__11276\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__896\ : InMux
    port map (
            O => \N__11271\,
            I => \un1_M_this_map_address_q_cry_3\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__11268\,
            I => \N__11265\
        );

    \I__894\ : CascadeBuf
    port map (
            O => \N__11265\,
            I => \N__11262\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__11262\,
            I => \N__11259\
        );

    \I__892\ : InMux
    port map (
            O => \N__11259\,
            I => \N__11256\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__11256\,
            I => \N__11252\
        );

    \I__890\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11249\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__11252\,
            I => \N__11246\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__11249\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__887\ : Odrv4
    port map (
            O => \N__11246\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__886\ : InMux
    port map (
            O => \N__11241\,
            I => \un1_M_this_map_address_q_cry_4\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__11238\,
            I => \this_vga_signals.vsync_1_3_cascade_\
        );

    \I__884\ : IoInMux
    port map (
            O => \N__11235\,
            I => \N__11232\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__11232\,
            I => \N__11229\
        );

    \I__882\ : IoSpan4Mux
    port map (
            O => \N__11229\,
            I => \N__11226\
        );

    \I__881\ : Sp12to4
    port map (
            O => \N__11226\,
            I => \N__11223\
        );

    \I__880\ : Span12Mux_v
    port map (
            O => \N__11223\,
            I => \N__11220\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__11220\,
            I => this_vga_signals_vsync_1_i
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__11217\,
            I => \this_vga_signals.g0_2_0_cascade_\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__11214\,
            I => \this_vga_signals.N_43_1_cascade_\
        );

    \I__876\ : InMux
    port map (
            O => \N__11211\,
            I => \N__11208\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__11208\,
            I => \this_vga_signals.un2_vsynclt8\
        );

    \I__874\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11202\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__11202\,
            I => \this_vga_signals.vsync_1_2\
        );

    \I__872\ : InMux
    port map (
            O => \N__11199\,
            I => \N__11196\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__11196\,
            I => \this_vga_signals.g1_1\
        );

    \I__870\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11190\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__11190\,
            I => \N__11187\
        );

    \I__868\ : Span12Mux_h
    port map (
            O => \N__11187\,
            I => \N__11184\
        );

    \I__867\ : Odrv12
    port map (
            O => \N__11184\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__11181\,
            I => \this_vga_signals.g0_0_0_0_cascade_\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__11178\,
            I => \this_vga_signals.g1_1_1_cascade_\
        );

    \I__864\ : InMux
    port map (
            O => \N__11175\,
            I => \N__11172\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__11172\,
            I => \N__11169\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__11169\,
            I => \this_vga_signals.g1_1_0\
        );

    \I__861\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11163\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__11163\,
            I => \this_vga_signals.N_4_0_0\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__11160\,
            I => \this_vga_signals.mult1_un47_sum_c3_0_cascade_\
        );

    \I__858\ : InMux
    port map (
            O => \N__11157\,
            I => \N__11154\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__11154\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_1\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__11151\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_1_cascade_\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__11148\,
            I => \this_vga_signals.g2_1_cascade_\
        );

    \I__854\ : InMux
    port map (
            O => \N__11145\,
            I => \N__11142\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__11142\,
            I => \this_vga_signals.g2\
        );

    \I__852\ : IoInMux
    port map (
            O => \N__11139\,
            I => \N__11136\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__11136\,
            I => \N__11133\
        );

    \I__850\ : Span12Mux_s8_h
    port map (
            O => \N__11133\,
            I => \N__11130\
        );

    \I__849\ : Span12Mux_v
    port map (
            O => \N__11130\,
            I => \N__11127\
        );

    \I__848\ : Odrv12
    port map (
            O => \N__11127\,
            I => rgb_c_0
        );

    \I__847\ : IoInMux
    port map (
            O => \N__11124\,
            I => \N__11121\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__11121\,
            I => \N__11118\
        );

    \I__845\ : Odrv12
    port map (
            O => \N__11118\,
            I => rgb_c_1
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__11115\,
            I => \N__11112\
        );

    \I__843\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11109\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__11109\,
            I => \M_this_vga_signals_address_2\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__11106\,
            I => \N__11103\
        );

    \I__840\ : InMux
    port map (
            O => \N__11103\,
            I => \N__11100\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__11100\,
            I => \N__11097\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__11097\,
            I => \M_this_vga_signals_address_6\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__11094\,
            I => \N__11091\
        );

    \I__836\ : InMux
    port map (
            O => \N__11091\,
            I => \N__11088\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__11088\,
            I => \M_this_vga_signals_address_4\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__11085\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__11082\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_0_cascade_\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__11079\,
            I => \N__11076\
        );

    \I__831\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11073\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__11073\,
            I => \M_this_vga_signals_address_7\
        );

    \I__829\ : IoInMux
    port map (
            O => \N__11070\,
            I => \N__11067\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__11067\,
            I => \this_vga_signals.N_692_0\
        );

    \I__827\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11061\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__11061\,
            I => port_clk_c
        );

    \I__825\ : IoInMux
    port map (
            O => \N__11058\,
            I => \N__11055\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__11055\,
            I => port_data_rw_0_i
        );

    \I__823\ : IoInMux
    port map (
            O => \N__11052\,
            I => \N__11049\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__11049\,
            I => \N__11046\
        );

    \I__821\ : Span4Mux_s2_h
    port map (
            O => \N__11046\,
            I => \N__11043\
        );

    \I__820\ : Span4Mux_v
    port map (
            O => \N__11043\,
            I => \N__11040\
        );

    \I__819\ : Odrv4
    port map (
            O => \N__11040\,
            I => port_nmib_0_i
        );

    \I__818\ : IoInMux
    port map (
            O => \N__11037\,
            I => \N__11034\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__11034\,
            I => \N__11031\
        );

    \I__816\ : Span12Mux_s2_v
    port map (
            O => \N__11031\,
            I => \N__11028\
        );

    \I__815\ : Odrv12
    port map (
            O => \N__11028\,
            I => this_vga_signals_vvisibility_i
        );

    \IN_MUX_bfv_24_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_22_0_\
        );

    \IN_MUX_bfv_24_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_external_address_q_cry_7\,
            carryinitout => \bfn_24_23_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_23_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_19_0_\
        );

    \IN_MUX_bfv_23_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_vaddress_q_cry_7\,
            carryinitout => \bfn_23_20_0_\
        );

    \IN_MUX_bfv_22_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_19_0_\
        );

    \IN_MUX_bfv_22_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_haddress_q_cry_7\,
            carryinitout => \bfn_22_20_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_data_count_q_cry_7\,
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_23_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_16_0_\
        );

    \IN_MUX_bfv_21_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_16_0_\
        );

    \IN_MUX_bfv_22_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_17_0_\
        );

    \IN_MUX_bfv_22_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_vaddress_q_3_cry_7\,
            carryinitout => \bfn_22_18_0_\
        );

    \IN_MUX_bfv_21_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_18_0_\
        );

    \IN_MUX_bfv_21_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_haddress_q_2_cry_7\,
            carryinitout => \bfn_21_19_0_\
        );

    \IN_MUX_bfv_19_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_22_0_\
        );

    \IN_MUX_bfv_19_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_sprites_address_q_cry_7\,
            carryinitout => \bfn_19_23_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_map_address_q_cry_7\,
            carryinitout => \bfn_9_24_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIR1G77_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11070\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_692_0_g\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI67JU6_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__16293\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_988_g\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__22858\,
            GLOBALBUFFEROUTPUT => \M_this_reset_cond_out_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19056\,
            in2 => \_gnd_net_\,
            in3 => \N__14736\,
            lcout => \this_vga_signals.N_692_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11064\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.port_data_rw_0_i_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__21710\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22923\,
            lcout => port_data_rw_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIKCDU5_9_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22931\,
            in2 => \_gnd_net_\,
            in3 => \N__22989\,
            lcout => port_nmib_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_9_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22978\,
            lcout => this_vga_signals_vvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15818\,
            in2 => \_gnd_net_\,
            in3 => \N__14898\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15663\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15819\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIGJMLD1_9_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15590\,
            in2 => \_gnd_net_\,
            in3 => \N__13131\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111101"
        )
    port map (
            in0 => \N__18858\,
            in1 => \N__18813\,
            in2 => \N__18759\,
            in3 => \N__18702\,
            lcout => \this_vga_ramdac.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNILR5N4_8_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__11772\,
            in1 => \N__15587\,
            in2 => \_gnd_net_\,
            in3 => \N__14691\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI9V9QB_9_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15588\,
            in2 => \_gnd_net_\,
            in3 => \N__13476\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12795\,
            in1 => \N__12477\,
            in2 => \N__15403\,
            in3 => \N__12336\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_m2_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011000101"
        )
    port map (
            in0 => \N__15485\,
            in1 => \N__12459\,
            in2 => \N__11085\,
            in3 => \N__12981\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIOIKI4Q_1_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15589\,
            in1 => \N__11175\,
            in2 => \N__11082\,
            in3 => \N__11898\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14205\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34541\,
            ce => \N__14762\,
            sr => \N__14732\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__11445\,
            in1 => \N__11157\,
            in2 => \_gnd_net_\,
            in3 => \N__13387\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_2_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001101"
        )
    port map (
            in0 => \N__11166\,
            in1 => \N__11145\,
            in2 => \N__11181\,
            in3 => \N__13299\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIO70OS4_1_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110111010100"
        )
    port map (
            in0 => \N__15481\,
            in1 => \N__15392\,
            in2 => \N__11178\,
            in3 => \N__11640\,
            lcout => \this_vga_signals.g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13386\,
            in1 => \N__16483\,
            in2 => \N__15306\,
            in3 => \N__13297\,
            lcout => \this_vga_signals.N_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_19_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000111011001"
        )
    port map (
            in0 => \N__12967\,
            in1 => \N__12206\,
            in2 => \N__11718\,
            in3 => \N__12881\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16703\,
            in1 => \N__16482\,
            in2 => \N__11160\,
            in3 => \N__12724\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_3_d_1\,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_3_d_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_1_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011110101"
        )
    port map (
            in0 => \N__11694\,
            in1 => \_gnd_net_\,
            in2 => \N__11151\,
            in3 => \N__13385\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010001001101"
        )
    port map (
            in0 => \N__15391\,
            in1 => \N__15295\,
            in2 => \N__11148\,
            in3 => \N__13298\,
            lcout => \this_vga_signals.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17172\,
            in1 => \N__20108\,
            in2 => \N__16779\,
            in3 => \N__16475\,
            lcout => OPEN,
            ltout => \this_vga_signals.vsync_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__11211\,
            in1 => \N__11205\,
            in2 => \N__11238\,
            in3 => \N__16601\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000010101"
        )
    port map (
            in0 => \N__16600\,
            in1 => \N__16473\,
            in2 => \N__16778\,
            in3 => \N__17066\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110111110000"
        )
    port map (
            in0 => \N__11607\,
            in1 => \N__11421\,
            in2 => \N__11217\,
            in3 => \N__13025\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_43_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__16771\,
            in1 => \N__11199\,
            in2 => \N__11214\,
            in3 => \N__12969\,
            lcout => \this_vga_signals.i6_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010101"
        )
    port map (
            in0 => \N__16474\,
            in1 => \N__15394\,
            in2 => \N__15486\,
            in3 => \N__15296\,
            lcout => \this_vga_signals.un2_vsynclt8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNICSHP_2_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__15395\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17067\,
            lcout => \this_vga_signals.vsync_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110001101"
        )
    port map (
            in0 => \N__12968\,
            in1 => \N__16767\,
            in2 => \N__16490\,
            in3 => \N__12882\,
            lcout => \this_vga_signals.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11427\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11193\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11433\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIP5821_9_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__20103\,
            in1 => \N__17167\,
            in2 => \_gnd_net_\,
            in3 => \N__16609\,
            lcout => \this_vga_signals.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_0_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11402\,
            in2 => \N__18260\,
            in3 => \N__18255\,
            lcout => \M_this_map_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \un1_M_this_map_address_q_cry_0\,
            clk => \N__34575\,
            ce => 'H',
            sr => \N__11739\
        );

    \M_this_map_address_q_1_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11375\,
            in2 => \_gnd_net_\,
            in3 => \N__11361\,
            lcout => \M_this_map_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_0\,
            carryout => \un1_M_this_map_address_q_cry_1\,
            clk => \N__34575\,
            ce => 'H',
            sr => \N__11739\
        );

    \M_this_map_address_q_2_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11345\,
            in2 => \_gnd_net_\,
            in3 => \N__11331\,
            lcout => \M_this_map_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_1\,
            carryout => \un1_M_this_map_address_q_cry_2\,
            clk => \N__34575\,
            ce => 'H',
            sr => \N__11739\
        );

    \M_this_map_address_q_3_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11315\,
            in2 => \_gnd_net_\,
            in3 => \N__11301\,
            lcout => \M_this_map_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_2\,
            carryout => \un1_M_this_map_address_q_cry_3\,
            clk => \N__34575\,
            ce => 'H',
            sr => \N__11739\
        );

    \M_this_map_address_q_4_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11285\,
            in2 => \_gnd_net_\,
            in3 => \N__11271\,
            lcout => \M_this_map_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_3\,
            carryout => \un1_M_this_map_address_q_cry_4\,
            clk => \N__34575\,
            ce => 'H',
            sr => \N__11739\
        );

    \M_this_map_address_q_5_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11255\,
            in2 => \_gnd_net_\,
            in3 => \N__11241\,
            lcout => \M_this_map_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_4\,
            carryout => \un1_M_this_map_address_q_cry_5\,
            clk => \N__34575\,
            ce => 'H',
            sr => \N__11739\
        );

    \M_this_map_address_q_6_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11576\,
            in2 => \_gnd_net_\,
            in3 => \N__11562\,
            lcout => \M_this_map_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_5\,
            carryout => \un1_M_this_map_address_q_cry_6\,
            clk => \N__34575\,
            ce => 'H',
            sr => \N__11739\
        );

    \M_this_map_address_q_7_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11546\,
            in2 => \_gnd_net_\,
            in3 => \N__11532\,
            lcout => \M_this_map_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_6\,
            carryout => \un1_M_this_map_address_q_cry_7\,
            clk => \N__34575\,
            ce => 'H',
            sr => \N__11739\
        );

    \M_this_map_address_q_8_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11516\,
            in2 => \_gnd_net_\,
            in3 => \N__11502\,
            lcout => \M_this_map_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \un1_M_this_map_address_q_cry_8\,
            clk => \N__34580\,
            ce => 'H',
            sr => \N__11735\
        );

    \M_this_map_address_q_9_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11483\,
            in2 => \_gnd_net_\,
            in3 => \N__11499\,
            lcout => \M_this_map_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34580\,
            ce => 'H',
            sr => \N__11735\
        );

    \this_vga_signals.M_this_map_ram_write_data_i_3_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32833\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18256\,
            lcout => \N_89_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_i_6_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18249\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32408\,
            lcout => \N_83_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_i_5_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34766\,
            in2 => \_gnd_net_\,
            in3 => \N__18248\,
            lcout => \N_85_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16753\,
            in2 => \_gnd_net_\,
            in3 => \N__16491\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_3_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_11_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__12875\,
            in1 => \N__11634\,
            in2 => \N__11448\,
            in3 => \N__12938\,
            lcout => \this_vga_signals.g0_6_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14241\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34506\,
            ce => \N__14764\,
            sr => \N__14729\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14838\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34506\,
            ce => \N__14764\,
            sr => \N__14729\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14868\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34506\,
            ce => \N__14764\,
            sr => \N__14729\
        );

    \this_vga_signals.un5_vaddress_g0_5_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100110011111"
        )
    port map (
            in0 => \N__17120\,
            in1 => \N__16534\,
            in2 => \N__20090\,
            in3 => \N__17019\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100110011111"
        )
    port map (
            in0 => \N__17136\,
            in1 => \N__16548\,
            in2 => \N__20078\,
            in3 => \N__17017\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14201\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34514\,
            ce => \N__14761\,
            sr => \N__14726\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100110011111"
        )
    port map (
            in0 => \N__12019\,
            in1 => \N__11954\,
            in2 => \N__11992\,
            in3 => \N__17016\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14837\,
            lcout => \this_vga_signals.M_vcounter_q_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34514\,
            ce => \N__14761\,
            sr => \N__14726\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14233\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34514\,
            ce => \N__14761\,
            sr => \N__14726\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14867\,
            lcout => \this_vga_signals.M_vcounter_q_9_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34514\,
            ce => \N__14761\,
            sr => \N__14726\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_0_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__11866\,
            in1 => \N__12156\,
            in2 => \_gnd_net_\,
            in3 => \N__11955\,
            lcout => \this_vga_signals.vaddress_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34514\,
            ce => \N__14761\,
            sr => \N__14726\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_RNI79KC_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110001"
        )
    port map (
            in0 => \N__11958\,
            in1 => \N__11917\,
            in2 => \N__11616\,
            in3 => \N__11994\,
            lcout => \this_vga_signals.SUM_2_i_1_1_3\,
            ltout => \this_vga_signals.SUM_2_i_1_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__17018\,
            in1 => \N__13043\,
            in2 => \N__11619\,
            in3 => \N__13004\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11785\,
            in2 => \_gnd_net_\,
            in3 => \N__11800\,
            lcout => \this_vga_signals.vaddress_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__11595\,
            in1 => \N__12042\,
            in2 => \_gnd_net_\,
            in3 => \N__14813\,
            lcout => \this_vga_signals.SUM_2_i_1_1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_4_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__12041\,
            in1 => \N__11786\,
            in2 => \_gnd_net_\,
            in3 => \N__11801\,
            lcout => \this_vga_signals.N_1_3_1\,
            ltout => \this_vga_signals.N_1_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_RNICPER_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001111"
        )
    port map (
            in0 => \N__11993\,
            in1 => \N__12020\,
            in2 => \N__11598\,
            in3 => \N__11957\,
            lcout => \this_vga_signals.SUM_2_i_1_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14866\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__14765\,
            sr => \N__14730\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14796\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__14765\,
            sr => \N__14730\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16686\,
            in2 => \_gnd_net_\,
            in3 => \N__16476\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_1_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_25_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011000000110"
        )
    port map (
            in0 => \N__12854\,
            in1 => \N__12945\,
            in2 => \N__11622\,
            in3 => \N__11841\,
            lcout => \this_vga_signals.g0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_24_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001111001011"
        )
    port map (
            in0 => \N__12606\,
            in1 => \N__12207\,
            in2 => \N__12964\,
            in3 => \N__12855\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14264\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34534\,
            ce => \N__14766\,
            sr => \N__14731\
        );

    \this_vga_signals.un5_vaddress_g1_0_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010000111"
        )
    port map (
            in0 => \N__12176\,
            in1 => \N__16685\,
            in2 => \N__16602\,
            in3 => \N__12853\,
            lcout => \this_vga_signals.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14265\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34534\,
            ce => \N__14766\,
            sr => \N__14731\
        );

    \this_vga_signals.un5_vaddress_g0_7_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__16488\,
            in1 => \N__12717\,
            in2 => \N__16736\,
            in3 => \N__12651\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__12652\,
            in1 => \N__12605\,
            in2 => \N__12725\,
            in3 => \N__12177\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_3_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16691\,
            in2 => \_gnd_net_\,
            in3 => \N__16459\,
            lcout => \this_vga_signals.vaddress_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_9_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000011"
        )
    port map (
            in0 => \N__17169\,
            in1 => \N__20104\,
            in2 => \N__11679\,
            in3 => \N__11922\,
            lcout => this_vga_signals_vvisibility,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__16598\,
            in1 => \N__16690\,
            in2 => \_gnd_net_\,
            in3 => \N__16458\,
            lcout => OPEN,
            ltout => \this_vga_signals.un6_vvisibilitylt8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI81G42_8_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000011001"
        )
    port map (
            in0 => \N__17051\,
            in1 => \N__17168\,
            in2 => \N__11682\,
            in3 => \N__16599\,
            lcout => \this_vga_signals.vvisibility_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100110011111"
        )
    port map (
            in0 => \N__16597\,
            in1 => \N__17170\,
            in2 => \N__20114\,
            in3 => \N__17050\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m8_0_a3_1_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_0_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__12879\,
            in1 => \N__11670\,
            in2 => \N__11664\,
            in3 => \N__12949\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100010111"
        )
    port map (
            in0 => \N__16469\,
            in1 => \N__15282\,
            in2 => \N__11661\,
            in3 => \N__11658\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_a2_1_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11652\,
            in1 => \N__13383\,
            in2 => \N__11643\,
            in3 => \N__13307\,
            lcout => \this_vga_signals.g0_i_x4_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_23_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100110011111"
        )
    port map (
            in0 => \N__17166\,
            in1 => \N__16596\,
            in2 => \N__20115\,
            in3 => \N__17049\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19025\,
            in2 => \_gnd_net_\,
            in3 => \N__19102\,
            lcout => \this_vga_signals.M_vcounter_q_379_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIS6TO_9_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000101"
        )
    port map (
            in0 => \N__13938\,
            in1 => \_gnd_net_\,
            in2 => \N__14606\,
            in3 => \N__14174\,
            lcout => \this_vga_signals.SUM_3_1_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19064\,
            in2 => \N__12288\,
            in3 => \N__13980\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34555\,
            ce => 'H',
            sr => \N__12374\
        );

    \this_vga_signals.M_hcounter_q_0_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__19065\,
            in1 => \N__12283\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34555\,
            ce => 'H',
            sr => \N__12374\
        );

    \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12363\,
            in2 => \_gnd_net_\,
            in3 => \N__19055\,
            lcout => \this_vga_signals.N_692_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__14172\,
            in1 => \N__14592\,
            in2 => \_gnd_net_\,
            in3 => \N__14678\,
            lcout => this_vga_signals_hvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_RNIC68K4_9_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18282\,
            in2 => \_gnd_net_\,
            in3 => \N__34113\,
            lcout => \M_stage_q_RNIC68K4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_0_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11873\,
            lcout => \this_vga_signals.vaddress_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_20_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100110011111"
        )
    port map (
            in0 => \N__17122\,
            in1 => \N__16549\,
            in2 => \N__20092\,
            in3 => \N__17020\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m8_0_a3_1_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_18_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__11711\,
            in1 => \N__12937\,
            in2 => \N__11697\,
            in3 => \N__12862\,
            lcout => \this_vga_signals.g0_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__11871\,
            in1 => \N__12166\,
            in2 => \_gnd_net_\,
            in3 => \N__11956\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14258\,
            lcout => \this_vga_signals.M_vcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34507\,
            ce => \N__14763\,
            sr => \N__14725\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11870\,
            in2 => \_gnd_net_\,
            in3 => \N__12165\,
            lcout => \this_vga_signals.vaddress_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_1_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11872\,
            lcout => \this_vga_signals.vaddress_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_21_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100110011111"
        )
    port map (
            in0 => \N__17121\,
            in1 => \N__16550\,
            in2 => \N__20091\,
            in3 => \N__17021\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010011111100"
        )
    port map (
            in0 => \N__11982\,
            in1 => \N__11952\,
            in2 => \N__12021\,
            in3 => \N__12039\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16583\,
            in2 => \_gnd_net_\,
            in3 => \N__12852\,
            lcout => \this_vga_signals.N_5_i_0\,
            ltout => \this_vga_signals.N_5_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_0_5_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010001011"
        )
    port map (
            in0 => \N__11820\,
            in1 => \N__16743\,
            in2 => \N__11811\,
            in3 => \N__16489\,
            lcout => \this_vga_signals.g1_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14240\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34515\,
            ce => \N__14767\,
            sr => \N__14727\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__11808\,
            in1 => \N__11802\,
            in2 => \N__14814\,
            in3 => \N__11787\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100011011"
        )
    port map (
            in0 => \N__12040\,
            in1 => \N__12015\,
            in2 => \N__11997\,
            in3 => \N__11983\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011010000"
        )
    port map (
            in0 => \N__11964\,
            in1 => \N__11953\,
            in2 => \N__11925\,
            in3 => \N__11918\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111001010101"
        )
    port map (
            in0 => \N__12944\,
            in1 => \N__12581\,
            in2 => \N__11901\,
            in3 => \N__12203\,
            lcout => \this_vga_signals.mult1_un47_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIC2H0Q9_1_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110000010"
        )
    port map (
            in0 => \N__12426\,
            in1 => \N__12243\,
            in2 => \N__12093\,
            in3 => \N__13056\,
            lcout => \this_vga_signals.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_15_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010110101101"
        )
    port map (
            in0 => \N__12205\,
            in1 => \N__11886\,
            in2 => \N__12963\,
            in3 => \N__12851\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12646\,
            in1 => \N__12180\,
            in2 => \N__12604\,
            in3 => \N__12541\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__12542\,
            in1 => \_gnd_net_\,
            in2 => \N__11877\,
            in3 => \N__12712\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__11874\,
            in1 => \N__12178\,
            in2 => \_gnd_net_\,
            in3 => \N__11840\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001110"
        )
    port map (
            in0 => \N__12939\,
            in1 => \N__12589\,
            in2 => \N__11823\,
            in3 => \N__12849\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010100101"
        )
    port map (
            in0 => \N__12850\,
            in1 => \N__12943\,
            in2 => \N__12603\,
            in3 => \N__12204\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i\,
            ltout => \this_vga_signals.mult1_un54_sum_axb2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_571_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111001111000"
        )
    port map (
            in0 => \N__12179\,
            in1 => \N__12593\,
            in2 => \N__12132\,
            in3 => \N__12645\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_571\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_5_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100001110001"
        )
    port map (
            in0 => \N__16711\,
            in1 => \N__16426\,
            in2 => \N__12129\,
            in3 => \N__12114\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_2_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIOV1AF_3_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011010100"
        )
    port map (
            in0 => \N__16427\,
            in1 => \N__15275\,
            in2 => \N__12105\,
            in3 => \N__12060\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI5FISK_2_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16712\,
            in1 => \N__15396\,
            in2 => \N__12102\,
            in3 => \N__12099\,
            lcout => \this_vga_signals.g1_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__16424\,
            in1 => \N__16707\,
            in2 => \N__12081\,
            in3 => \N__12066\,
            lcout => \this_vga_signals.g0_1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_17_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__12713\,
            in1 => \N__16425\,
            in2 => \N__16742\,
            in3 => \N__12654\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0\,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIHM8LF_3_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001010101"
        )
    port map (
            in0 => \N__15298\,
            in1 => \_gnd_net_\,
            in2 => \N__12054\,
            in3 => \N__12051\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQC7Q91_2_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__15393\,
            in1 => \N__13377\,
            in2 => \N__12045\,
            in3 => \N__13293\,
            lcout => OPEN,
            ltout => \this_vga_signals.g3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_0_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001111000000"
        )
    port map (
            in0 => \N__15297\,
            in1 => \N__13211\,
            in2 => \N__12246\,
            in3 => \N__12747\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNII65L3_9_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__14597\,
            in1 => \N__14680\,
            in2 => \N__14181\,
            in3 => \N__22956\,
            lcout => \M_this_vga_ramdac_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__12280\,
            in1 => \N__12321\,
            in2 => \N__13998\,
            in3 => \N__13826\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_d7lt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__12327\,
            in1 => \N__14596\,
            in2 => \N__12237\,
            in3 => \N__14679\,
            lcout => \this_vga_signals.M_hcounter_d7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m2_0_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001001000"
        )
    port map (
            in0 => \N__14040\,
            in1 => \N__13827\,
            in2 => \N__14101\,
            in3 => \N__13463\,
            lcout => \this_vga_signals.if_m2_0\,
            ltout => \this_vga_signals.if_m2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010001001101"
        )
    port map (
            in0 => \N__13464\,
            in1 => \N__14093\,
            in2 => \N__12234\,
            in3 => \N__13830\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_0_1_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__12281\,
            in1 => \N__13088\,
            in2 => \N__13999\,
            in3 => \N__13147\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un89_sum_c3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNII3DE13_2_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110100110"
        )
    port map (
            in0 => \N__13148\,
            in1 => \N__14041\,
            in2 => \N__12231\,
            in3 => \N__13120\,
            lcout => OPEN,
            ltout => \this_vga_signals.haddress_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI7BUL75_2_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__13155\,
            in1 => \N__15558\,
            in2 => \N__12228\,
            in3 => \N__13089\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__13880\,
            in1 => \N__14158\,
            in2 => \_gnd_net_\,
            in3 => \N__13932\,
            lcout => \this_vga_signals.M_hcounter_d7lto7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14027\,
            in2 => \_gnd_net_\,
            in3 => \N__14073\,
            lcout => \this_vga_signals.un2_hsynclto3_0\,
            ltout => \this_vga_signals.un2_hsynclto3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__13990\,
            in1 => \N__12287\,
            in2 => \N__12315\,
            in3 => \N__13825\,
            lcout => OPEN,
            ltout => \this_vga_signals.un2_hsynclto6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__13881\,
            in1 => \N__14159\,
            in2 => \N__12312\,
            in3 => \N__13933\,
            lcout => \this_vga_signals.un2_hsynclt8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15618\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15817\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12282\,
            in2 => \N__13994\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19060\,
            in1 => \N__14038\,
            in2 => \_gnd_net_\,
            in3 => \N__12255\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__34556\,
            ce => 'H',
            sr => \N__12378\
        );

    \this_vga_signals.M_hcounter_q_3_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19057\,
            in1 => \N__14088\,
            in2 => \_gnd_net_\,
            in3 => \N__12252\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__34556\,
            ce => 'H',
            sr => \N__12378\
        );

    \this_vga_signals.M_hcounter_q_4_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19061\,
            in1 => \N__13824\,
            in2 => \_gnd_net_\,
            in3 => \N__12249\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__34556\,
            ce => 'H',
            sr => \N__12378\
        );

    \this_vga_signals.M_hcounter_q_5_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19058\,
            in1 => \N__13882\,
            in2 => \_gnd_net_\,
            in3 => \N__12405\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__34556\,
            ce => 'H',
            sr => \N__12378\
        );

    \this_vga_signals.M_hcounter_q_6_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19062\,
            in1 => \N__13937\,
            in2 => \_gnd_net_\,
            in3 => \N__12402\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__34556\,
            ce => 'H',
            sr => \N__12378\
        );

    \this_vga_signals.M_hcounter_q_7_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19059\,
            in1 => \N__14171\,
            in2 => \_gnd_net_\,
            in3 => \N__12399\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__34556\,
            ce => 'H',
            sr => \N__12378\
        );

    \this_vga_signals.M_hcounter_q_8_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19063\,
            in1 => \N__14671\,
            in2 => \_gnd_net_\,
            in3 => \N__12396\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__34556\,
            ce => 'H',
            sr => \N__12378\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14591\,
            in2 => \_gnd_net_\,
            in3 => \N__12393\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34567\,
            ce => \N__12390\,
            sr => \N__12373\
        );

    \this_vga_signals.un5_vaddress_g0_26_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__16477\,
            in1 => \N__12726\,
            in2 => \N__16776\,
            in3 => \N__12653\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_3_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__16478\,
            in1 => \N__12678\,
            in2 => \_gnd_net_\,
            in3 => \N__12546\,
            lcout => \this_vga_signals.g0_i_x4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_x0_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111011000011"
        )
    port map (
            in0 => \N__15263\,
            in1 => \N__12782\,
            in2 => \N__13308\,
            in3 => \N__12420\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_3_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_ns_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13389\,
            in2 => \N__12339\,
            in3 => \N__12411\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13388\,
            in1 => \N__12783\,
            in2 => \N__15291\,
            in3 => \N__13306\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_1_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__15361\,
            in1 => \N__13070\,
            in2 => \_gnd_net_\,
            in3 => \N__12738\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011101000"
        )
    port map (
            in0 => \N__15463\,
            in1 => \N__15425\,
            in2 => \N__12468\,
            in3 => \N__12465\,
            lcout => \this_vga_signals.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIMRO4P_3_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010011001"
        )
    port map (
            in0 => \N__13369\,
            in1 => \N__15234\,
            in2 => \N__12450\,
            in3 => \N__12441\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIUC6F91_1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__15405\,
            in1 => \N__15456\,
            in2 => \N__12429\,
            in3 => \N__13294\,
            lcout => \this_vga_signals.g0_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000100001"
        )
    port map (
            in0 => \N__13367\,
            in1 => \N__15230\,
            in2 => \N__12776\,
            in3 => \N__13270\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__16455\,
            in1 => \_gnd_net_\,
            in2 => \N__13296\,
            in3 => \N__15226\,
            lcout => \this_vga_signals.g0_2_0_a2_1\,
            ltout => \this_vga_signals.g0_2_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_x1_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111101101001"
        )
    port map (
            in0 => \N__12772\,
            in1 => \N__13275\,
            in2 => \N__12414\,
            in3 => \N__15235\,
            lcout => \this_vga_signals.g0_3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_13_x0_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100100111100"
        )
    port map (
            in0 => \N__12674\,
            in1 => \N__13368\,
            in2 => \N__15271\,
            in3 => \N__12538\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_13_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_13_ns_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12660\,
            in2 => \N__12741\,
            in3 => \N__13274\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010011100101"
        )
    port map (
            in0 => \N__12582\,
            in1 => \N__15225\,
            in2 => \N__16484\,
            in3 => \N__12537\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_14_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__16394\,
            in1 => \N__12732\,
            in2 => \N__16775\,
            in3 => \N__12711\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_3_d_2\,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_3_d_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_13_x1_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011000111001"
        )
    port map (
            in0 => \N__12540\,
            in1 => \N__15240\,
            in2 => \N__12663\,
            in3 => \N__13361\,
            lcout => \this_vga_signals.g0_13_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12647\,
            in2 => \N__12510\,
            in3 => \N__12615\,
            lcout => \this_vga_signals.mult1_un61_sum_c3\,
            ltout => \this_vga_signals.mult1_un61_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIANU4Q_3_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15241\,
            in2 => \N__12609\,
            in3 => \N__13362\,
            lcout => \this_vga_signals.M_vcounter_q_RNIANU4QZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x1_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010011100110"
        )
    port map (
            in0 => \N__12597\,
            in1 => \N__16366\,
            in2 => \N__15272\,
            in3 => \N__12539\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNITVMCU_3_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12501\,
            in1 => \N__13363\,
            in2 => \N__15302\,
            in3 => \N__13276\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_RNITVMCUZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI2KDQ22_3_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12495\,
            in2 => \N__12486\,
            in3 => \N__12483\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI0FHHA4_2_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111001010001"
        )
    port map (
            in0 => \N__13071\,
            in1 => \N__15387\,
            in2 => \N__13059\,
            in3 => \N__13212\,
            lcout => \this_vga_signals.g0_0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__13050\,
            in1 => \N__17068\,
            in2 => \N__13032\,
            in3 => \N__13011\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_axb1_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111001001"
        )
    port map (
            in0 => \N__12966\,
            in1 => \N__16764\,
            in2 => \N__12993\,
            in3 => \N__12801\,
            lcout => \this_vga_signals.g0_i_x4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_4_1_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011111101000"
        )
    port map (
            in0 => \N__15267\,
            in1 => \N__12768\,
            in2 => \N__16451\,
            in3 => \N__13384\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_x4_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_4_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15404\,
            in1 => \N__12990\,
            in2 => \N__12984\,
            in3 => \N__13269\,
            lcout => \this_vga_signals.g0_i_x4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_0_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100011011110"
        )
    port map (
            in0 => \N__16385\,
            in1 => \N__12965\,
            in2 => \N__16777\,
            in3 => \N__12880\,
            lcout => \this_vga_signals.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15274\,
            in1 => \N__13366\,
            in2 => \N__16481\,
            in3 => \N__13268\,
            lcout => \this_vga_signals.g0_2_0_a2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__13365\,
            in1 => \_gnd_net_\,
            in2 => \N__13295\,
            in3 => \N__12767\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_0_a2_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15273\,
            in1 => \N__13364\,
            in2 => \N__16480\,
            in3 => \N__13264\,
            lcout => \this_vga_signals.N_4_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100101100011"
        )
    port map (
            in0 => \N__13828\,
            in1 => \N__13492\,
            in2 => \N__14102\,
            in3 => \N__13465\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010011011011"
        )
    port map (
            in0 => \N__14100\,
            in1 => \N__14042\,
            in2 => \N__13197\,
            in3 => \N__13440\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI49VKF_9_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15559\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100011110"
        )
    port map (
            in0 => \N__13179\,
            in1 => \N__13172\,
            in2 => \N__13497\,
            in3 => \N__13164\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001110001"
        )
    port map (
            in0 => \N__14043\,
            in1 => \N__14000\,
            in2 => \N__13158\,
            in3 => \N__13087\,
            lcout => \this_vga_signals.mult1_un82_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIIHKHP3_9_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__15560\,
            in1 => \N__13149\,
            in2 => \N__13134\,
            in3 => \N__13121\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011001101100"
        )
    port map (
            in0 => \N__13829\,
            in1 => \N__13493\,
            in2 => \N__14103\,
            in3 => \N__13466\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010001010"
        )
    port map (
            in0 => \N__14120\,
            in1 => \N__13413\,
            in2 => \N__13884\,
            in3 => \N__13931\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13878\,
            in2 => \N__13500\,
            in3 => \N__13809\,
            lcout => \this_vga_signals.mult1_un68_sum_axb2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111110001100"
        )
    port map (
            in0 => \N__13808\,
            in1 => \N__13412\,
            in2 => \N__13883\,
            in3 => \N__13930\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14121\,
            in2 => \N__13482\,
            in3 => \N__13401\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010010"
        )
    port map (
            in0 => \N__13877\,
            in1 => \N__13395\,
            in2 => \N__13479\,
            in3 => \N__14109\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14087\,
            in2 => \N__13443\,
            in3 => \N__13810\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI18DB6_9_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13434\,
            in2 => \_gnd_net_\,
            in3 => \N__15561\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010111010111"
        )
    port map (
            in0 => \N__14663\,
            in1 => \N__14160\,
            in2 => \N__14601\,
            in3 => \N__13924\,
            lcout => \this_vga_signals.SUM_3\,
            ltout => \this_vga_signals.SUM_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000010010"
        )
    port map (
            in0 => \N__13926\,
            in1 => \N__13869\,
            in2 => \N__13404\,
            in3 => \N__13805\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__14665\,
            in1 => \N__14164\,
            in2 => \N__14602\,
            in3 => \N__13927\,
            lcout => \this_vga_signals.N_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010010101"
        )
    port map (
            in0 => \N__13925\,
            in1 => \N__14587\,
            in2 => \N__14173\,
            in3 => \N__14664\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\,
            ltout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001110"
        )
    port map (
            in0 => \N__13806\,
            in1 => \N__13879\,
            in2 => \N__14112\,
            in3 => \N__13928\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14089\,
            in1 => \N__14039\,
            in2 => \_gnd_net_\,
            in3 => \N__14001\,
            lcout => OPEN,
            ltout => \this_vga_signals.un4_hsynclt4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIFPJM1_5_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__13929\,
            in1 => \N__13870\,
            in2 => \N__13833\,
            in3 => \N__13807\,
            lcout => \this_vga_signals.un4_hsynclt8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a3_3_0_0_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__33492\,
            in1 => \N__34757\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals_N_419_i_i_0_a3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_i_2_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33443\,
            lcout => \N_91_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_i_1_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32912\,
            in2 => \_gnd_net_\,
            in3 => \N__18240\,
            lcout => \N_93_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI43UU_6_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__13740\,
            in1 => \N__29990\,
            in2 => \N__30164\,
            in3 => \N__31089\,
            lcout => \M_this_ppu_sprites_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI43UU_2_6_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__14523\,
            in1 => \N__30000\,
            in2 => \N__30162\,
            in3 => \N__31116\,
            lcout => \M_this_ppu_sprites_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18997\,
            in1 => \N__15429\,
            in2 => \N__19131\,
            in3 => \N__19123\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__34487\,
            ce => 'H',
            sr => \N__14723\
        );

    \this_vga_signals.M_vcounter_q_1_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18999\,
            in1 => \N__15457\,
            in2 => \_gnd_net_\,
            in3 => \N__14277\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__34487\,
            ce => 'H',
            sr => \N__14723\
        );

    \this_vga_signals.M_vcounter_q_2_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18998\,
            in1 => \N__15360\,
            in2 => \_gnd_net_\,
            in3 => \N__14274\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__34487\,
            ce => 'H',
            sr => \N__14723\
        );

    \this_vga_signals.M_vcounter_q_3_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19000\,
            in1 => \N__15236\,
            in2 => \_gnd_net_\,
            in3 => \N__14271\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__34487\,
            ce => 'H',
            sr => \N__14723\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16479\,
            in2 => \_gnd_net_\,
            in3 => \N__14268\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16760\,
            in2 => \_gnd_net_\,
            in3 => \N__14244\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16608\,
            in2 => \_gnd_net_\,
            in3 => \N__14208\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17072\,
            in2 => \_gnd_net_\,
            in3 => \N__14184\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17171\,
            in2 => \_gnd_net_\,
            in3 => \N__14874\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20102\,
            in2 => \_gnd_net_\,
            in3 => \N__14871\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14825\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34498\,
            ce => \N__14768\,
            sr => \N__14724\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14795\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34516\,
            ce => \N__14769\,
            sr => \N__14728\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__14690\,
            in1 => \N__14631\,
            in2 => \N__14622\,
            in3 => \N__14607\,
            lcout => this_vga_signals_hsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__15832\,
            in1 => \N__15895\,
            in2 => \N__15875\,
            in3 => \N__19113\,
            lcout => \this_vga_signals.M_pcounter_q_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_1_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__15834\,
            in1 => \N__15896\,
            in2 => \N__15876\,
            in3 => \N__19115\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34526\,
            ce => \N__19009\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_0_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__19114\,
            in1 => \N__15833\,
            in2 => \_gnd_net_\,
            in3 => \N__15714\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34526\,
            ce => \N__19009\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__15831\,
            in1 => \N__15713\,
            in2 => \_gnd_net_\,
            in3 => \N__19112\,
            lcout => \this_vga_signals.M_pcounter_q_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15805\,
            in2 => \_gnd_net_\,
            in3 => \N__16233\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_i_0_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33750\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18239\,
            lcout => \N_95_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000100110"
        )
    port map (
            in0 => \N__18730\,
            in1 => \N__18773\,
            in2 => \N__18840\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_ramdac.N_24_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__15455\,
            in1 => \N__15421\,
            in2 => \N__15365\,
            in3 => \N__15197\,
            lcout => \this_vga_signals.M_vcounter_d7lt8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI43UU_0_6_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__15150\,
            in1 => \N__29941\,
            in2 => \N__30163\,
            in3 => \N__31161\,
            lcout => \M_this_ppu_sprites_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010100101011"
        )
    port map (
            in0 => \N__18883\,
            in1 => \N__18832\,
            in2 => \N__18784\,
            in3 => \N__18729\,
            lcout => \this_vga_ramdac.m19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100101111"
        )
    port map (
            in0 => \N__18731\,
            in1 => \N__18884\,
            in2 => \N__18839\,
            in3 => \N__18777\,
            lcout => \this_vga_ramdac.m6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__14904\,
            in1 => \N__16263\,
            in2 => \N__14891\,
            in3 => \N__22870\,
            lcout => \this_vga_ramdac.N_2862_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.G_330_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15701\,
            in1 => \N__16279\,
            in2 => \_gnd_net_\,
            in3 => \N__34104\,
            lcout => \this_vga_signals.GZ0Z_330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100100101"
        )
    port map (
            in0 => \N__18871\,
            in1 => \N__18820\,
            in2 => \N__18785\,
            in3 => \N__18715\,
            lcout => \this_vga_ramdac.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__15702\,
            in1 => \N__16280\,
            in2 => \_gnd_net_\,
            in3 => \N__34105\,
            lcout => \this_pixel_clk_M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16110\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15791\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__15672\,
            in1 => \N__16255\,
            in2 => \N__15653\,
            in3 => \N__22859\,
            lcout => \this_vga_ramdac.N_2863_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__15728\,
            in1 => \_gnd_net_\,
            in2 => \N__15849\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_this_vga_signals_pixel_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__22862\,
            in1 => \N__15761\,
            in2 => \N__16266\,
            in3 => \N__15636\,
            lcout => \this_vga_ramdac.N_2867_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__15627\,
            in1 => \N__16259\,
            in2 => \N__15614\,
            in3 => \N__22861\,
            lcout => \this_vga_ramdac.N_2866_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15597\,
            in1 => \N__15845\,
            in2 => \_gnd_net_\,
            in3 => \N__15727\,
            lcout => \M_pcounter_q_ret_2_RNIH7PG8\,
            ltout => \M_pcounter_q_ret_2_RNIH7PG8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_ret_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__15790\,
            in1 => \N__15591\,
            in2 => \N__15525\,
            in3 => \N__22863\,
            lcout => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__22860\,
            in1 => \N__16109\,
            in2 => \N__16265\,
            in3 => \N__16125\,
            lcout => \this_vga_ramdac.N_2864_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI0F523_0_6_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22901\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => dma_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15897\,
            in1 => \N__15882\,
            in2 => \_gnd_net_\,
            in3 => \N__19007\,
            lcout => \this_vga_signals.N_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15874\,
            in1 => \N__15855\,
            in2 => \_gnd_net_\,
            in3 => \N__19008\,
            lcout => \this_vga_signals.N_3_0\,
            ltout => \this_vga_signals.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15837\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_pcounter_q_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15804\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15765\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15729\,
            lcout => \this_vga_signals.M_pcounter_q_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__18586\,
            in1 => \N__20463\,
            in2 => \N__16182\,
            in3 => \N__34125\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34535\,
            ce => \N__18483\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_10_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__18585\,
            in1 => \N__18280\,
            in2 => \N__16206\,
            in3 => \N__34124\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34542\,
            ce => \N__18476\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_c_0_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18339\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \M_this_data_count_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17705\,
            in2 => \N__18411\,
            in3 => \N__16149\,
            lcout => \M_this_data_count_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_0\,
            carryout => \M_this_data_count_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18428\,
            in2 => \N__17805\,
            in3 => \N__16146\,
            lcout => \M_this_data_count_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_1\,
            carryout => \M_this_data_count_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17709\,
            in2 => \N__18450\,
            in3 => \N__16143\,
            lcout => \M_this_data_count_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_2\,
            carryout => \M_this_data_count_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16947\,
            in2 => \N__17806\,
            in3 => \N__16140\,
            lcout => \M_this_data_count_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_3\,
            carryout => \M_this_data_count_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17713\,
            in2 => \N__16923\,
            in3 => \N__16137\,
            lcout => \M_this_data_count_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_4\,
            carryout => \M_this_data_count_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_6_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16965\,
            in2 => \N__17804\,
            in3 => \N__16134\,
            lcout => \M_this_data_count_q_s_6\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_5\,
            carryout => \M_this_data_count_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17714\,
            in2 => \N__16899\,
            in3 => \N__16131\,
            lcout => \M_this_data_count_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_6\,
            carryout => \M_this_data_count_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_7_THRU_LUT4_0_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16821\,
            in2 => \N__17897\,
            in3 => \N__16128\,
            lcout => \M_this_data_count_q_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => \M_this_data_count_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17817\,
            in2 => \N__17454\,
            in3 => \N__16209\,
            lcout => \M_this_data_count_q_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_8\,
            carryout => \M_this_data_count_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_10_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18386\,
            in2 => \N__17895\,
            in3 => \N__16194\,
            lcout => \M_this_data_count_q_s_10\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_9\,
            carryout => \M_this_data_count_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17810\,
            in2 => \N__18365\,
            in3 => \N__16191\,
            lcout => \M_this_data_count_q_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_10\,
            carryout => \M_this_data_count_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16860\,
            in2 => \N__17896\,
            in3 => \N__16188\,
            lcout => \M_this_data_count_q_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_11\,
            carryout => \M_this_data_count_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_13_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__16844\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16185\,
            lcout => \M_this_data_count_q_s_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_610_0_i_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__20600\,
            in1 => \N__19409\,
            in2 => \_gnd_net_\,
            in3 => \N__34109\,
            lcout => \N_610_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_i_4_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18237\,
            lcout => \N_87_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_i_7_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33657\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18238\,
            lcout => \N_81_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010101"
        )
    port map (
            in0 => \N__16611\,
            in1 => \N__16766\,
            in2 => \N__16506\,
            in3 => \N__16456\,
            lcout => \this_vga_signals.un4_lvisibility_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_7_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30152\,
            in2 => \_gnd_net_\,
            in3 => \N__34118\,
            lcout => \this_ppu.M_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16765\,
            in1 => \N__16610\,
            in2 => \N__17178\,
            in3 => \N__17047\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_d7lto8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__16502\,
            in1 => \N__20110\,
            in2 => \N__16494\,
            in3 => \N__16457\,
            lcout => \this_vga_signals.M_vcounter_d8\,
            ltout => \this_vga_signals.M_vcounter_d8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18974\,
            in2 => \N__16296\,
            in3 => \N__19119\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_0_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16281\,
            lcout => \this_pixel_clk_M_counter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34482\,
            ce => 'H',
            sr => \N__34024\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__18684\,
            in1 => \N__16264\,
            in2 => \N__16229\,
            in3 => \N__22826\,
            lcout => \this_vga_ramdac.N_2865_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIDU2V1_6_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__16794\,
            in1 => \N__16806\,
            in2 => \N__20496\,
            in3 => \N__23703\,
            lcout => OPEN,
            ltout => \dma_ac0_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI0F523_6_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16800\,
            in2 => \N__16212\,
            in3 => \N__19317\,
            lcout => dma_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_tr27_i_o3_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18306\,
            in2 => \_gnd_net_\,
            in3 => \N__35793\,
            lcout => \N_160_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIOE1S_11_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19691\,
            in1 => \N__18304\,
            in2 => \N__24965\,
            in3 => \N__20342\,
            lcout => \M_this_state_q_RNIOE1SZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un20_i_a2_x_3_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000001"
        )
    port map (
            in0 => \N__18305\,
            in1 => \N__28120\,
            in2 => \N__23750\,
            in3 => \_gnd_net_\,
            lcout => un20_i_a2_x_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIG01L_12_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__35579\,
            in1 => \N__28119\,
            in2 => \_gnd_net_\,
            in3 => \N__20410\,
            lcout => \M_this_state_q_RNIG01LZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_326_i_i_a2_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19313\,
            in2 => \_gnd_net_\,
            in3 => \N__20492\,
            lcout => \N_278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_419_i_i_0_1_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000110011"
        )
    port map (
            in0 => \N__19872\,
            in1 => \N__19395\,
            in2 => \N__19436\,
            in3 => \N__20416\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_419_i_i_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qe_0_i_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110000"
        )
    port map (
            in0 => \N__19396\,
            in1 => \N__20512\,
            in2 => \N__16788\,
            in3 => \N__34114\,
            lcout => \M_this_data_count_qe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_a3_0_9_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__33487\,
            in1 => \N__20415\,
            in2 => \N__34770\,
            in3 => \N__19871\,
            lcout => \N_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_6_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__16785\,
            in1 => \N__18568\,
            in2 => \N__19569\,
            in3 => \N__34123\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34543\,
            ce => \N__18477\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d55_9_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16964\,
            in1 => \N__16918\,
            in2 => \N__16898\,
            in3 => \N__16945\,
            lcout => \this_vga_signals.M_this_state_d55Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_4_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__16946\,
            in1 => \N__16953\,
            in2 => \_gnd_net_\,
            in3 => \N__18566\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34543\,
            ce => \N__18477\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_5_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__16932\,
            in1 => \N__18565\,
            in2 => \_gnd_net_\,
            in3 => \N__16919\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34543\,
            ce => \N__18477\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_7_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__16905\,
            in1 => \N__18567\,
            in2 => \_gnd_net_\,
            in3 => \N__16894\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34543\,
            ce => \N__18477\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_3_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__16878\,
            in1 => \N__18564\,
            in2 => \_gnd_net_\,
            in3 => \N__18449\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34543\,
            ce => \N__18477\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_11_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__18366\,
            in1 => \N__18558\,
            in2 => \_gnd_net_\,
            in3 => \N__16872\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34549\,
            ce => \N__18491\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_12_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__18559\,
            in1 => \N__16866\,
            in2 => \_gnd_net_\,
            in3 => \N__16859\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34549\,
            ce => \N__18491\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d55_8_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16858\,
            in1 => \N__17449\,
            in2 => \N__16845\,
            in3 => \N__16819\,
            lcout => \this_vga_signals.M_this_state_d55Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_8_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100001001"
        )
    port map (
            in0 => \N__16820\,
            in1 => \N__16827\,
            in2 => \N__18579\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34549\,
            ce => \N__18491\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_2_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000101"
        )
    port map (
            in0 => \N__18560\,
            in1 => \_gnd_net_\,
            in2 => \N__17469\,
            in3 => \N__18429\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34549\,
            ce => \N__18491\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_9_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__17460\,
            in1 => \N__18569\,
            in2 => \_gnd_net_\,
            in3 => \N__17453\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34557\,
            ce => \N__18498\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI43UU_1_6_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__17433\,
            in1 => \N__29978\,
            in2 => \N__30145\,
            in3 => \N__31137\,
            lcout => \M_this_ppu_sprites_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011010000"
        )
    port map (
            in0 => \N__17190\,
            in1 => \N__17177\,
            in2 => \N__20004\,
            in3 => \N__17048\,
            lcout => \this_ppu.M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIKM001_1_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__19150\,
            in1 => \N__18057\,
            in2 => \N__19227\,
            in3 => \N__18633\,
            lcout => \this_ppu.M_count_d_0_sqmuxa_1_7\,
            ltout => \this_ppu.M_count_d_0_sqmuxa_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_7_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111101001100"
        )
    port map (
            in0 => \N__25931\,
            in1 => \N__17496\,
            in2 => \N__17193\,
            in3 => \N__28642\,
            lcout => \this_ppu.M_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34475\,
            ce => 'H',
            sr => \N__34021\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011010000"
        )
    port map (
            in0 => \N__17189\,
            in1 => \N__17176\,
            in2 => \N__20000\,
            in3 => \N__17073\,
            lcout => \M_this_vga_signals_line_clk_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19191\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19151\,
            in2 => \N__17602\,
            in3 => \N__16968\,
            lcout => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17550\,
            in2 => \N__18075\,
            in3 => \N__18033\,
            lcout => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19219\,
            in2 => \N__17603\,
            in3 => \N__18030\,
            lcout => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17554\,
            in2 => \N__18120\,
            in3 => \N__18027\,
            lcout => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18137\,
            in2 => \N__17604\,
            in3 => \N__18024\,
            lcout => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17558\,
            in2 => \N__18102\,
            in3 => \N__17502\,
            lcout => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_7_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110110"
        )
    port map (
            in0 => \N__25925\,
            in1 => \N__18645\,
            in2 => \N__28668\,
            in3 => \N__17499\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_5_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000010"
        )
    port map (
            in0 => \N__19253\,
            in1 => \N__17490\,
            in2 => \N__18138\,
            in3 => \N__19288\,
            lcout => \this_ppu.M_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_6_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000010"
        )
    port map (
            in0 => \N__19254\,
            in1 => \N__17484\,
            in2 => \N__18098\,
            in3 => \N__19289\,
            lcout => \this_ppu.M_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_4_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000010"
        )
    port map (
            in0 => \N__19252\,
            in1 => \N__17478\,
            in2 => \N__19290\,
            in3 => \N__18116\,
            lcout => \this_ppu.M_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_2_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__18071\,
            in1 => \N__19284\,
            in2 => \N__18147\,
            in3 => \N__19251\,
            lcout => \this_ppu.M_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIDE0G_2_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18133\,
            in1 => \N__18115\,
            in2 => \N__18097\,
            in3 => \N__18070\,
            lcout => \this_ppu.M_count_d_1_sqmuxa_1_i_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_9_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__21023\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18666\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_i_o3_0_2_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__21678\,
            in1 => \N__21727\,
            in2 => \_gnd_net_\,
            in3 => \N__21634\,
            lcout => \N_465_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_i_o3_0_10_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21635\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19344\,
            lcout => \this_vga_signals_M_this_state_q_ns_i_o3_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18048\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__26373\,
            in1 => \N__21213\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_8_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__20865\,
            in1 => \N__23702\,
            in2 => \N__20937\,
            in3 => \N__20809\,
            lcout => \M_this_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34505\,
            ce => 'H',
            sr => \N__34012\
        );

    \this_vga_signals.un20_i_a2_sx_3_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18302\,
            in1 => \N__19338\,
            in2 => \N__19692\,
            in3 => \N__23728\,
            lcout => OPEN,
            ltout => \this_vga_signals.un20_i_a2_sxZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un20_i_a2_3_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18036\,
            in3 => \N__28118\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_11_0_i_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__19296\,
            in1 => \N__23729\,
            in2 => \N__18318\,
            in3 => \N__35713\,
            lcout => \un1_M_this_state_q_11_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_10_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100010000"
        )
    port map (
            in0 => \N__35714\,
            in1 => \N__20610\,
            in2 => \N__18315\,
            in3 => \N__18303\,
            lcout => \M_this_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34505\,
            ce => 'H',
            sr => \N__34012\
        );

    \M_this_state_q_2_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__18627\,
            in1 => \N__28567\,
            in2 => \N__24995\,
            in3 => \N__35812\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__34011\
        );

    \M_this_substate_q_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__19545\,
            in1 => \N__19526\,
            in2 => \N__18615\,
            in3 => \N__24228\,
            lcout => \M_this_substate_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__34011\
        );

    \M_this_state_q_9_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__18281\,
            in1 => \N__20519\,
            in2 => \N__18251\,
            in3 => \N__19343\,
            lcout => \M_this_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__34011\
        );

    \M_this_state_q_11_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__19668\,
            in1 => \N__19562\,
            in2 => \N__35248\,
            in3 => \N__21650\,
            lcout => \M_this_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__34011\
        );

    \M_this_state_q_5_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__35810\,
            in1 => \N__19361\,
            in2 => \N__26670\,
            in3 => \N__20420\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__34011\
        );

    \M_this_state_q_1_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__19360\,
            in1 => \N__26318\,
            in2 => \N__19527\,
            in3 => \N__35811\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__34011\
        );

    \M_this_state_q_12_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__35809\,
            in1 => \N__19667\,
            in2 => \N__21654\,
            in3 => \N__28126\,
            lcout => \M_this_state_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__34011\
        );

    \M_this_state_q_RNO_0_2_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__26725\,
            in1 => \N__19543\,
            in2 => \N__28415\,
            in3 => \N__18610\,
            lcout => \M_this_state_qc_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_1_4_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__26726\,
            in1 => \_gnd_net_\,
            in2 => \N__28416\,
            in3 => \N__18611\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001100"
        )
    port map (
            in0 => \N__35813\,
            in1 => \N__28579\,
            in2 => \N__18618\,
            in3 => \N__35578\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34524\,
            ce => 'H',
            sr => \N__34010\
        );

    \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__26727\,
            in1 => \N__28414\,
            in2 => \N__28584\,
            in3 => \N__18609\,
            lcout => \N_484_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_419_i_i_0_a2_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__21649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20579\,
            lcout => \this_vga_signals.N_279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18587\,
            in2 => \_gnd_net_\,
            in3 => \N__18338\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34533\,
            ce => \N__18484\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_1_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000101"
        )
    port map (
            in0 => \N__18588\,
            in1 => \_gnd_net_\,
            in2 => \N__18510\,
            in3 => \N__18407\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34533\,
            ce => \N__18484\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d55_6_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18445\,
            in2 => \_gnd_net_\,
            in3 => \N__18427\,
            lcout => \this_vga_signals.M_this_state_d55Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d55_7_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18403\,
            in1 => \N__18387\,
            in2 => \N__18364\,
            in3 => \N__18334\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_d55Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d55_LC_16_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18906\,
            in1 => \N__18900\,
            in2 => \N__18894\,
            in3 => \N__18891\,
            lcout => \M_this_state_d55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20988\,
            in2 => \_gnd_net_\,
            in3 => \N__21042\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110010111"
        )
    port map (
            in0 => \N__18885\,
            in1 => \N__18831\,
            in2 => \N__18789\,
            in3 => \N__18732\,
            lcout => \this_vga_ramdac.m16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_6_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20990\,
            in2 => \_gnd_net_\,
            in3 => \N__18672\,
            lcout => \this_reset_cond.M_stage_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_5_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20989\,
            in2 => \_gnd_net_\,
            in3 => \N__19740\,
            lcout => \this_reset_cond.M_stage_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_8_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__20992\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18651\,
            lcout => \this_reset_cond.M_stage_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_7_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20991\,
            in2 => \_gnd_net_\,
            in3 => \N__18657\,
            lcout => \this_reset_cond.M_stage_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIL508_7_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18644\,
            in2 => \_gnd_net_\,
            in3 => \N__19189\,
            lcout => \this_ppu.M_count_d_1_sqmuxa_1_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_0_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011111111"
        )
    port map (
            in0 => \N__29358\,
            in1 => \N__29403\,
            in2 => \N__29471\,
            in3 => \N__18921\,
            lcout => \this_ppu.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI4GQN4_0_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__29402\,
            in1 => \N__29456\,
            in2 => \_gnd_net_\,
            in3 => \N__29357\,
            lcout => \this_ppu.N_132_0\,
            ltout => \this_ppu.N_132_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_0_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000000000"
        )
    port map (
            in0 => \N__19190\,
            in1 => \N__25930\,
            in2 => \N__19194\,
            in3 => \N__18920\,
            lcout => \this_ppu.M_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__19133\,
            in1 => \N__19176\,
            in2 => \_gnd_net_\,
            in3 => \N__20147\,
            lcout => \this_vga_signals.un1_M_hcounter_d7_1_0\,
            ltout => \this_vga_signals.un1_M_hcounter_d7_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_0_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011000101010"
        )
    port map (
            in0 => \N__20133\,
            in1 => \N__19054\,
            in2 => \N__19164\,
            in3 => \N__19134\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_1_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__19152\,
            in1 => \N__19283\,
            in2 => \N__19161\,
            in3 => \N__19250\,
            lcout => \this_ppu.M_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI01PG1_0_1_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__25846\,
            in1 => \N__25921\,
            in2 => \_gnd_net_\,
            in3 => \N__34106\,
            lcout => \this_ppu.N_1157_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20132\,
            in2 => \_gnd_net_\,
            in3 => \N__19132\,
            lcout => OPEN,
            ltout => \this_vga_signals.CO0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_1_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100100000"
        )
    port map (
            in0 => \N__19053\,
            in1 => \N__18930\,
            in2 => \N__18924\,
            in3 => \N__20148\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI4HJ86_0_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__29472\,
            in1 => \N__18919\,
            in2 => \N__29434\,
            in3 => \N__29370\,
            lcout => \this_ppu.N_1157_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI4L615_0_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__29371\,
            in1 => \N__29427\,
            in2 => \N__25932\,
            in3 => \N__29473\,
            lcout => \this_ppu.un16_0\,
            ltout => \this_ppu.un16_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_3_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100100000000"
        )
    port map (
            in0 => \N__19263\,
            in1 => \N__19220\,
            in2 => \N__19257\,
            in3 => \N__19249\,
            lcout => \this_ppu.M_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__26138\,
            in1 => \N__24984\,
            in2 => \N__32971\,
            in3 => \N__35755\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_start_data_delay_out_m_0_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__23690\,
            in1 => \N__20924\,
            in2 => \N__20893\,
            in3 => \N__20801\,
            lcout => \this_vga_signals.M_this_state_q_ns_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o2_0_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__20800\,
            in1 => \_gnd_net_\,
            in2 => \N__20934\,
            in3 => \N__20885\,
            lcout => \N_459_0\,
            ltout => \N_459_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o3_0_0_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__21728\,
            in1 => \_gnd_net_\,
            in2 => \N__19200\,
            in3 => \_gnd_net_\,
            lcout => \N_462_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__20802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20881\,
            lcout => \this_start_data_delay_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__20886\,
            in1 => \N__20920\,
            in2 => \_gnd_net_\,
            in3 => \N__20799\,
            lcout => \N_458_0\,
            ltout => \N_458_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_419_i_i_0_o2_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__32954\,
            in1 => \N__20552\,
            in2 => \N__19197\,
            in3 => \N__33670\,
            lcout => \this_vga_signals.N_169_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o3_2_0_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20334\,
            in1 => \N__24961\,
            in2 => \N__35609\,
            in3 => \N__26292\,
            lcout => OPEN,
            ltout => \N_496_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_1_0_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111110101"
        )
    port map (
            in0 => \N__35716\,
            in1 => \N__19440\,
            in2 => \N__19413\,
            in3 => \N__20414\,
            lcout => OPEN,
            ltout => \M_this_state_qsr_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_0_0_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__19659\,
            in1 => \N__19410\,
            in2 => \N__19380\,
            in3 => \N__20609\,
            lcout => OPEN,
            ltout => \M_this_state_qsr_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101111100001111"
        )
    port map (
            in0 => \N__19377\,
            in1 => \N__21744\,
            in2 => \N__19371\,
            in3 => \N__21679\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34518\,
            ce => 'H',
            sr => \N__34014\
        );

    \M_this_state_q_3_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__20335\,
            in1 => \N__19368\,
            in2 => \N__26760\,
            in3 => \N__35717\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34518\,
            ce => 'H',
            sr => \N__34014\
        );

    \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_3_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23673\,
            in2 => \_gnd_net_\,
            in3 => \N__20333\,
            lcout => \this_vga_signals.N_159_0\,
            ltout => \this_vga_signals.N_159_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_12_0_m2_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__24933\,
            in1 => \N__26291\,
            in2 => \N__19347\,
            in3 => \N__35715\,
            lcout => \this_vga_signals.N_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un22_i_a2_0_o2_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19689\,
            in2 => \_gnd_net_\,
            in3 => \N__19339\,
            lcout => \N_168_0\,
            ltout => \N_168_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_2_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__20409\,
            in1 => \N__26290\,
            in2 => \N__19299\,
            in3 => \N__20270\,
            lcout => \this_vga_signals.M_this_external_address_d_0_sqmuxa_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o3_1_11_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20607\,
            in2 => \_gnd_net_\,
            in3 => \N__19690\,
            lcout => \N_456_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__32916\,
            in1 => \N__33672\,
            in2 => \N__20553\,
            in3 => \N__24199\,
            lcout => \N_500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_0_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__33800\,
            in1 => \N__27399\,
            in2 => \N__32598\,
            in3 => \N__27350\,
            lcout => \M_this_sprites_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d_2_sqmuxa_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24218\,
            in1 => \N__34740\,
            in2 => \_gnd_net_\,
            in3 => \N__24200\,
            lcout => \M_this_state_d_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a3_0_0_1_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__28407\,
            in1 => \N__26708\,
            in2 => \N__28583\,
            in3 => \N__19544\,
            lcout => \this_vga_signals_M_this_state_q_ns_0_a3_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__35781\,
            in1 => \N__22133\,
            in2 => \N__33491\,
            in3 => \N__24960\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3_0_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33799\,
            in1 => \N__32799\,
            in2 => \N__32409\,
            in3 => \N__32588\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19512\,
            in1 => \N__19491\,
            in2 => \_gnd_net_\,
            in3 => \N__30458\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30455\,
            in1 => \N__19476\,
            in2 => \_gnd_net_\,
            in3 => \N__19455\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19851\,
            in1 => \N__19833\,
            in2 => \_gnd_net_\,
            in3 => \N__30457\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30456\,
            in1 => \N__19815\,
            in2 => \_gnd_net_\,
            in3 => \N__19797\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__28999\,
            in1 => \N__24588\,
            in2 => \N__19776\,
            in3 => \N__19773\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__24589\,
            in1 => \N__19767\,
            in2 => \N__19761\,
            in3 => \N__19758\,
            lcout => \M_this_ppu_vram_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21021\,
            in2 => \_gnd_net_\,
            in3 => \N__19752\,
            lcout => \this_reset_cond.M_stage_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_4_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21022\,
            in2 => \_gnd_net_\,
            in3 => \N__19746\,
            lcout => \this_reset_cond.M_stage_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30418\,
            in1 => \N__19734\,
            in2 => \_gnd_net_\,
            in3 => \N__19716\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__29003\,
            in1 => \N__24593\,
            in2 => \N__19695\,
            in3 => \N__25038\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__24594\,
            in1 => \N__20154\,
            in2 => \N__20223\,
            in3 => \N__20631\,
            lcout => \M_this_ppu_vram_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_13_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__31002\,
            in1 => \N__30108\,
            in2 => \N__20220\,
            in3 => \N__29999\,
            lcout => \this_sprites_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30419\,
            in1 => \N__20193\,
            in2 => \_gnd_net_\,
            in3 => \N__20172\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_7_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__20622\,
            in1 => \N__25135\,
            in2 => \N__25258\,
            in3 => \N__25185\,
            lcout => \M_this_ppu_map_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34491\,
            ce => 'H',
            sr => \N__23129\
        );

    \this_ppu.M_haddress_q_5_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25243\,
            in2 => \_gnd_net_\,
            in3 => \N__20620\,
            lcout => \M_this_ppu_map_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34491\,
            ce => 'H',
            sr => \N__23129\
        );

    \this_ppu.M_haddress_q_6_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__20621\,
            in1 => \_gnd_net_\,
            in2 => \N__25257\,
            in3 => \N__25184\,
            lcout => \M_this_ppu_map_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34491\,
            ce => 'H',
            sr => \N__23129\
        );

    \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20146\,
            in1 => \N__20131\,
            in2 => \_gnd_net_\,
            in3 => \N__20109\,
            lcout => \this_vga_signals.line_clk_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_3_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__32800\,
            in1 => \N__27404\,
            in2 => \N__33658\,
            in3 => \N__27368\,
            lcout => \M_this_sprites_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_a3_0_6_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33471\,
            in1 => \N__20433\,
            in2 => \N__34705\,
            in3 => \N__19862\,
            lcout => \N_210\,
            ltout => \N_210_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_12_0_o3_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001111"
        )
    port map (
            in0 => \N__20434\,
            in1 => \_gnd_net_\,
            in2 => \N__20274\,
            in3 => \N__20354\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_167_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_12_0_i_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001111"
        )
    port map (
            in0 => \N__20435\,
            in1 => \N__20271\,
            in2 => \N__20259\,
            in3 => \N__23763\,
            lcout => \un1_M_this_state_q_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__35765\,
            in1 => \N__21168\,
            in2 => \N__25014\,
            in3 => \N__32393\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__31783\,
            in1 => \N__26357\,
            in2 => \N__32403\,
            in3 => \N__35763\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__35764\,
            in1 => \N__21427\,
            in2 => \N__25013\,
            in3 => \N__34684\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_0_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26358\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24332\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21428\,
            in2 => \_gnd_net_\,
            in3 => \N__26356\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_5_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__20256\,
            in1 => \N__27721\,
            in2 => \N__20250\,
            in3 => \N__21369\,
            lcout => \M_this_sprites_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34527\,
            ce => 'H',
            sr => \N__34017\
        );

    \M_this_sprites_address_q_6_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__27722\,
            in1 => \N__20247\,
            in2 => \N__20241\,
            in3 => \N__21135\,
            lcout => \M_this_sprites_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34527\,
            ce => 'H',
            sr => \N__34017\
        );

    \this_vga_signals.M_this_state_q_ns_i_o3_0_7_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20487\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21648\,
            lcout => OPEN,
            ltout => \this_vga_signals_M_this_state_q_ns_i_o3_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011100"
        )
    port map (
            in0 => \N__20608\,
            in1 => \N__23697\,
            in2 => \N__20556\,
            in3 => \N__35782\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34536\,
            ce => 'H',
            sr => \N__34015\
        );

    \this_vga_signals.M_this_state_d_0_sqmuxa_i_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__20429\,
            in1 => \N__20936\,
            in2 => \N__20895\,
            in3 => \N__20816\,
            lcout => \N_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d_2_sqmuxa_0_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__32917\,
            in1 => \N__33671\,
            in2 => \N__33483\,
            in3 => \N__20551\,
            lcout => \this_vga_signals_M_this_state_d_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__20488\,
            in1 => \N__20459\,
            in2 => \N__23769\,
            in3 => \N__20523\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34536\,
            ce => 'H',
            sr => \N__34015\
        );

    \this_vga_signals.un1_M_this_state_q_14_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__20458\,
            in1 => \N__20436\,
            in2 => \N__27360\,
            in3 => \N__20358\,
            lcout => \this_vga_signals.un1_M_this_state_q_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__27445\,
            in1 => \N__35779\,
            in2 => \N__32594\,
            in3 => \N__25002\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__22377\,
            in1 => \N__35780\,
            in2 => \N__33482\,
            in3 => \N__26375\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000111"
        )
    port map (
            in0 => \N__23677\,
            in1 => \N__35778\,
            in2 => \N__23767\,
            in3 => \N__20343\,
            lcout => \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20313\,
            in1 => \N__20292\,
            in2 => \_gnd_net_\,
            in3 => \N__30459\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_11_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__30081\,
            in1 => \N__30021\,
            in2 => \N__20760\,
            in3 => \N__30978\,
            lcout => \this_sprites_ram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__21048\,
            in1 => \N__30372\,
            in2 => \N__24600\,
            in3 => \N__20673\,
            lcout => \M_this_ppu_vram_data_3\,
            ltout => \M_this_ppu_vram_data_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vram_en_i_a2_0_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20708\,
            in1 => \N__21776\,
            in2 => \N__20697\,
            in3 => \N__20687\,
            lcout => \this_ppu.N_156\,
            ltout => \this_ppu.N_156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI22N1G_5_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30006\,
            in2 => \N__20676\,
            in3 => \N__23504\,
            lcout => \M_this_ppu_vram_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_6_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__23505\,
            in1 => \N__23365\,
            in2 => \N__23784\,
            in3 => \N__22871\,
            lcout => \this_ppu.M_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__24595\,
            in1 => \N__21093\,
            in2 => \N__29004\,
            in3 => \N__22995\,
            lcout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30424\,
            in1 => \N__20667\,
            in2 => \_gnd_net_\,
            in3 => \N__20649\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIRHU1G_1_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25517\,
            in1 => \N__25569\,
            in2 => \_gnd_net_\,
            in3 => \N__22605\,
            lcout => \this_ppu.un1_M_haddress_q_3_c2\,
            ltout => \this_ppu.un1_M_haddress_q_3_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI81A2G_4_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25302\,
            in1 => \N__25382\,
            in2 => \N__20625\,
            in3 => \N__25464\,
            lcout => \this_ppu.un1_M_haddress_q_3_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30423\,
            in1 => \N__21126\,
            in2 => \_gnd_net_\,
            in3 => \N__21108\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21087\,
            in1 => \N__21066\,
            in2 => \_gnd_net_\,
            in3 => \N__30425\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21030\,
            in2 => \_gnd_net_\,
            in3 => \N__20943\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21029\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIGL6V4_0_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__29474\,
            in1 => \N__29372\,
            in2 => \N__29435\,
            in3 => \N__34111\,
            lcout => \this_ppu.M_state_q_RNIGL6V4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_4_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32593\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34519\,
            ce => \N__34163\,
            sr => \N__34025\
        );

    \this_vga_signals.M_this_state_q_tr32_i_o3_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__28133\,
            in1 => \N__20935\,
            in2 => \N__20894\,
            in3 => \N__20817\,
            lcout => \N_156_0\,
            ltout => \N_156_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35435\,
            in1 => \N__34750\,
            in2 => \N__20775\,
            in3 => \N__34987\,
            lcout => \N_35_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_RNO_1_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21732\,
            in1 => \N__21689\,
            in2 => \_gnd_net_\,
            in3 => \N__21639\,
            lcout => \M_this_substate_q_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI13IA1_1_1_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__35080\,
            in1 => \N__34986\,
            in2 => \N__35467\,
            in3 => \N__34115\,
            lcout => \N_1142_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNIQ61C7_0_LC_19_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24281\,
            in2 => \N__21606\,
            in3 => \N__21605\,
            lcout => \M_this_sprites_address_q_RNIQ61C7Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_19_22_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26097\,
            in2 => \_gnd_net_\,
            in3 => \N__21591\,
            lcout => \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_0\,
            carryout => \un1_M_this_sprites_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22132\,
            in2 => \_gnd_net_\,
            in3 => \N__21588\,
            lcout => \un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_1\,
            carryout => \un1_M_this_sprites_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24038\,
            in3 => \N__21585\,
            lcout => \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_2\,
            carryout => \un1_M_this_sprites_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27466\,
            in2 => \_gnd_net_\,
            in3 => \N__21582\,
            lcout => \un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_3\,
            carryout => \un1_M_this_sprites_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21401\,
            in2 => \_gnd_net_\,
            in3 => \N__21363\,
            lcout => \un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_4\,
            carryout => \un1_M_this_sprites_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21186\,
            in3 => \N__21129\,
            lcout => \un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_5\,
            carryout => \un1_M_this_sprites_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21860\,
            in2 => \_gnd_net_\,
            in3 => \N__21765\,
            lcout => \un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_6\,
            carryout => \un1_M_this_sprites_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26433\,
            in2 => \_gnd_net_\,
            in3 => \N__21762\,
            lcout => \un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0\,
            ltout => OPEN,
            carryin => \bfn_19_23_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22373\,
            in2 => \_gnd_net_\,
            in3 => \N__21759\,
            lcout => \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_8\,
            carryout => \un1_M_this_sprites_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24688\,
            in2 => \_gnd_net_\,
            in3 => \N__21756\,
            lcout => \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_9\,
            carryout => \un1_M_this_sprites_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31861\,
            in3 => \N__21753\,
            lcout => \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_10\,
            carryout => \un1_M_this_sprites_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31940\,
            in2 => \_gnd_net_\,
            in3 => \N__21750\,
            lcout => \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_11\,
            carryout => \un1_M_this_sprites_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31724\,
            in2 => \_gnd_net_\,
            in3 => \N__21747\,
            lcout => \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_a3_5_220_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000111"
        )
    port map (
            in0 => \N__26735\,
            in1 => \N__28561\,
            in2 => \N__26666\,
            in3 => \N__28394\,
            lcout => \M_this_state_d25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_9_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22418\,
            in2 => \_gnd_net_\,
            in3 => \N__25003\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_9_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__27685\,
            in1 => \N__22587\,
            in2 => \N__22581\,
            in3 => \N__22578\,
            lcout => \M_this_sprites_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34550\,
            ce => 'H',
            sr => \N__34016\
        );

    \this_vga_signals.M_this_sprites_address_q_m_2_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22111\,
            in2 => \_gnd_net_\,
            in3 => \N__26376\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_2_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__22314\,
            in1 => \N__27683\,
            in2 => \N__22305\,
            in3 => \N__22302\,
            lcout => \M_this_sprites_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34550\,
            ce => 'H',
            sr => \N__34016\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__35851\,
            in1 => \N__24029\,
            in2 => \N__32832\,
            in3 => \N__25004\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_3_LC_19_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__27684\,
            in1 => \N__23940\,
            in2 => \N__22056\,
            in3 => \N__22053\,
            lcout => \M_this_sprites_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34550\,
            ce => 'H',
            sr => \N__34016\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__35852\,
            in1 => \N__21839\,
            in2 => \N__33818\,
            in3 => \N__26374\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_7_LC_19_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__21798\,
            in1 => \N__27702\,
            in2 => \N__22044\,
            in3 => \N__22041\,
            lcout => \M_this_sprites_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34558\,
            ce => 'H',
            sr => \N__34013\
        );

    \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21838\,
            in2 => \_gnd_net_\,
            in3 => \N__25005\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__23034\,
            in1 => \N__21792\,
            in2 => \N__24599\,
            in3 => \N__24546\,
            lcout => \M_this_ppu_vram_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_wclke_3_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31970\,
            in1 => \N__31863\,
            in2 => \N__31779\,
            in3 => \N__31649\,
            lcout => \this_sprites_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23061\,
            in1 => \N__23046\,
            in2 => \_gnd_net_\,
            in3 => \N__30460\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30464\,
            in1 => \N__23028\,
            in2 => \_gnd_net_\,
            in3 => \N__23013\,
            lcout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI42KTA_0_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100101010"
        )
    port map (
            in0 => \N__28663\,
            in1 => \N__22988\,
            in2 => \N__22930\,
            in3 => \N__34112\,
            lcout => \this_ppu.M_state_q_RNI42KTAZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_1_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__30019\,
            in1 => \N__23506\,
            in2 => \_gnd_net_\,
            in3 => \N__28664\,
            lcout => OPEN,
            ltout => \this_ppu.N_150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_1_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__23507\,
            in1 => \N__23366\,
            in2 => \N__22875\,
            in3 => \N__22872\,
            lcout => \this_ppu.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI70261_2_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__29997\,
            in1 => \N__25098\,
            in2 => \N__30082\,
            in3 => \N__25462\,
            lcout => \M_this_ppu_sprites_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_2_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__22607\,
            in1 => \N__25468\,
            in2 => \N__25580\,
            in3 => \N__25520\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34502\,
            ce => 'H',
            sr => \N__23130\
        );

    \this_ppu.M_haddress_q_1_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__25519\,
            in1 => \N__25573\,
            in2 => \_gnd_net_\,
            in3 => \N__22606\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34502\,
            ce => 'H',
            sr => \N__23130\
        );

    \this_ppu.M_haddress_q_0_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001010110"
        )
    port map (
            in0 => \N__25572\,
            in1 => \N__23508\,
            in2 => \N__30018\,
            in3 => \N__23370\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34502\,
            ce => 'H',
            sr => \N__23130\
        );

    \this_ppu.M_haddress_q_RNI88B5_0_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__28031\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25570\,
            lcout => OPEN,
            ltout => \this_ppu.un2_hscroll_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIVK7O_0_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001011"
        )
    port map (
            in0 => \N__25571\,
            in1 => \N__30055\,
            in2 => \N__23349\,
            in3 => \N__29998\,
            lcout => \M_this_ppu_sprites_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_3_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__25383\,
            in1 => \N__25463\,
            in2 => \_gnd_net_\,
            in3 => \N__23138\,
            lcout => \M_this_ppu_map_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34502\,
            ce => 'H',
            sr => \N__23130\
        );

    \this_ppu.M_haddress_q_4_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__23139\,
            in1 => \N__25384\,
            in2 => \N__25312\,
            in3 => \N__25469\,
            lcout => \M_this_ppu_map_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34502\,
            ce => 'H',
            sr => \N__23130\
        );

    \this_sprites_ram.mem_mem_3_0_wclke_3_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__31969\,
            in1 => \N__31862\,
            in2 => \N__31790\,
            in3 => \N__31645\,
            lcout => \this_sprites_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_4_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000010100000"
        )
    port map (
            in0 => \N__23393\,
            in1 => \N__23820\,
            in2 => \N__23910\,
            in3 => \N__23478\,
            lcout => \this_ppu.M_oam_idx_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_2_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010100000"
        )
    port map (
            in0 => \N__23906\,
            in1 => \N__23864\,
            in2 => \N__23456\,
            in3 => \N__23886\,
            lcout => \M_this_ppu_oam_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_1_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010100000"
        )
    port map (
            in0 => \N__30682\,
            in1 => \N__35189\,
            in2 => \N__35418\,
            in3 => \N__34982\,
            lcout => \M_this_oam_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI01PG1_1_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__25910\,
            in1 => \N__25856\,
            in2 => \_gnd_net_\,
            in3 => \N__34108\,
            lcout => \this_ppu.N_1046_0\,
            ltout => \this_ppu.N_1046_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_3_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23819\,
            in2 => \N__23511\,
            in3 => \N__23477\,
            lcout => \M_this_ppu_oam_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_0_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010000000000"
        )
    port map (
            in0 => \N__26012\,
            in1 => \N__25951\,
            in2 => \N__23420\,
            in3 => \N__23905\,
            lcout => \M_this_ppu_oam_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_5_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__34120\,
            in1 => \_gnd_net_\,
            in2 => \N__25953\,
            in3 => \N__26011\,
            lcout => \this_ppu.M_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_3_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23376\,
            in2 => \_gnd_net_\,
            in3 => \N__34119\,
            lcout => \this_ppu.M_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIGJUB2_3_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__25947\,
            in1 => \N__23413\,
            in2 => \_gnd_net_\,
            in3 => \N__26010\,
            lcout => \this_ppu.un1_M_oam_idx_q_1_c1\,
            ltout => \this_ppu.un1_M_oam_idx_q_1_c1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__23862\,
            in1 => \_gnd_net_\,
            in2 => \N__23481\,
            in3 => \N__23449\,
            lcout => \this_ppu.un1_M_oam_idx_q_1_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_RNI3VF_4_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__23448\,
            in1 => \N__23412\,
            in2 => \N__23394\,
            in3 => \N__23861\,
            lcout => \this_ppu.N_144_4\,
            ltout => \this_ppu.N_144_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_4_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__25994\,
            in1 => \N__23821\,
            in2 => \N__23379\,
            in3 => \N__34121\,
            lcout => \this_ppu.M_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_1_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__23904\,
            in1 => \N__23863\,
            in2 => \_gnd_net_\,
            in3 => \N__23885\,
            lcout => \M_this_ppu_oam_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_6_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__23825\,
            in1 => \N__23790\,
            in2 => \N__25995\,
            in3 => \N__34110\,
            lcout => \this_ppu.N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_en_iv_0_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__23768\,
            in1 => \N__23701\,
            in2 => \_gnd_net_\,
            in3 => \N__35783\,
            lcout => \M_this_sprites_ram_write_en_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__35784\,
            in1 => \N__31967\,
            in2 => \N__34761\,
            in3 => \N__26379\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_2_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__33454\,
            in1 => \N__27400\,
            in2 => \N__32389\,
            in3 => \N__27369\,
            lcout => \M_this_sprites_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__24282\,
            in1 => \N__25012\,
            in2 => \N__33833\,
            in3 => \N__35785\,
            lcout => \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_4_0_wclke_3_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31947\,
            in1 => \N__31626\,
            in2 => \N__31753\,
            in3 => \N__31845\,
            lcout => \this_sprites_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_11_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__26748\,
            in1 => \N__27725\,
            in2 => \N__24249\,
            in3 => \N__23535\,
            lcout => \M_this_sprites_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34544\,
            ce => 'H',
            sr => \N__34022\
        );

    \M_this_sprites_address_q_13_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__27727\,
            in1 => \N__23529\,
            in2 => \N__23922\,
            in3 => \N__23517\,
            lcout => \M_this_sprites_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34544\,
            ce => 'H',
            sr => \N__34022\
        );

    \M_this_sprites_address_q_12_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__24507\,
            in1 => \N__27726\,
            in2 => \N__23934\,
            in3 => \N__24501\,
            lcout => \M_this_sprites_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34544\,
            ce => 'H',
            sr => \N__34022\
        );

    \M_this_sprites_address_q_0_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__24495\,
            in1 => \N__24489\,
            in2 => \N__24483\,
            in3 => \N__27724\,
            lcout => \M_this_sprites_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34544\,
            ce => 'H',
            sr => \N__34022\
        );

    \this_vga_signals.M_this_sprites_address_q_m_11_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24985\,
            in2 => \_gnd_net_\,
            in3 => \N__31844\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_RNO_0_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__28557\,
            in1 => \N__28464\,
            in2 => \N__24648\,
            in3 => \N__24237\,
            lcout => \M_this_substate_q_s_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_8_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24986\,
            in2 => \_gnd_net_\,
            in3 => \N__26419\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_ibuf_RNIC68K4_5_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__24219\,
            in1 => \N__24204\,
            in2 => \N__34762\,
            in3 => \N__34107\,
            lcout => \N_1152_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_3_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23999\,
            in2 => \_gnd_net_\,
            in3 => \N__26384\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__24997\,
            in1 => \N__31968\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_13_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24996\,
            in2 => \_gnd_net_\,
            in3 => \N__31749\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_10_LC_20_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__24998\,
            in1 => \N__24690\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_10_LC_20_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__24654\,
            in1 => \N__27703\,
            in2 => \N__24888\,
            in3 => \N__24885\,
            lcout => \M_this_sprites_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34559\,
            ce => 'H',
            sr => \N__34018\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_20_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__24689\,
            in1 => \N__32823\,
            in2 => \N__26385\,
            in3 => \N__35850\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_RNO_3_LC_20_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__26731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28364\,
            lcout => \M_this_substate_q_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_m_4_LC_20_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27441\,
            in2 => \_gnd_net_\,
            in3 => \N__26383\,
            lcout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30453\,
            in1 => \N__24636\,
            in2 => \_gnd_net_\,
            in3 => \N__24621\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__28989\,
            in1 => \N__24587\,
            in2 => \N__24549\,
            in3 => \N__24513\,
            lcout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30454\,
            in1 => \N__24540\,
            in2 => \_gnd_net_\,
            in3 => \N__24525\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_hscroll_cry_0_c_inv_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25568\,
            in2 => \N__25113\,
            in3 => \N__28030\,
            lcout => \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_21_16_0_\,
            carryout => \this_ppu.un2_hscroll_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25502\,
            in2 => \N__25029\,
            in3 => \N__25104\,
            lcout => \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un2_hscroll_cry_0\,
            carryout => \this_ppu.un2_hscroll_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__27931\,
            in1 => \N__25461\,
            in2 => \_gnd_net_\,
            in3 => \N__25101\,
            lcout => \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_wclke_3_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__31988\,
            in1 => \N__31886\,
            in2 => \N__31799\,
            in3 => \N__31660\,
            lcout => \this_sprites_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIPG425_1_LC_21_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__28672\,
            in1 => \N__28715\,
            in2 => \_gnd_net_\,
            in3 => \N__29327\,
            lcout => \this_ppu.un1_M_vaddress_q_2_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30449\,
            in1 => \N__25068\,
            in2 => \_gnd_net_\,
            in3 => \N__25050\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30927\,
            lcout => \M_this_oam_ram_read_data_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27980\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_oam_ram_read_data_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc1_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30871\,
            in2 => \_gnd_net_\,
            in3 => \N__30928\,
            lcout => \this_ppu.un1_M_haddress_q_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI4S061_1_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__29991\,
            in1 => \N__25020\,
            in2 => \N__30153\,
            in3 => \N__25518\,
            lcout => \M_this_ppu_sprites_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28044\,
            in2 => \N__28032\,
            in3 => \N__25567\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_0\,
            ltout => OPEN,
            carryin => \bfn_21_18_0_\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27993\,
            in2 => \N__27981\,
            in3 => \N__25501\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_0\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27948\,
            in2 => \N__27936\,
            in3 => \N__25460\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_1\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27896\,
            in2 => \N__25425\,
            in3 => \N__25381\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_2\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28283\,
            in2 => \N__25347\,
            in3 => \N__25301\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_3\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28269\,
            in2 => \N__28083\,
            in3 => \N__25256\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_4\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28257\,
            in2 => \N__31056\,
            in3 => \N__25192\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_3\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_5\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25139\,
            in1 => \N__30747\,
            in2 => \N__28245\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_4\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_6\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__28227\,
            in1 => \N__28089\,
            in2 => \_gnd_net_\,
            in3 => \N__26016\,
            lcout => \this_ppu.vscroll8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_2_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__25830\,
            in1 => \N__34122\,
            in2 => \N__25926\,
            in3 => \N__26013\,
            lcout => \this_ppu.M_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34528\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35340\,
            in1 => \N__35165\,
            in2 => \N__25824\,
            in3 => \N__34994\,
            lcout => \N_48_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_28_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35341\,
            in1 => \N__35164\,
            in2 => \N__32592\,
            in3 => \N__34995\,
            lcout => \M_this_oam_ram_write_data_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_2_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__25952\,
            in1 => \N__25911\,
            in2 => \_gnd_net_\,
            in3 => \N__25857\,
            lcout => \this_ppu.N_148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_20_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32578\,
            lcout => \M_this_data_tmp_qZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34537\,
            ce => \N__31449\,
            sr => \N__34027\
        );

    \M_this_oam_address_q_RNI13IA1_0_1_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__35119\,
            in1 => \N__35400\,
            in2 => \N__35003\,
            in3 => \N__34116\,
            lcout => \N_1134_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__26434\,
            in1 => \N__26378\,
            in2 => \N__32985\,
            in3 => \N__35787\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d21_6_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28527\,
            in1 => \N__28214\,
            in2 => \N__28167\,
            in3 => \N__28191\,
            lcout => \this_vga_signals.M_this_state_d21Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_5_0_wclke_3_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31627\,
            in1 => \N__31948\,
            in2 => \N__31754\,
            in3 => \N__31846\,
            lcout => \this_sprites_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d22_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__28502\,
            in1 => \N__28395\,
            in2 => \N__26682\,
            in3 => \N__28454\,
            lcout => \M_this_state_d22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__31843\,
            in1 => \N__26377\,
            in2 => \N__32568\,
            in3 => \N__35846\,
            lcout => \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d24_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26739\,
            in1 => \N__26681\,
            in2 => \N__28329\,
            in3 => \N__28503\,
            lcout => \this_vga_signals.M_this_state_dZ0Z24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_9_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__35610\,
            in1 => \N__32019\,
            in2 => \N__35871\,
            in3 => \N__32926\,
            lcout => \M_this_external_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34560\,
            ce => 'H',
            sr => \N__34023\
        );

    \M_this_sprites_address_q_8_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__27729\,
            in1 => \N__26640\,
            in2 => \N__26631\,
            in3 => \N__26622\,
            lcout => \M_this_sprites_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34560\,
            ce => 'H',
            sr => \N__34023\
        );

    \this_vga_signals.M_this_sprites_address_q_m_1_LC_21_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26044\,
            in2 => \_gnd_net_\,
            in3 => \N__26352\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_q_mZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_1_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__26250\,
            in1 => \N__27728\,
            in2 => \N__26238\,
            in3 => \N__26235\,
            lcout => \M_this_sprites_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34560\,
            ce => 'H',
            sr => \N__34023\
        );

    \M_this_sprites_address_q_4_LC_21_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__27738\,
            in1 => \N__27723\,
            in2 => \N__27654\,
            in3 => \N__27645\,
            lcout => \M_this_sprites_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34568\,
            ce => 'H',
            sr => \N__34020\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_1_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__32955\,
            in1 => \N__27405\,
            in2 => \N__34739\,
            in3 => \N__27361\,
            lcout => \M_this_sprites_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_7_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34493\,
            ce => \N__34198\,
            sr => \N__34036\
        );

    \this_ppu.M_state_q_RNI53UU_6_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__27222\,
            in1 => \N__30017\,
            in2 => \N__31041\,
            in3 => \N__30112\,
            lcout => \M_this_ppu_sprites_addr_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__30016\,
            in1 => \N__29040\,
            in2 => \N__30136\,
            in3 => \N__28711\,
            lcout => \M_this_ppu_sprites_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_1_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__29326\,
            in1 => \_gnd_net_\,
            in2 => \N__28721\,
            in3 => \N__28676\,
            lcout => \this_ppu.M_vaddress_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34503\,
            ce => 'H',
            sr => \N__29264\
        );

    \this_ppu.M_vaddress_q_5_LC_22_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27851\,
            lcout => \M_this_ppu_map_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34503\,
            ce => 'H',
            sr => \N__29264\
        );

    \this_ppu.M_vaddress_q_6_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27882\,
            in1 => \N__27801\,
            in2 => \_gnd_net_\,
            in3 => \N__27852\,
            lcout => \M_this_ppu_map_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34503\,
            ce => 'H',
            sr => \N__29264\
        );

    \this_ppu.M_vaddress_q_7_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__27853\,
            in1 => \N__27880\,
            in2 => \N__27809\,
            in3 => \N__27760\,
            lcout => \M_this_ppu_map_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34503\,
            ce => 'H',
            sr => \N__29264\
        );

    \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_22_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29506\,
            in1 => \N__29556\,
            in2 => \N__29594\,
            in3 => \N__29630\,
            lcout => \this_ppu.un1_M_vaddress_q_2_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29213\,
            in2 => \N__29198\,
            in3 => \N__29302\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_7\,
            ltout => OPEN,
            carryin => \bfn_22_17_0_\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29147\,
            in2 => \N__31206\,
            in3 => \N__28716\,
            lcout => \this_ppu.M_vaddress_q_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_0\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29132\,
            in2 => \N__29118\,
            in3 => \N__29628\,
            lcout => \this_ppu.M_vaddress_q_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_1\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30332\,
            in2 => \N__31509\,
            in3 => \N__29555\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_2\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30314\,
            in2 => \N__30945\,
            in3 => \N__29505\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_6\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_3\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30296\,
            in2 => \N__31221\,
            in3 => \N__27857\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_7\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_4\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30278\,
            in2 => \N__31347\,
            in3 => \N__27808\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_8\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_5\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31392\,
            in2 => \N__30264\,
            in3 => \N__27764\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_9\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_6\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28092\,
            lcout => \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc2_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__30782\,
            in1 => \N__30879\,
            in2 => \_gnd_net_\,
            in3 => \N__30930\,
            lcout => \this_ppu.un1_M_haddress_q_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNO_0_4_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35398\,
            in1 => \N__35175\,
            in2 => \N__34996\,
            in3 => \N__30590\,
            lcout => OPEN,
            ltout => \un1_M_this_oam_address_q_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_4_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__30689\,
            in1 => \N__30181\,
            in2 => \N__28071\,
            in3 => \N__30634\,
            lcout => \M_this_oam_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35397\,
            in1 => \N__35174\,
            in2 => \N__28068\,
            in3 => \N__34922\,
            lcout => \N_65_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_0_c_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28043\,
            in2 => \N__28026\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_19_0_\,
            carryout => \this_ppu.un1_M_haddress_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_1_c_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27992\,
            in2 => \N__27976\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_0\,
            carryout => \this_ppu.un1_M_haddress_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_2_c_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27947\,
            in2 => \N__27932\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_1\,
            carryout => \this_ppu.un1_M_haddress_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_3_c_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30929\,
            in2 => \N__27897\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_2\,
            carryout => \this_ppu.un1_M_haddress_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_4_c_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30878\,
            in2 => \N__28284\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_3\,
            carryout => \this_ppu.un1_M_haddress_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_5_c_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28268\,
            in2 => \N__30786\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_4\,
            carryout => \this_ppu.un1_M_haddress_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_6_c_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28256\,
            in2 => \N__30819\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_5\,
            carryout => \this_ppu.un1_M_haddress_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_7_c_LC_22_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28241\,
            in2 => \N__30840\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_6\,
            carryout => \this_ppu.un1_M_haddress_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__30957\,
            in1 => \N__31068\,
            in2 => \N__30243\,
            in3 => \N__28230\,
            lcout => \this_ppu.vscroll8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_2_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__30585\,
            in1 => \N__30683\,
            in2 => \_gnd_net_\,
            in3 => \N__30552\,
            lcout => \M_this_oam_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d21_6_x_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__28221\,
            in1 => \N__28187\,
            in2 => \_gnd_net_\,
            in3 => \N__28160\,
            lcout => \M_this_state_d21_6_x\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNILT531_12_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34935\,
            in1 => \N__28137\,
            in2 => \N__35469\,
            in3 => \N__35786\,
            lcout => \un1_M_this_oam_address_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_13_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35452\,
            in1 => \N__35098\,
            in2 => \N__28593\,
            in3 => \N__34936\,
            lcout => \N_56_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_13_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34695\,
            lcout => \M_this_data_tmp_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34561\,
            ce => \N__32188\,
            sr => \N__34026\
        );

    \this_vga_signals.M_this_state_d21_1_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__28501\,
            in1 => \N__28478\,
            in2 => \N__28455\,
            in3 => \N__28520\,
            lcout => \M_this_state_d21_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_RNO_2_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__28519\,
            in1 => \N__28500\,
            in2 => \N__28479\,
            in3 => \N__28450\,
            lcout => \M_this_substate_q_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d24_1_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__28441\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28382\,
            lcout => \this_vga_signals.M_this_state_d24Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_7_0_wclke_3_LC_22_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__31983\,
            in1 => \N__31875\,
            in2 => \N__31791\,
            in3 => \N__31659\,
            lcout => \this_sprites_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_3_LC_22_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32801\,
            lcout => \M_this_data_tmp_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34581\,
            ce => \N__34187\,
            sr => \N__34019\
        );

    \M_this_data_tmp_q_esr_15_LC_23_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33629\,
            lcout => \M_this_data_tmp_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34494\,
            ce => \N__32189\,
            sr => \N__34039\
        );

    \M_this_data_tmp_q_esr_6_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34504\,
            ce => \N__34199\,
            sr => \N__34037\
        );

    \this_vga_signals.M_this_oam_ram_write_data_15_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35466\,
            in1 => \N__35230\,
            in2 => \N__29076\,
            in3 => \N__34962\,
            lcout => \M_this_oam_ram_write_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_vscroll_cry_0_c_inv_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29303\,
            in2 => \N__29049\,
            in3 => \N__29199\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_16\,
            ltout => OPEN,
            carryin => \bfn_23_16_0_\,
            carryout => \this_ppu.un2_vscroll_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31167\,
            in2 => \N__28722\,
            in3 => \N__29034\,
            lcout => \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un2_vscroll_cry_0\,
            carryout => \this_ppu.un2_vscroll_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__29116\,
            in1 => \N__29629\,
            in2 => \_gnd_net_\,
            in3 => \N__29031\,
            lcout => \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_12_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__30161\,
            in1 => \N__30020\,
            in2 => \N__29028\,
            in3 => \N__31020\,
            lcout => \this_sprites_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__30002\,
            in1 => \N__28956\,
            in2 => \N__30165\,
            in3 => \N__29631\,
            lcout => \M_this_ppu_sprites_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_2_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__29633\,
            in1 => \N__28720\,
            in2 => \N__28677\,
            in3 => \N__29306\,
            lcout => \this_ppu.M_vaddress_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34530\,
            ce => 'H',
            sr => \N__29265\
        );

    \this_ppu.M_vaddress_q_3_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29600\,
            in1 => \N__29557\,
            in2 => \_gnd_net_\,
            in3 => \N__29632\,
            lcout => \M_this_ppu_map_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34530\,
            ce => 'H',
            sr => \N__29265\
        );

    \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29193\,
            in2 => \_gnd_net_\,
            in3 => \N__29304\,
            lcout => OPEN,
            ltout => \this_ppu.un2_vscroll_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIS5A21_0_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001101"
        )
    port map (
            in0 => \N__30160\,
            in1 => \N__29319\,
            in2 => \N__30024\,
            in3 => \N__30001\,
            lcout => \M_this_ppu_sprites_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_4_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__29634\,
            in1 => \N__29601\,
            in2 => \N__29564\,
            in3 => \N__29507\,
            lcout => \M_this_ppu_map_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34530\,
            ce => 'H',
            sr => \N__29265\
        );

    \this_ppu.M_vaddress_q_0_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010011010101010"
        )
    port map (
            in0 => \N__29305\,
            in1 => \N__29481\,
            in2 => \N__29436\,
            in3 => \N__29379\,
            lcout => \M_this_ppu_vram_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34530\,
            ce => 'H',
            sr => \N__29265\
        );

    \M_this_oam_address_q_0_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__34921\,
            in1 => \_gnd_net_\,
            in2 => \N__35229\,
            in3 => \N__30690\,
            lcout => \M_this_oam_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35399\,
            in1 => \N__35176\,
            in2 => \N__29241\,
            in3 => \N__34920\,
            lcout => \N_71_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_0_c_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29214\,
            in2 => \N__29197\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_23_19_0_\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_1_c_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29148\,
            in2 => \N__31205\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_0\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_2_c_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29133\,
            in2 => \N__29117\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_1\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_3_c_LC_23_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31545\,
            in2 => \N__30336\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_2\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_4_c_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31257\,
            in2 => \N__30318\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_3\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_5_c_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31290\,
            in2 => \N__30300\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_4\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_6_c_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31373\,
            in2 => \N__30282\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_5\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_7_c_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30263\,
            in2 => \N__31416\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_6\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30246\,
            lcout => \this_ppu.un1_M_vaddress_q_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_10_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35430\,
            in1 => \N__35169\,
            in2 => \N__30501\,
            in3 => \N__34937\,
            lcout => \N_61_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34938\,
            in1 => \N__30222\,
            in2 => \N__35228\,
            in3 => \N__35444\,
            lcout => \N_73_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_5_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010100000"
        )
    port map (
            in0 => \N__30685\,
            in1 => \N__30191\,
            in2 => \N__30710\,
            in3 => \N__30537\,
            lcout => \M_this_oam_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_3_LC_23_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__30551\,
            in1 => \N__30586\,
            in2 => \N__30635\,
            in3 => \N__30684\,
            lcout => \M_this_oam_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNO_0_5_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30621\,
            in1 => \N__30581\,
            in2 => \_gnd_net_\,
            in3 => \N__30550\,
            lcout => \un1_M_this_oam_address_q_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_19_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35445\,
            in1 => \N__35170\,
            in2 => \N__31488\,
            in3 => \N__34939\,
            lcout => \N_50_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_21_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35431\,
            in1 => \N__35120\,
            in2 => \N__30510\,
            in3 => \N__34950\,
            lcout => \N_46_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_21_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34706\,
            lcout => \M_this_data_tmp_qZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34562\,
            ce => \N__31445\,
            sr => \N__34029\
        );

    \M_this_data_tmp_q_esr_10_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33444\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34569\,
            ce => \N__32183\,
            sr => \N__34028\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30489\,
            in1 => \N__30477\,
            in2 => \_gnd_net_\,
            in3 => \N__30465\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__31989\,
            in1 => \N__31890\,
            in2 => \N__31800\,
            in3 => \N__31671\,
            lcout => \this_sprites_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31201\,
            lcout => \M_this_oam_ram_read_data_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un9lto7_5_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31148\,
            in1 => \N__31127\,
            in2 => \N__31109\,
            in3 => \N__31079\,
            lcout => \this_ppu.un9lto7Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc3_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__30774\,
            in1 => \N__30870\,
            in2 => \N__30815\,
            in3 => \N__30915\,
            lcout => \this_ppu.un1_M_haddress_q_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un9lto7_4_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31031\,
            in1 => \N__31013\,
            in2 => \N__30995\,
            in3 => \N__30968\,
            lcout => \this_ppu.un9lto7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc1_LC_24_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__31541\,
            in1 => \_gnd_net_\,
            in2 => \N__31256\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.un1_M_vaddress_q_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_ac0_1_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30905\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30861\,
            lcout => OPEN,
            ltout => \this_ppu.un1_oam_data_1_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc4_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__30830\,
            in1 => \N__30811\,
            in2 => \N__30789\,
            in3 => \N__30775\,
            lcout => \this_ppu.un1_M_haddress_q_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_24_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35439\,
            in1 => \N__35184\,
            in2 => \N__30738\,
            in3 => \N__34923\,
            lcout => \N_67_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_ac0_1_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31249\,
            in2 => \_gnd_net_\,
            in3 => \N__31540\,
            lcout => OPEN,
            ltout => \this_ppu.un1_oam_data_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc4_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__31415\,
            in1 => \N__31374\,
            in2 => \N__31395\,
            in3 => \N__31289\,
            lcout => \this_ppu.un1_M_vaddress_q_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_22_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34892\,
            in1 => \N__31470\,
            in2 => \N__35233\,
            in3 => \N__35423\,
            lcout => \M_this_oam_ram_write_data_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc3_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__31248\,
            in1 => \N__31282\,
            in2 => \N__31372\,
            in3 => \N__31536\,
            lcout => \this_ppu.un1_M_vaddress_q_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_31_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34890\,
            in1 => \N__33668\,
            in2 => \N__35231\,
            in3 => \N__35421\,
            lcout => \M_this_oam_ram_write_data_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_18_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35420\,
            in1 => \N__35200\,
            in2 => \N__31479\,
            in3 => \N__34893\,
            lcout => \N_52_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_16_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34891\,
            in1 => \N__31494\,
            in2 => \N__35232\,
            in3 => \N__35422\,
            lcout => \M_this_oam_ram_write_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o3_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35419\,
            in1 => \N__35190\,
            in2 => \_gnd_net_\,
            in3 => \N__34889\,
            lcout => \N_158_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc2_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__31535\,
            in1 => \N__31278\,
            in2 => \_gnd_net_\,
            in3 => \N__31247\,
            lcout => \this_ppu.un1_M_vaddress_q_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31534\,
            lcout => \M_this_oam_ram_read_data_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_16_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33825\,
            lcout => \M_this_data_tmp_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34563\,
            ce => \N__31438\,
            sr => \N__34031\
        );

    \M_this_data_tmp_q_esr_19_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34563\,
            ce => \N__31438\,
            sr => \N__34031\
        );

    \M_this_data_tmp_q_esr_18_LC_24_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33472\,
            lcout => \M_this_data_tmp_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34563\,
            ce => \N__31438\,
            sr => \N__34031\
        );

    \M_this_data_tmp_q_esr_22_LC_24_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32331\,
            lcout => \M_this_data_tmp_qZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34563\,
            ce => \N__31438\,
            sr => \N__34031\
        );

    \M_this_data_tmp_q_esr_23_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33669\,
            lcout => \M_this_data_tmp_qZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34563\,
            ce => \N__31438\,
            sr => \N__34031\
        );

    \M_this_data_tmp_q_esr_17_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32981\,
            lcout => \M_this_data_tmp_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34563\,
            ce => \N__31438\,
            sr => \N__34031\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35429\,
            in1 => \N__35122\,
            in2 => \N__31464\,
            in3 => \N__34953\,
            lcout => \N_54_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI13IA1_1_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__34951\,
            in1 => \N__35427\,
            in2 => \N__35183\,
            in3 => \N__34117\,
            lcout => \N_1126_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_30_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35428\,
            in1 => \N__35121\,
            in2 => \N__32352\,
            in3 => \N__34952\,
            lcout => \M_this_oam_ram_write_data_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_0_c_LC_24_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33296\,
            in2 => \N__33272\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_24_22_0_\,
            carryout => \un1_M_this_external_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_0_THRU_LUT4_0_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33222\,
            in2 => \_gnd_net_\,
            in3 => \N__31566\,
            lcout => \un1_M_this_external_address_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_0\,
            carryout => \un1_M_this_external_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_1_THRU_LUT4_0_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33173\,
            in2 => \_gnd_net_\,
            in3 => \N__31563\,
            lcout => \un1_M_this_external_address_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_1\,
            carryout => \un1_M_this_external_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_2_THRU_LUT4_0_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33125\,
            in2 => \_gnd_net_\,
            in3 => \N__31560\,
            lcout => \un1_M_this_external_address_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_2\,
            carryout => \un1_M_this_external_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_3_THRU_LUT4_0_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33084\,
            in2 => \_gnd_net_\,
            in3 => \N__31557\,
            lcout => \un1_M_this_external_address_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_3\,
            carryout => \un1_M_this_external_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_4_THRU_LUT4_0_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33038\,
            in2 => \_gnd_net_\,
            in3 => \N__31554\,
            lcout => \un1_M_this_external_address_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_4\,
            carryout => \un1_M_this_external_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_5_THRU_LUT4_0_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35519\,
            in2 => \_gnd_net_\,
            in3 => \N__31551\,
            lcout => \un1_M_this_external_address_q_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_5\,
            carryout => \un1_M_this_external_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_6_THRU_LUT4_0_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32635\,
            in2 => \_gnd_net_\,
            in3 => \N__31548\,
            lcout => \un1_M_this_external_address_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_6\,
            carryout => \un1_M_this_external_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33695\,
            in2 => \_gnd_net_\,
            in3 => \N__32046\,
            lcout => \un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0\,
            ltout => OPEN,
            carryin => \bfn_24_23_0_\,
            carryout => \un1_M_this_external_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32033\,
            in2 => \_gnd_net_\,
            in3 => \N__32010\,
            lcout => \un1_M_this_external_address_q_cry_8_c_RNI09PBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_8\,
            carryout => \un1_M_this_external_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33317\,
            in2 => \_gnd_net_\,
            in3 => \N__32007\,
            lcout => \un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_9\,
            carryout => \un1_M_this_external_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32684\,
            in2 => \_gnd_net_\,
            in3 => \N__32004\,
            lcout => \un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_10\,
            carryout => \un1_M_this_external_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32480\,
            in2 => \_gnd_net_\,
            in3 => \N__32001\,
            lcout => \un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_11\,
            carryout => \un1_M_this_external_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32444\,
            in2 => \_gnd_net_\,
            in3 => \N__31998\,
            lcout => \un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_12\,
            carryout => \un1_M_this_external_address_q_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32270\,
            in2 => \_gnd_net_\,
            in3 => \N__31995\,
            lcout => \un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_13\,
            carryout => \un1_M_this_external_address_q_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33524\,
            in2 => \_gnd_net_\,
            in3 => \N__31992\,
            lcout => \un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__31984\,
            in1 => \N__31885\,
            in2 => \N__31795\,
            in3 => \N__31667\,
            lcout => \this_sprites_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_8_LC_26_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35247\,
            in1 => \N__35483\,
            in2 => \N__32109\,
            in3 => \N__35002\,
            lcout => \M_this_oam_ram_write_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_8_LC_26_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34548\,
            ce => \N__32184\,
            sr => \N__34040\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_26_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35486\,
            in1 => \N__35239\,
            in2 => \N__32094\,
            in3 => \N__34990\,
            lcout => \N_79_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_0_LC_26_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34552\,
            ce => \N__34200\,
            sr => \N__34038\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_26_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35484\,
            in1 => \N__35246\,
            in2 => \N__35004\,
            in3 => \N__33814\,
            lcout => \N_43_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_26_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34988\,
            in1 => \N__32064\,
            in2 => \N__35250\,
            in3 => \N__35485\,
            lcout => \N_77_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_1_LC_26_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32987\,
            lcout => \M_this_data_tmp_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34552\,
            ce => \N__34200\,
            sr => \N__34038\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_26_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34989\,
            in1 => \N__32220\,
            in2 => \N__35249\,
            in3 => \N__35487\,
            lcout => \N_58_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_14_LC_26_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35441\,
            in1 => \N__35186\,
            in2 => \N__32202\,
            in3 => \N__34980\,
            lcout => \M_this_oam_ram_write_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_26_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34978\,
            in1 => \N__35443\,
            in2 => \N__32211\,
            in3 => \N__35188\,
            lcout => \N_63_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_26_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35442\,
            in1 => \N__35187\,
            in2 => \N__32859\,
            in3 => \N__34981\,
            lcout => \N_75_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_11_LC_26_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35440\,
            in1 => \N__35185\,
            in2 => \N__32229\,
            in3 => \N__34979\,
            lcout => \M_this_oam_ram_write_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_11_LC_26_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32831\,
            lcout => \M_this_data_tmp_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34570\,
            ce => \N__32190\,
            sr => \N__34034\
        );

    \M_this_data_tmp_q_esr_12_LC_26_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34570\,
            ce => \N__32190\,
            sr => \N__34034\
        );

    \M_this_data_tmp_q_esr_9_LC_26_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32988\,
            lcout => \M_this_data_tmp_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34570\,
            ce => \N__32190\,
            sr => \N__34034\
        );

    \M_this_data_tmp_q_esr_14_LC_26_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32388\,
            lcout => \M_this_data_tmp_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34570\,
            ce => \N__32190\,
            sr => \N__34034\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_26_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35237\,
            in1 => \N__35481\,
            in2 => \N__33421\,
            in3 => \N__35001\,
            lcout => \N_39_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_27_LC_26_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35235\,
            in1 => \N__35480\,
            in2 => \N__32830\,
            in3 => \N__35000\,
            lcout => \M_this_oam_ram_write_data_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_23_LC_26_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35234\,
            in1 => \N__35479\,
            in2 => \N__33006\,
            in3 => \N__34999\,
            lcout => \M_this_oam_ram_write_data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_26_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34998\,
            in1 => \N__35482\,
            in2 => \N__32986\,
            in3 => \N__35236\,
            lcout => \N_41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_2_LC_26_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33394\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34576\,
            ce => \N__34162\,
            sr => \N__34033\
        );

    \M_this_external_address_q_11_LC_26_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__35634\,
            in1 => \N__32847\,
            in2 => \N__32834\,
            in3 => \N__35856\,
            lcout => \M_this_external_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__34032\
        );

    \M_this_external_address_q_7_LC_26_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__35855\,
            in1 => \N__35640\,
            in2 => \N__32636\,
            in3 => \N__32661\,
            lcout => \M_this_external_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__34032\
        );

    \M_this_external_address_q_12_LC_26_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__35635\,
            in1 => \N__32610\,
            in2 => \N__32547\,
            in3 => \N__35857\,
            lcout => \M_this_external_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__34032\
        );

    \M_this_external_address_q_13_LC_26_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35853\,
            in1 => \N__35638\,
            in2 => \N__34694\,
            in3 => \N__32457\,
            lcout => \M_this_external_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__34032\
        );

    \M_this_external_address_q_14_LC_26_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__35636\,
            in1 => \N__32421\,
            in2 => \N__32407\,
            in3 => \N__35858\,
            lcout => \M_this_external_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__34032\
        );

    \M_this_external_address_q_8_LC_26_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__35637\,
            in1 => \N__33846\,
            in2 => \N__33834\,
            in3 => \N__35859\,
            lcout => \M_this_external_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__34032\
        );

    \M_this_external_address_q_15_LC_26_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35854\,
            in1 => \N__35639\,
            in2 => \N__33637\,
            in3 => \N__33546\,
            lcout => \M_this_external_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__34032\
        );

    \M_this_external_address_q_10_LC_26_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__35611\,
            in1 => \N__33501\,
            in2 => \N__33420\,
            in3 => \N__35864\,
            lcout => \M_this_external_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__34030\
        );

    \M_this_external_address_q_0_LC_26_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__35860\,
            in1 => \N__35615\,
            in2 => \N__33262\,
            in3 => \N__33303\,
            lcout => \M_this_external_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__34030\
        );

    \M_this_external_address_q_1_LC_26_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000111100"
        )
    port map (
            in0 => \N__35612\,
            in1 => \N__33234\,
            in2 => \N__33220\,
            in3 => \N__35865\,
            lcout => \M_this_external_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__34030\
        );

    \M_this_external_address_q_2_LC_26_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__35861\,
            in1 => \N__35616\,
            in2 => \N__33172\,
            in3 => \N__33192\,
            lcout => \M_this_external_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__34030\
        );

    \M_this_external_address_q_3_LC_26_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000111100"
        )
    port map (
            in0 => \N__35613\,
            in1 => \N__33144\,
            in2 => \N__33124\,
            in3 => \N__35866\,
            lcout => \M_this_external_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__34030\
        );

    \M_this_external_address_q_4_LC_26_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__35862\,
            in1 => \N__35617\,
            in2 => \N__33082\,
            in3 => \N__33096\,
            lcout => \M_this_external_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__34030\
        );

    \M_this_external_address_q_5_LC_26_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000111100"
        )
    port map (
            in0 => \N__35614\,
            in1 => \N__33054\,
            in2 => \N__33034\,
            in3 => \N__35867\,
            lcout => \M_this_external_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__34030\
        );

    \M_this_external_address_q_6_LC_26_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__35863\,
            in1 => \N__35618\,
            in2 => \N__35515\,
            in3 => \N__35538\,
            lcout => \M_this_external_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__34030\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_27_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35468\,
            in1 => \N__35238\,
            in2 => \N__34605\,
            in3 => \N__34997\,
            lcout => \N_69_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_5_LC_27_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34664\,
            lcout => \M_this_data_tmp_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34577\,
            ce => \N__34188\,
            sr => \N__34035\
        );
end \INTERFACE\;
