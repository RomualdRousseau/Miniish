// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 30 2022 08:36:04

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    led,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output [7:0] led;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__35922;
    wire N__35921;
    wire N__35920;
    wire N__35911;
    wire N__35910;
    wire N__35909;
    wire N__35902;
    wire N__35901;
    wire N__35900;
    wire N__35893;
    wire N__35892;
    wire N__35891;
    wire N__35884;
    wire N__35883;
    wire N__35882;
    wire N__35875;
    wire N__35874;
    wire N__35873;
    wire N__35866;
    wire N__35865;
    wire N__35864;
    wire N__35857;
    wire N__35856;
    wire N__35855;
    wire N__35848;
    wire N__35847;
    wire N__35846;
    wire N__35839;
    wire N__35838;
    wire N__35837;
    wire N__35830;
    wire N__35829;
    wire N__35828;
    wire N__35821;
    wire N__35820;
    wire N__35819;
    wire N__35812;
    wire N__35811;
    wire N__35810;
    wire N__35803;
    wire N__35802;
    wire N__35801;
    wire N__35794;
    wire N__35793;
    wire N__35792;
    wire N__35785;
    wire N__35784;
    wire N__35783;
    wire N__35776;
    wire N__35775;
    wire N__35774;
    wire N__35767;
    wire N__35766;
    wire N__35765;
    wire N__35758;
    wire N__35757;
    wire N__35756;
    wire N__35749;
    wire N__35748;
    wire N__35747;
    wire N__35740;
    wire N__35739;
    wire N__35738;
    wire N__35731;
    wire N__35730;
    wire N__35729;
    wire N__35722;
    wire N__35721;
    wire N__35720;
    wire N__35713;
    wire N__35712;
    wire N__35711;
    wire N__35704;
    wire N__35703;
    wire N__35702;
    wire N__35695;
    wire N__35694;
    wire N__35693;
    wire N__35686;
    wire N__35685;
    wire N__35684;
    wire N__35677;
    wire N__35676;
    wire N__35675;
    wire N__35668;
    wire N__35667;
    wire N__35666;
    wire N__35659;
    wire N__35658;
    wire N__35657;
    wire N__35650;
    wire N__35649;
    wire N__35648;
    wire N__35641;
    wire N__35640;
    wire N__35639;
    wire N__35632;
    wire N__35631;
    wire N__35630;
    wire N__35623;
    wire N__35622;
    wire N__35621;
    wire N__35614;
    wire N__35613;
    wire N__35612;
    wire N__35605;
    wire N__35604;
    wire N__35603;
    wire N__35596;
    wire N__35595;
    wire N__35594;
    wire N__35587;
    wire N__35586;
    wire N__35585;
    wire N__35578;
    wire N__35577;
    wire N__35576;
    wire N__35569;
    wire N__35568;
    wire N__35567;
    wire N__35560;
    wire N__35559;
    wire N__35558;
    wire N__35551;
    wire N__35550;
    wire N__35549;
    wire N__35542;
    wire N__35541;
    wire N__35540;
    wire N__35533;
    wire N__35532;
    wire N__35531;
    wire N__35524;
    wire N__35523;
    wire N__35522;
    wire N__35515;
    wire N__35514;
    wire N__35513;
    wire N__35506;
    wire N__35505;
    wire N__35504;
    wire N__35497;
    wire N__35496;
    wire N__35495;
    wire N__35488;
    wire N__35487;
    wire N__35486;
    wire N__35479;
    wire N__35478;
    wire N__35477;
    wire N__35470;
    wire N__35469;
    wire N__35468;
    wire N__35461;
    wire N__35460;
    wire N__35459;
    wire N__35442;
    wire N__35439;
    wire N__35438;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35427;
    wire N__35426;
    wire N__35425;
    wire N__35422;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35410;
    wire N__35407;
    wire N__35406;
    wire N__35403;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35383;
    wire N__35380;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35345;
    wire N__35342;
    wire N__35337;
    wire N__35334;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35316;
    wire N__35313;
    wire N__35312;
    wire N__35311;
    wire N__35310;
    wire N__35309;
    wire N__35308;
    wire N__35307;
    wire N__35306;
    wire N__35305;
    wire N__35304;
    wire N__35303;
    wire N__35302;
    wire N__35301;
    wire N__35300;
    wire N__35299;
    wire N__35298;
    wire N__35289;
    wire N__35280;
    wire N__35271;
    wire N__35262;
    wire N__35261;
    wire N__35256;
    wire N__35251;
    wire N__35248;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35226;
    wire N__35223;
    wire N__35222;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35201;
    wire N__35200;
    wire N__35197;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35180;
    wire N__35175;
    wire N__35172;
    wire N__35169;
    wire N__35168;
    wire N__35165;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35148;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35132;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35108;
    wire N__35105;
    wire N__35102;
    wire N__35097;
    wire N__35096;
    wire N__35095;
    wire N__35094;
    wire N__35093;
    wire N__35092;
    wire N__35091;
    wire N__35090;
    wire N__35089;
    wire N__35088;
    wire N__35087;
    wire N__35086;
    wire N__35085;
    wire N__35084;
    wire N__35083;
    wire N__35082;
    wire N__35081;
    wire N__35080;
    wire N__35079;
    wire N__35078;
    wire N__35077;
    wire N__35076;
    wire N__35075;
    wire N__35074;
    wire N__35073;
    wire N__35072;
    wire N__35071;
    wire N__35070;
    wire N__35065;
    wire N__35058;
    wire N__35055;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35019;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35001;
    wire N__34996;
    wire N__34995;
    wire N__34994;
    wire N__34993;
    wire N__34992;
    wire N__34991;
    wire N__34990;
    wire N__34989;
    wire N__34988;
    wire N__34987;
    wire N__34986;
    wire N__34985;
    wire N__34984;
    wire N__34983;
    wire N__34982;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34850;
    wire N__34849;
    wire N__34848;
    wire N__34845;
    wire N__34838;
    wire N__34837;
    wire N__34832;
    wire N__34831;
    wire N__34830;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34781;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34746;
    wire N__34743;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34726;
    wire N__34725;
    wire N__34724;
    wire N__34723;
    wire N__34722;
    wire N__34721;
    wire N__34716;
    wire N__34705;
    wire N__34702;
    wire N__34701;
    wire N__34696;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34648;
    wire N__34641;
    wire N__34640;
    wire N__34639;
    wire N__34638;
    wire N__34637;
    wire N__34636;
    wire N__34635;
    wire N__34634;
    wire N__34633;
    wire N__34632;
    wire N__34631;
    wire N__34630;
    wire N__34629;
    wire N__34628;
    wire N__34627;
    wire N__34626;
    wire N__34625;
    wire N__34624;
    wire N__34623;
    wire N__34622;
    wire N__34621;
    wire N__34620;
    wire N__34619;
    wire N__34618;
    wire N__34617;
    wire N__34616;
    wire N__34615;
    wire N__34614;
    wire N__34613;
    wire N__34612;
    wire N__34611;
    wire N__34610;
    wire N__34609;
    wire N__34608;
    wire N__34607;
    wire N__34606;
    wire N__34605;
    wire N__34604;
    wire N__34603;
    wire N__34602;
    wire N__34601;
    wire N__34600;
    wire N__34599;
    wire N__34598;
    wire N__34597;
    wire N__34596;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34592;
    wire N__34591;
    wire N__34590;
    wire N__34589;
    wire N__34588;
    wire N__34587;
    wire N__34586;
    wire N__34585;
    wire N__34584;
    wire N__34583;
    wire N__34582;
    wire N__34581;
    wire N__34580;
    wire N__34579;
    wire N__34578;
    wire N__34577;
    wire N__34576;
    wire N__34575;
    wire N__34574;
    wire N__34573;
    wire N__34572;
    wire N__34571;
    wire N__34570;
    wire N__34569;
    wire N__34568;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34564;
    wire N__34563;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34557;
    wire N__34556;
    wire N__34555;
    wire N__34554;
    wire N__34553;
    wire N__34552;
    wire N__34551;
    wire N__34550;
    wire N__34549;
    wire N__34548;
    wire N__34547;
    wire N__34546;
    wire N__34545;
    wire N__34544;
    wire N__34543;
    wire N__34542;
    wire N__34541;
    wire N__34540;
    wire N__34539;
    wire N__34538;
    wire N__34537;
    wire N__34536;
    wire N__34535;
    wire N__34534;
    wire N__34533;
    wire N__34532;
    wire N__34531;
    wire N__34530;
    wire N__34529;
    wire N__34528;
    wire N__34527;
    wire N__34526;
    wire N__34525;
    wire N__34524;
    wire N__34523;
    wire N__34522;
    wire N__34521;
    wire N__34520;
    wire N__34519;
    wire N__34518;
    wire N__34517;
    wire N__34516;
    wire N__34515;
    wire N__34514;
    wire N__34257;
    wire N__34254;
    wire N__34251;
    wire N__34248;
    wire N__34245;
    wire N__34242;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34211;
    wire N__34208;
    wire N__34205;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34193;
    wire N__34192;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34174;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34159;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34097;
    wire N__34094;
    wire N__34091;
    wire N__34088;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34046;
    wire N__34043;
    wire N__34042;
    wire N__34041;
    wire N__34038;
    wire N__34037;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34020;
    wire N__34017;
    wire N__34016;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33980;
    wire N__33979;
    wire N__33974;
    wire N__33971;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33955;
    wire N__33952;
    wire N__33947;
    wire N__33944;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33912;
    wire N__33909;
    wire N__33908;
    wire N__33905;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33897;
    wire N__33896;
    wire N__33893;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33865;
    wire N__33862;
    wire N__33859;
    wire N__33854;
    wire N__33851;
    wire N__33846;
    wire N__33845;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33796;
    wire N__33793;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33761;
    wire N__33756;
    wire N__33753;
    wire N__33750;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33732;
    wire N__33731;
    wire N__33730;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33705;
    wire N__33702;
    wire N__33701;
    wire N__33698;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33662;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33612;
    wire N__33609;
    wire N__33608;
    wire N__33607;
    wire N__33606;
    wire N__33605;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33585;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33502;
    wire N__33499;
    wire N__33492;
    wire N__33489;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33471;
    wire N__33468;
    wire N__33467;
    wire N__33464;
    wire N__33463;
    wire N__33460;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33416;
    wire N__33413;
    wire N__33406;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33348;
    wire N__33345;
    wire N__33344;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33312;
    wire N__33309;
    wire N__33306;
    wire N__33305;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33270;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33246;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33129;
    wire N__33126;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33071;
    wire N__33068;
    wire N__33067;
    wire N__33066;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33047;
    wire N__33042;
    wire N__33041;
    wire N__33038;
    wire N__33035;
    wire N__33034;
    wire N__33031;
    wire N__33030;
    wire N__33029;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33004;
    wire N__32997;
    wire N__32996;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32967;
    wire N__32966;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32950;
    wire N__32949;
    wire N__32944;
    wire N__32943;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32924;
    wire N__32917;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32894;
    wire N__32893;
    wire N__32892;
    wire N__32887;
    wire N__32882;
    wire N__32881;
    wire N__32880;
    wire N__32879;
    wire N__32878;
    wire N__32877;
    wire N__32876;
    wire N__32871;
    wire N__32866;
    wire N__32865;
    wire N__32864;
    wire N__32863;
    wire N__32862;
    wire N__32861;
    wire N__32860;
    wire N__32859;
    wire N__32858;
    wire N__32857;
    wire N__32856;
    wire N__32855;
    wire N__32854;
    wire N__32853;
    wire N__32852;
    wire N__32851;
    wire N__32850;
    wire N__32849;
    wire N__32848;
    wire N__32847;
    wire N__32846;
    wire N__32845;
    wire N__32844;
    wire N__32843;
    wire N__32842;
    wire N__32837;
    wire N__32832;
    wire N__32827;
    wire N__32820;
    wire N__32817;
    wire N__32808;
    wire N__32803;
    wire N__32798;
    wire N__32789;
    wire N__32780;
    wire N__32779;
    wire N__32778;
    wire N__32775;
    wire N__32774;
    wire N__32773;
    wire N__32770;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32754;
    wire N__32747;
    wire N__32744;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32721;
    wire N__32710;
    wire N__32707;
    wire N__32694;
    wire N__32693;
    wire N__32692;
    wire N__32691;
    wire N__32690;
    wire N__32689;
    wire N__32688;
    wire N__32687;
    wire N__32686;
    wire N__32685;
    wire N__32684;
    wire N__32683;
    wire N__32682;
    wire N__32681;
    wire N__32680;
    wire N__32679;
    wire N__32678;
    wire N__32677;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32669;
    wire N__32668;
    wire N__32667;
    wire N__32666;
    wire N__32665;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32657;
    wire N__32656;
    wire N__32655;
    wire N__32654;
    wire N__32653;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32641;
    wire N__32638;
    wire N__32633;
    wire N__32628;
    wire N__32623;
    wire N__32618;
    wire N__32613;
    wire N__32606;
    wire N__32601;
    wire N__32598;
    wire N__32591;
    wire N__32588;
    wire N__32587;
    wire N__32586;
    wire N__32583;
    wire N__32582;
    wire N__32575;
    wire N__32574;
    wire N__32573;
    wire N__32572;
    wire N__32571;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32557;
    wire N__32538;
    wire N__32533;
    wire N__32524;
    wire N__32521;
    wire N__32516;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32502;
    wire N__32495;
    wire N__32490;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32462;
    wire N__32461;
    wire N__32460;
    wire N__32459;
    wire N__32458;
    wire N__32457;
    wire N__32456;
    wire N__32455;
    wire N__32454;
    wire N__32453;
    wire N__32444;
    wire N__32443;
    wire N__32442;
    wire N__32441;
    wire N__32440;
    wire N__32439;
    wire N__32438;
    wire N__32437;
    wire N__32436;
    wire N__32435;
    wire N__32434;
    wire N__32433;
    wire N__32432;
    wire N__32431;
    wire N__32430;
    wire N__32429;
    wire N__32428;
    wire N__32427;
    wire N__32426;
    wire N__32421;
    wire N__32414;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32394;
    wire N__32385;
    wire N__32384;
    wire N__32383;
    wire N__32378;
    wire N__32377;
    wire N__32376;
    wire N__32375;
    wire N__32374;
    wire N__32373;
    wire N__32368;
    wire N__32359;
    wire N__32356;
    wire N__32349;
    wire N__32340;
    wire N__32337;
    wire N__32336;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32323;
    wire N__32320;
    wire N__32315;
    wire N__32310;
    wire N__32303;
    wire N__32296;
    wire N__32287;
    wire N__32280;
    wire N__32277;
    wire N__32270;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32178;
    wire N__32175;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32010;
    wire N__32009;
    wire N__32006;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31991;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31959;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31925;
    wire N__31922;
    wire N__31919;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31874;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31858;
    wire N__31853;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31825;
    wire N__31820;
    wire N__31817;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31790;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31774;
    wire N__31771;
    wire N__31766;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31682;
    wire N__31679;
    wire N__31678;
    wire N__31677;
    wire N__31674;
    wire N__31673;
    wire N__31672;
    wire N__31671;
    wire N__31668;
    wire N__31667;
    wire N__31664;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31653;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31582;
    wire N__31579;
    wire N__31578;
    wire N__31571;
    wire N__31566;
    wire N__31563;
    wire N__31556;
    wire N__31553;
    wire N__31552;
    wire N__31549;
    wire N__31546;
    wire N__31543;
    wire N__31536;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31520;
    wire N__31517;
    wire N__31512;
    wire N__31503;
    wire N__31502;
    wire N__31501;
    wire N__31500;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31482;
    wire N__31481;
    wire N__31480;
    wire N__31479;
    wire N__31478;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31457;
    wire N__31454;
    wire N__31453;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31441;
    wire N__31438;
    wire N__31437;
    wire N__31434;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31418;
    wire N__31415;
    wire N__31412;
    wire N__31407;
    wire N__31404;
    wire N__31399;
    wire N__31396;
    wire N__31393;
    wire N__31388;
    wire N__31383;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31356;
    wire N__31353;
    wire N__31346;
    wire N__31335;
    wire N__31334;
    wire N__31331;
    wire N__31330;
    wire N__31329;
    wire N__31326;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31315;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31262;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31248;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31227;
    wire N__31224;
    wire N__31219;
    wire N__31216;
    wire N__31213;
    wire N__31210;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31190;
    wire N__31187;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31156;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31133;
    wire N__31130;
    wire N__31125;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31109;
    wire N__31106;
    wire N__31101;
    wire N__31098;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31067;
    wire N__31064;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31050;
    wire N__31047;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31026;
    wire N__31025;
    wire N__31022;
    wire N__31021;
    wire N__31018;
    wire N__31013;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31002;
    wire N__30999;
    wire N__30994;
    wire N__30991;
    wire N__30988;
    wire N__30985;
    wire N__30978;
    wire N__30975;
    wire N__30974;
    wire N__30971;
    wire N__30970;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30945;
    wire N__30944;
    wire N__30943;
    wire N__30942;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30930;
    wire N__30927;
    wire N__30922;
    wire N__30919;
    wire N__30918;
    wire N__30915;
    wire N__30910;
    wire N__30907;
    wire N__30902;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30842;
    wire N__30841;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30824;
    wire N__30823;
    wire N__30822;
    wire N__30821;
    wire N__30818;
    wire N__30813;
    wire N__30812;
    wire N__30809;
    wire N__30802;
    wire N__30799;
    wire N__30794;
    wire N__30791;
    wire N__30780;
    wire N__30779;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30766;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30715;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30695;
    wire N__30694;
    wire N__30691;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30676;
    wire N__30671;
    wire N__30668;
    wire N__30663;
    wire N__30660;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30635;
    wire N__30634;
    wire N__30633;
    wire N__30632;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30624;
    wire N__30617;
    wire N__30614;
    wire N__30609;
    wire N__30606;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30590;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30566;
    wire N__30563;
    wire N__30560;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30515;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30494;
    wire N__30493;
    wire N__30490;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30475;
    wire N__30474;
    wire N__30471;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30453;
    wire N__30452;
    wire N__30449;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30428;
    wire N__30427;
    wire N__30426;
    wire N__30425;
    wire N__30420;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30395;
    wire N__30394;
    wire N__30391;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30367;
    wire N__30364;
    wire N__30355;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30334;
    wire N__30331;
    wire N__30324;
    wire N__30321;
    wire N__30320;
    wire N__30319;
    wire N__30318;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30303;
    wire N__30296;
    wire N__30295;
    wire N__30294;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30280;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30243;
    wire N__30242;
    wire N__30241;
    wire N__30240;
    wire N__30239;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30221;
    wire N__30220;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30198;
    wire N__30197;
    wire N__30194;
    wire N__30189;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30162;
    wire N__30161;
    wire N__30160;
    wire N__30159;
    wire N__30158;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30102;
    wire N__30099;
    wire N__30096;
    wire N__30093;
    wire N__30088;
    wire N__30085;
    wire N__30084;
    wire N__30081;
    wire N__30076;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30054;
    wire N__30053;
    wire N__30052;
    wire N__30051;
    wire N__30050;
    wire N__30049;
    wire N__30048;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__29999;
    wire N__29990;
    wire N__29985;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29973;
    wire N__29970;
    wire N__29969;
    wire N__29966;
    wire N__29965;
    wire N__29962;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29951;
    wire N__29950;
    wire N__29949;
    wire N__29948;
    wire N__29947;
    wire N__29944;
    wire N__29939;
    wire N__29936;
    wire N__29931;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29906;
    wire N__29901;
    wire N__29898;
    wire N__29897;
    wire N__29896;
    wire N__29895;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29866;
    wire N__29863;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29837;
    wire N__29836;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29826;
    wire N__29821;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29804;
    wire N__29801;
    wire N__29796;
    wire N__29793;
    wire N__29792;
    wire N__29789;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29773;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29743;
    wire N__29742;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29727;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29707;
    wire N__29704;
    wire N__29699;
    wire N__29694;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29657;
    wire N__29656;
    wire N__29653;
    wire N__29652;
    wire N__29651;
    wire N__29650;
    wire N__29649;
    wire N__29648;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29633;
    wire N__29632;
    wire N__29631;
    wire N__29630;
    wire N__29629;
    wire N__29628;
    wire N__29627;
    wire N__29624;
    wire N__29623;
    wire N__29618;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29584;
    wire N__29581;
    wire N__29574;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29543;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29522;
    wire N__29521;
    wire N__29520;
    wire N__29519;
    wire N__29516;
    wire N__29511;
    wire N__29508;
    wire N__29507;
    wire N__29504;
    wire N__29503;
    wire N__29500;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29492;
    wire N__29491;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29419;
    wire N__29414;
    wire N__29409;
    wire N__29406;
    wire N__29401;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29380;
    wire N__29373;
    wire N__29370;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29343;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29324;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29316;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29299;
    wire N__29298;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29277;
    wire N__29274;
    wire N__29273;
    wire N__29272;
    wire N__29269;
    wire N__29268;
    wire N__29265;
    wire N__29258;
    wire N__29255;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29237;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29229;
    wire N__29224;
    wire N__29221;
    wire N__29216;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29191;
    wire N__29188;
    wire N__29185;
    wire N__29180;
    wire N__29173;
    wire N__29170;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29146;
    wire N__29141;
    wire N__29138;
    wire N__29127;
    wire N__29126;
    wire N__29125;
    wire N__29122;
    wire N__29117;
    wire N__29116;
    wire N__29115;
    wire N__29114;
    wire N__29113;
    wire N__29112;
    wire N__29111;
    wire N__29106;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29092;
    wire N__29091;
    wire N__29088;
    wire N__29087;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29057;
    wire N__29054;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29021;
    wire N__29020;
    wire N__29019;
    wire N__29018;
    wire N__29017;
    wire N__29016;
    wire N__29013;
    wire N__29012;
    wire N__29011;
    wire N__29010;
    wire N__29009;
    wire N__29008;
    wire N__29007;
    wire N__29004;
    wire N__29003;
    wire N__29000;
    wire N__28999;
    wire N__28996;
    wire N__28995;
    wire N__28994;
    wire N__28993;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28973;
    wire N__28968;
    wire N__28963;
    wire N__28956;
    wire N__28951;
    wire N__28948;
    wire N__28947;
    wire N__28946;
    wire N__28943;
    wire N__28942;
    wire N__28941;
    wire N__28938;
    wire N__28933;
    wire N__28928;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28914;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28881;
    wire N__28878;
    wire N__28869;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28861;
    wire N__28860;
    wire N__28859;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28838;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28824;
    wire N__28821;
    wire N__28820;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28806;
    wire N__28805;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28765;
    wire N__28764;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28730;
    wire N__28727;
    wire N__28722;
    wire N__28715;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28668;
    wire N__28667;
    wire N__28666;
    wire N__28665;
    wire N__28664;
    wire N__28663;
    wire N__28662;
    wire N__28661;
    wire N__28660;
    wire N__28659;
    wire N__28658;
    wire N__28657;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28604;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28593;
    wire N__28592;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28578;
    wire N__28575;
    wire N__28574;
    wire N__28571;
    wire N__28570;
    wire N__28565;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28555;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28540;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28504;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28458;
    wire N__28453;
    wire N__28450;
    wire N__28445;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28426;
    wire N__28421;
    wire N__28418;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28328;
    wire N__28327;
    wire N__28326;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28217;
    wire N__28214;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28187;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28100;
    wire N__28099;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28091;
    wire N__28090;
    wire N__28087;
    wire N__28086;
    wire N__28085;
    wire N__28084;
    wire N__28083;
    wire N__28080;
    wire N__28079;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28065;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27968;
    wire N__27963;
    wire N__27956;
    wire N__27953;
    wire N__27946;
    wire N__27943;
    wire N__27938;
    wire N__27929;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27890;
    wire N__27889;
    wire N__27888;
    wire N__27887;
    wire N__27886;
    wire N__27885;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27877;
    wire N__27876;
    wire N__27873;
    wire N__27872;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27833;
    wire N__27832;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27776;
    wire N__27771;
    wire N__27770;
    wire N__27767;
    wire N__27766;
    wire N__27757;
    wire N__27754;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27740;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27721;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27700;
    wire N__27693;
    wire N__27684;
    wire N__27683;
    wire N__27682;
    wire N__27681;
    wire N__27680;
    wire N__27679;
    wire N__27678;
    wire N__27677;
    wire N__27676;
    wire N__27673;
    wire N__27670;
    wire N__27669;
    wire N__27668;
    wire N__27667;
    wire N__27666;
    wire N__27663;
    wire N__27658;
    wire N__27653;
    wire N__27648;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27636;
    wire N__27633;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27625;
    wire N__27622;
    wire N__27611;
    wire N__27608;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27585;
    wire N__27584;
    wire N__27581;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27555;
    wire N__27554;
    wire N__27553;
    wire N__27552;
    wire N__27551;
    wire N__27550;
    wire N__27549;
    wire N__27548;
    wire N__27547;
    wire N__27546;
    wire N__27545;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27539;
    wire N__27538;
    wire N__27537;
    wire N__27536;
    wire N__27533;
    wire N__27528;
    wire N__27527;
    wire N__27522;
    wire N__27521;
    wire N__27520;
    wire N__27519;
    wire N__27518;
    wire N__27515;
    wire N__27514;
    wire N__27511;
    wire N__27506;
    wire N__27505;
    wire N__27504;
    wire N__27503;
    wire N__27498;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27478;
    wire N__27475;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27461;
    wire N__27460;
    wire N__27459;
    wire N__27458;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27443;
    wire N__27440;
    wire N__27435;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27419;
    wire N__27418;
    wire N__27417;
    wire N__27416;
    wire N__27409;
    wire N__27406;
    wire N__27401;
    wire N__27394;
    wire N__27391;
    wire N__27378;
    wire N__27371;
    wire N__27362;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27333;
    wire N__27330;
    wire N__27329;
    wire N__27328;
    wire N__27327;
    wire N__27324;
    wire N__27319;
    wire N__27316;
    wire N__27309;
    wire N__27306;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27298;
    wire N__27297;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27283;
    wire N__27276;
    wire N__27275;
    wire N__27274;
    wire N__27273;
    wire N__27270;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27252;
    wire N__27251;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27203;
    wire N__27200;
    wire N__27193;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27172;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27161;
    wire N__27160;
    wire N__27159;
    wire N__27156;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27137;
    wire N__27134;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27098;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27062;
    wire N__27061;
    wire N__27058;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27046;
    wire N__27043;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26968;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26822;
    wire N__26821;
    wire N__26820;
    wire N__26817;
    wire N__26816;
    wire N__26815;
    wire N__26812;
    wire N__26811;
    wire N__26810;
    wire N__26809;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26801;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26750;
    wire N__26749;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26698;
    wire N__26695;
    wire N__26690;
    wire N__26683;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26662;
    wire N__26655;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26633;
    wire N__26630;
    wire N__26623;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26556;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26498;
    wire N__26497;
    wire N__26496;
    wire N__26493;
    wire N__26492;
    wire N__26491;
    wire N__26484;
    wire N__26483;
    wire N__26480;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26458;
    wire N__26455;
    wire N__26450;
    wire N__26445;
    wire N__26442;
    wire N__26441;
    wire N__26438;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26411;
    wire N__26408;
    wire N__26407;
    wire N__26406;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26389;
    wire N__26382;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26309;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26298;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26286;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26259;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26230;
    wire N__26229;
    wire N__26228;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26183;
    wire N__26182;
    wire N__26181;
    wire N__26180;
    wire N__26179;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26150;
    wire N__26147;
    wire N__26144;
    wire N__26143;
    wire N__26142;
    wire N__26141;
    wire N__26134;
    wire N__26129;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26062;
    wire N__26055;
    wire N__26052;
    wire N__26051;
    wire N__26050;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26021;
    wire N__26020;
    wire N__26019;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26008;
    wire N__26007;
    wire N__26006;
    wire N__26005;
    wire N__26004;
    wire N__26001;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25984;
    wire N__25983;
    wire N__25982;
    wire N__25981;
    wire N__25978;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25914;
    wire N__25911;
    wire N__25902;
    wire N__25899;
    wire N__25896;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25884;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25863;
    wire N__25858;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25840;
    wire N__25837;
    wire N__25832;
    wire N__25829;
    wire N__25828;
    wire N__25823;
    wire N__25816;
    wire N__25813;
    wire N__25808;
    wire N__25805;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25784;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25776;
    wire N__25773;
    wire N__25772;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25751;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25726;
    wire N__25725;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25713;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25694;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25682;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25620;
    wire N__25613;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25595;
    wire N__25590;
    wire N__25589;
    wire N__25588;
    wire N__25585;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25577;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25547;
    wire N__25546;
    wire N__25545;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25531;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25512;
    wire N__25511;
    wire N__25508;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25471;
    wire N__25468;
    wire N__25463;
    wire N__25460;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25429;
    wire N__25424;
    wire N__25415;
    wire N__25412;
    wire N__25411;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25370;
    wire N__25367;
    wire N__25366;
    wire N__25363;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25349;
    wire N__25348;
    wire N__25343;
    wire N__25342;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25303;
    wire N__25300;
    wire N__25295;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25260;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25247;
    wire N__25246;
    wire N__25245;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25234;
    wire N__25233;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25225;
    wire N__25222;
    wire N__25217;
    wire N__25210;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25194;
    wire N__25191;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25172;
    wire N__25171;
    wire N__25170;
    wire N__25169;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25158;
    wire N__25157;
    wire N__25156;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25130;
    wire N__25129;
    wire N__25128;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25114;
    wire N__25113;
    wire N__25110;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25022;
    wire N__25019;
    wire N__25018;
    wire N__25013;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24978;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24960;
    wire N__24955;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24834;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24707;
    wire N__24706;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24691;
    wire N__24690;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24679;
    wire N__24678;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24643;
    wire N__24642;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24607;
    wire N__24604;
    wire N__24603;
    wire N__24596;
    wire N__24593;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24562;
    wire N__24557;
    wire N__24554;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24533;
    wire N__24526;
    wire N__24525;
    wire N__24524;
    wire N__24521;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24494;
    wire N__24491;
    wire N__24490;
    wire N__24489;
    wire N__24486;
    wire N__24485;
    wire N__24484;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24465;
    wire N__24462;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24438;
    wire N__24437;
    wire N__24434;
    wire N__24433;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24422;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24404;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24365;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24357;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24343;
    wire N__24340;
    wire N__24339;
    wire N__24338;
    wire N__24337;
    wire N__24334;
    wire N__24333;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24319;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24307;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24297;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24242;
    wire N__24237;
    wire N__24234;
    wire N__24227;
    wire N__24224;
    wire N__24219;
    wire N__24216;
    wire N__24215;
    wire N__24210;
    wire N__24207;
    wire N__24198;
    wire N__24195;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24181;
    wire N__24178;
    wire N__24173;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23987;
    wire N__23986;
    wire N__23985;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23977;
    wire N__23976;
    wire N__23973;
    wire N__23972;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23964;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23925;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23855;
    wire N__23852;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23832;
    wire N__23825;
    wire N__23824;
    wire N__23819;
    wire N__23816;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23801;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23775;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23699;
    wire N__23698;
    wire N__23697;
    wire N__23696;
    wire N__23695;
    wire N__23692;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23670;
    wire N__23663;
    wire N__23660;
    wire N__23653;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23639;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23624;
    wire N__23621;
    wire N__23620;
    wire N__23619;
    wire N__23618;
    wire N__23617;
    wire N__23612;
    wire N__23609;
    wire N__23608;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23583;
    wire N__23582;
    wire N__23581;
    wire N__23580;
    wire N__23571;
    wire N__23568;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23553;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23538;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23523;
    wire N__23520;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23505;
    wire N__23502;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23487;
    wire N__23484;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23469;
    wire N__23466;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23451;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23433;
    wire N__23432;
    wire N__23431;
    wire N__23430;
    wire N__23429;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23360;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23345;
    wire N__23344;
    wire N__23343;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23316;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23304;
    wire N__23301;
    wire N__23294;
    wire N__23289;
    wire N__23286;
    wire N__23285;
    wire N__23284;
    wire N__23283;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23246;
    wire N__23245;
    wire N__23244;
    wire N__23241;
    wire N__23234;
    wire N__23229;
    wire N__23226;
    wire N__23223;
    wire N__23222;
    wire N__23221;
    wire N__23218;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23203;
    wire N__23202;
    wire N__23197;
    wire N__23194;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23175;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23144;
    wire N__23141;
    wire N__23140;
    wire N__23139;
    wire N__23138;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23099;
    wire N__23096;
    wire N__23095;
    wire N__23092;
    wire N__23091;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23077;
    wire N__23074;
    wire N__23073;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23044;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23005;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22993;
    wire N__22992;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22949;
    wire N__22938;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22930;
    wire N__22929;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22902;
    wire N__22893;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22882;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22870;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22817;
    wire N__22814;
    wire N__22813;
    wire N__22812;
    wire N__22811;
    wire N__22808;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22765;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22628;
    wire N__22625;
    wire N__22624;
    wire N__22621;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22535;
    wire N__22532;
    wire N__22531;
    wire N__22530;
    wire N__22529;
    wire N__22528;
    wire N__22527;
    wire N__22526;
    wire N__22525;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22511;
    wire N__22508;
    wire N__22507;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22364;
    wire N__22359;
    wire N__22354;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22333;
    wire N__22328;
    wire N__22323;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22269;
    wire N__22266;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22124;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22068;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22038;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22023;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22008;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21993;
    wire N__21992;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21934;
    wire N__21933;
    wire N__21932;
    wire N__21929;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21893;
    wire N__21892;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21845;
    wire N__21844;
    wire N__21843;
    wire N__21842;
    wire N__21839;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21802;
    wire N__21801;
    wire N__21798;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21758;
    wire N__21757;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21732;
    wire N__21731;
    wire N__21730;
    wire N__21729;
    wire N__21728;
    wire N__21723;
    wire N__21722;
    wire N__21721;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21703;
    wire N__21700;
    wire N__21687;
    wire N__21686;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21674;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21663;
    wire N__21662;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21648;
    wire N__21645;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21629;
    wire N__21628;
    wire N__21627;
    wire N__21624;
    wire N__21617;
    wire N__21616;
    wire N__21611;
    wire N__21608;
    wire N__21603;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21592;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21580;
    wire N__21577;
    wire N__21576;
    wire N__21575;
    wire N__21572;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21552;
    wire N__21551;
    wire N__21550;
    wire N__21549;
    wire N__21548;
    wire N__21543;
    wire N__21538;
    wire N__21535;
    wire N__21534;
    wire N__21533;
    wire N__21528;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21502;
    wire N__21495;
    wire N__21492;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21484;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21476;
    wire N__21471;
    wire N__21470;
    wire N__21469;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21453;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21404;
    wire N__21401;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21345;
    wire N__21342;
    wire N__21333;
    wire N__21332;
    wire N__21329;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21312;
    wire N__21309;
    wire N__21308;
    wire N__21305;
    wire N__21302;
    wire N__21301;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21285;
    wire N__21282;
    wire N__21281;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21258;
    wire N__21257;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21114;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21079;
    wire N__21078;
    wire N__21077;
    wire N__21074;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21024;
    wire N__21021;
    wire N__21020;
    wire N__21017;
    wire N__21016;
    wire N__21013;
    wire N__21012;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20995;
    wire N__20990;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20978;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20960;
    wire N__20957;
    wire N__20952;
    wire N__20947;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20900;
    wire N__20899;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20875;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20846;
    wire N__20843;
    wire N__20842;
    wire N__20839;
    wire N__20838;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20811;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20799;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20723;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20715;
    wire N__20712;
    wire N__20707;
    wire N__20704;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20618;
    wire N__20615;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20598;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20575;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20529;
    wire N__20528;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20501;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20454;
    wire N__20453;
    wire N__20450;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20370;
    wire N__20367;
    wire N__20366;
    wire N__20363;
    wire N__20362;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20350;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20324;
    wire N__20323;
    wire N__20320;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20282;
    wire N__20281;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20232;
    wire N__20231;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20216;
    wire N__20213;
    wire N__20206;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20147;
    wire N__20144;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20114;
    wire N__20113;
    wire N__20110;
    wire N__20105;
    wire N__20100;
    wire N__20099;
    wire N__20098;
    wire N__20097;
    wire N__20096;
    wire N__20093;
    wire N__20092;
    wire N__20091;
    wire N__20088;
    wire N__20087;
    wire N__20086;
    wire N__20085;
    wire N__20084;
    wire N__20083;
    wire N__20082;
    wire N__20081;
    wire N__20080;
    wire N__20077;
    wire N__20076;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20068;
    wire N__20067;
    wire N__20064;
    wire N__20061;
    wire N__20058;
    wire N__20057;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20046;
    wire N__20043;
    wire N__20042;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20034;
    wire N__20031;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20013;
    wire N__20012;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19987;
    wire N__19986;
    wire N__19979;
    wire N__19976;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19968;
    wire N__19965;
    wire N__19964;
    wire N__19957;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19924;
    wire N__19917;
    wire N__19914;
    wire N__19913;
    wire N__19912;
    wire N__19911;
    wire N__19910;
    wire N__19907;
    wire N__19902;
    wire N__19899;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19887;
    wire N__19884;
    wire N__19879;
    wire N__19878;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19866;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19854;
    wire N__19851;
    wire N__19850;
    wire N__19849;
    wire N__19846;
    wire N__19845;
    wire N__19842;
    wire N__19841;
    wire N__19838;
    wire N__19837;
    wire N__19836;
    wire N__19835;
    wire N__19828;
    wire N__19823;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19802;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19781;
    wire N__19766;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19758;
    wire N__19755;
    wire N__19750;
    wire N__19747;
    wire N__19746;
    wire N__19745;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19733;
    wire N__19730;
    wire N__19729;
    wire N__19724;
    wire N__19721;
    wire N__19714;
    wire N__19711;
    wire N__19706;
    wire N__19695;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19676;
    wire N__19671;
    wire N__19668;
    wire N__19667;
    wire N__19662;
    wire N__19659;
    wire N__19658;
    wire N__19655;
    wire N__19650;
    wire N__19647;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19606;
    wire N__19603;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19585;
    wire N__19582;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19543;
    wire N__19540;
    wire N__19535;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19457;
    wire N__19456;
    wire N__19455;
    wire N__19454;
    wire N__19453;
    wire N__19452;
    wire N__19451;
    wire N__19450;
    wire N__19449;
    wire N__19448;
    wire N__19447;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19428;
    wire N__19417;
    wire N__19414;
    wire N__19401;
    wire N__19398;
    wire N__19397;
    wire N__19396;
    wire N__19395;
    wire N__19394;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19362;
    wire N__19361;
    wire N__19360;
    wire N__19357;
    wire N__19352;
    wire N__19347;
    wire N__19344;
    wire N__19343;
    wire N__19342;
    wire N__19339;
    wire N__19334;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19316;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19271;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19184;
    wire N__19183;
    wire N__19180;
    wire N__19175;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19163;
    wire N__19158;
    wire N__19155;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19139;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19077;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19046;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19023;
    wire N__19020;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire N__18996;
    wire N__18995;
    wire N__18994;
    wire N__18993;
    wire N__18992;
    wire N__18989;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18969;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18954;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18941;
    wire N__18938;
    wire N__18937;
    wire N__18934;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18922;
    wire N__18919;
    wire N__18912;
    wire N__18909;
    wire N__18908;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18854;
    wire N__18853;
    wire N__18852;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18844;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18833;
    wire N__18832;
    wire N__18831;
    wire N__18830;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18790;
    wire N__18789;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18697;
    wire N__18692;
    wire N__18689;
    wire N__18682;
    wire N__18679;
    wire N__18674;
    wire N__18671;
    wire N__18666;
    wire N__18663;
    wire N__18658;
    wire N__18653;
    wire N__18648;
    wire N__18647;
    wire N__18644;
    wire N__18643;
    wire N__18642;
    wire N__18641;
    wire N__18640;
    wire N__18637;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18613;
    wire N__18612;
    wire N__18611;
    wire N__18610;
    wire N__18609;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18597;
    wire N__18596;
    wire N__18591;
    wire N__18590;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18541;
    wire N__18536;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18514;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18492;
    wire N__18489;
    wire N__18486;
    wire N__18483;
    wire N__18480;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18448;
    wire N__18443;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18426;
    wire N__18423;
    wire N__18420;
    wire N__18419;
    wire N__18414;
    wire N__18411;
    wire N__18410;
    wire N__18407;
    wire N__18406;
    wire N__18405;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18391;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18326;
    wire N__18325;
    wire N__18322;
    wire N__18321;
    wire N__18318;
    wire N__18317;
    wire N__18314;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18282;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18262;
    wire N__18261;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18249;
    wire N__18248;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18184;
    wire N__18181;
    wire N__18180;
    wire N__18177;
    wire N__18172;
    wire N__18167;
    wire N__18162;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18145;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18124;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18085;
    wire N__18082;
    wire N__18079;
    wire N__18076;
    wire N__18075;
    wire N__18070;
    wire N__18067;
    wire N__18064;
    wire N__18063;
    wire N__18058;
    wire N__18055;
    wire N__18052;
    wire N__18051;
    wire N__18050;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18038;
    wire N__18035;
    wire N__18034;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18022;
    wire N__18021;
    wire N__18020;
    wire N__18019;
    wire N__18018;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17955;
    wire N__17952;
    wire N__17947;
    wire N__17942;
    wire N__17939;
    wire N__17928;
    wire N__17925;
    wire N__17920;
    wire N__17917;
    wire N__17912;
    wire N__17907;
    wire N__17906;
    wire N__17901;
    wire N__17898;
    wire N__17895;
    wire N__17892;
    wire N__17889;
    wire N__17886;
    wire N__17883;
    wire N__17880;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17872;
    wire N__17869;
    wire N__17864;
    wire N__17859;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17838;
    wire N__17837;
    wire N__17836;
    wire N__17833;
    wire N__17832;
    wire N__17831;
    wire N__17828;
    wire N__17823;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17815;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17785;
    wire N__17782;
    wire N__17777;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17765;
    wire N__17762;
    wire N__17761;
    wire N__17758;
    wire N__17757;
    wire N__17756;
    wire N__17755;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17737;
    wire N__17734;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17715;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17682;
    wire N__17681;
    wire N__17680;
    wire N__17677;
    wire N__17672;
    wire N__17671;
    wire N__17670;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17658;
    wire N__17655;
    wire N__17652;
    wire N__17649;
    wire N__17646;
    wire N__17645;
    wire N__17642;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17618;
    wire N__17615;
    wire N__17610;
    wire N__17607;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17583;
    wire N__17582;
    wire N__17581;
    wire N__17580;
    wire N__17579;
    wire N__17578;
    wire N__17577;
    wire N__17576;
    wire N__17575;
    wire N__17574;
    wire N__17569;
    wire N__17560;
    wire N__17551;
    wire N__17550;
    wire N__17547;
    wire N__17542;
    wire N__17539;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17517;
    wire N__17514;
    wire N__17511;
    wire N__17508;
    wire N__17505;
    wire N__17502;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17445;
    wire N__17442;
    wire N__17439;
    wire N__17436;
    wire N__17435;
    wire N__17434;
    wire N__17433;
    wire N__17432;
    wire N__17429;
    wire N__17428;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17407;
    wire N__17406;
    wire N__17401;
    wire N__17398;
    wire N__17397;
    wire N__17394;
    wire N__17389;
    wire N__17386;
    wire N__17385;
    wire N__17384;
    wire N__17379;
    wire N__17376;
    wire N__17375;
    wire N__17368;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17349;
    wire N__17346;
    wire N__17341;
    wire N__17336;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17309;
    wire N__17308;
    wire N__17307;
    wire N__17306;
    wire N__17305;
    wire N__17302;
    wire N__17301;
    wire N__17300;
    wire N__17299;
    wire N__17296;
    wire N__17289;
    wire N__17288;
    wire N__17287;
    wire N__17286;
    wire N__17285;
    wire N__17284;
    wire N__17283;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17272;
    wire N__17271;
    wire N__17270;
    wire N__17269;
    wire N__17268;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17253;
    wire N__17248;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17229;
    wire N__17226;
    wire N__17217;
    wire N__17212;
    wire N__17207;
    wire N__17204;
    wire N__17195;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17177;
    wire N__17174;
    wire N__17169;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17147;
    wire N__17146;
    wire N__17143;
    wire N__17138;
    wire N__17133;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17118;
    wire N__17117;
    wire N__17116;
    wire N__17115;
    wire N__17112;
    wire N__17109;
    wire N__17108;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17094;
    wire N__17093;
    wire N__17088;
    wire N__17085;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17071;
    wire N__17068;
    wire N__17067;
    wire N__17062;
    wire N__17057;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__16998;
    wire N__16995;
    wire N__16992;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16980;
    wire N__16977;
    wire N__16974;
    wire N__16971;
    wire N__16968;
    wire N__16965;
    wire N__16962;
    wire N__16959;
    wire N__16956;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16932;
    wire N__16929;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16901;
    wire N__16900;
    wire N__16899;
    wire N__16898;
    wire N__16893;
    wire N__16888;
    wire N__16885;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16869;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16861;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16839;
    wire N__16836;
    wire N__16833;
    wire N__16830;
    wire N__16829;
    wire N__16824;
    wire N__16821;
    wire N__16820;
    wire N__16819;
    wire N__16816;
    wire N__16811;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16797;
    wire N__16794;
    wire N__16791;
    wire N__16790;
    wire N__16785;
    wire N__16782;
    wire N__16781;
    wire N__16780;
    wire N__16779;
    wire N__16778;
    wire N__16777;
    wire N__16776;
    wire N__16775;
    wire N__16772;
    wire N__16771;
    wire N__16770;
    wire N__16769;
    wire N__16768;
    wire N__16763;
    wire N__16762;
    wire N__16761;
    wire N__16760;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16746;
    wire N__16743;
    wire N__16738;
    wire N__16731;
    wire N__16728;
    wire N__16723;
    wire N__16718;
    wire N__16717;
    wire N__16716;
    wire N__16715;
    wire N__16712;
    wire N__16711;
    wire N__16710;
    wire N__16709;
    wire N__16708;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16692;
    wire N__16689;
    wire N__16684;
    wire N__16681;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16665;
    wire N__16660;
    wire N__16655;
    wire N__16642;
    wire N__16629;
    wire N__16628;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16620;
    wire N__16619;
    wire N__16616;
    wire N__16615;
    wire N__16614;
    wire N__16611;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16603;
    wire N__16602;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16573;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16542;
    wire N__16541;
    wire N__16540;
    wire N__16539;
    wire N__16538;
    wire N__16537;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16523;
    wire N__16518;
    wire N__16517;
    wire N__16516;
    wire N__16515;
    wire N__16512;
    wire N__16511;
    wire N__16510;
    wire N__16509;
    wire N__16508;
    wire N__16507;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16487;
    wire N__16486;
    wire N__16483;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16467;
    wire N__16458;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16442;
    wire N__16425;
    wire N__16424;
    wire N__16423;
    wire N__16420;
    wire N__16419;
    wire N__16418;
    wire N__16413;
    wire N__16412;
    wire N__16411;
    wire N__16410;
    wire N__16409;
    wire N__16408;
    wire N__16407;
    wire N__16404;
    wire N__16399;
    wire N__16396;
    wire N__16391;
    wire N__16388;
    wire N__16383;
    wire N__16380;
    wire N__16371;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16355;
    wire N__16350;
    wire N__16347;
    wire N__16346;
    wire N__16343;
    wire N__16342;
    wire N__16341;
    wire N__16338;
    wire N__16337;
    wire N__16336;
    wire N__16335;
    wire N__16332;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16320;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16306;
    wire N__16301;
    wire N__16298;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16278;
    wire N__16275;
    wire N__16274;
    wire N__16273;
    wire N__16272;
    wire N__16271;
    wire N__16270;
    wire N__16269;
    wire N__16268;
    wire N__16267;
    wire N__16266;
    wire N__16263;
    wire N__16258;
    wire N__16255;
    wire N__16250;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16234;
    wire N__16221;
    wire N__16218;
    wire N__16217;
    wire N__16216;
    wire N__16213;
    wire N__16208;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16175;
    wire N__16174;
    wire N__16171;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16156;
    wire N__16155;
    wire N__16152;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16128;
    wire N__16125;
    wire N__16116;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16105;
    wire N__16100;
    wire N__16097;
    wire N__16092;
    wire N__16091;
    wire N__16090;
    wire N__16089;
    wire N__16086;
    wire N__16085;
    wire N__16084;
    wire N__16083;
    wire N__16080;
    wire N__16079;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16071;
    wire N__16068;
    wire N__16063;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16048;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16036;
    wire N__16027;
    wire N__16024;
    wire N__16021;
    wire N__16018;
    wire N__16011;
    wire N__16008;
    wire N__15999;
    wire N__15998;
    wire N__15995;
    wire N__15994;
    wire N__15993;
    wire N__15992;
    wire N__15991;
    wire N__15990;
    wire N__15989;
    wire N__15988;
    wire N__15987;
    wire N__15986;
    wire N__15985;
    wire N__15984;
    wire N__15983;
    wire N__15982;
    wire N__15981;
    wire N__15980;
    wire N__15979;
    wire N__15976;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15942;
    wire N__15941;
    wire N__15936;
    wire N__15931;
    wire N__15926;
    wire N__15915;
    wire N__15910;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15879;
    wire N__15878;
    wire N__15877;
    wire N__15874;
    wire N__15869;
    wire N__15864;
    wire N__15861;
    wire N__15860;
    wire N__15859;
    wire N__15856;
    wire N__15853;
    wire N__15850;
    wire N__15843;
    wire N__15842;
    wire N__15841;
    wire N__15838;
    wire N__15835;
    wire N__15830;
    wire N__15825;
    wire N__15824;
    wire N__15821;
    wire N__15820;
    wire N__15817;
    wire N__15814;
    wire N__15811;
    wire N__15804;
    wire N__15803;
    wire N__15802;
    wire N__15799;
    wire N__15794;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15772;
    wire N__15771;
    wire N__15770;
    wire N__15769;
    wire N__15758;
    wire N__15755;
    wire N__15750;
    wire N__15747;
    wire N__15744;
    wire N__15741;
    wire N__15740;
    wire N__15739;
    wire N__15738;
    wire N__15737;
    wire N__15726;
    wire N__15723;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15645;
    wire N__15644;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15627;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15599;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15582;
    wire N__15579;
    wire N__15578;
    wire N__15573;
    wire N__15570;
    wire N__15567;
    wire N__15566;
    wire N__15565;
    wire N__15562;
    wire N__15557;
    wire N__15552;
    wire N__15549;
    wire N__15548;
    wire N__15547;
    wire N__15544;
    wire N__15539;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15513;
    wire N__15510;
    wire N__15509;
    wire N__15506;
    wire N__15505;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15476;
    wire N__15475;
    wire N__15474;
    wire N__15473;
    wire N__15472;
    wire N__15469;
    wire N__15456;
    wire N__15453;
    wire N__15450;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15420;
    wire N__15417;
    wire N__15414;
    wire N__15411;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15371;
    wire N__15370;
    wire N__15367;
    wire N__15366;
    wire N__15365;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15355;
    wire N__15350;
    wire N__15343;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15327;
    wire N__15326;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15304;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15272;
    wire N__15269;
    wire N__15264;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15252;
    wire N__15249;
    wire N__15246;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15234;
    wire N__15233;
    wire N__15232;
    wire N__15229;
    wire N__15224;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15216;
    wire N__15213;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15186;
    wire N__15183;
    wire N__15182;
    wire N__15179;
    wire N__15178;
    wire N__15177;
    wire N__15174;
    wire N__15171;
    wire N__15166;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15146;
    wire N__15143;
    wire N__15142;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15127;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15110;
    wire N__15107;
    wire N__15106;
    wire N__15105;
    wire N__15104;
    wire N__15101;
    wire N__15100;
    wire N__15099;
    wire N__15096;
    wire N__15093;
    wire N__15088;
    wire N__15085;
    wire N__15080;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15051;
    wire N__15050;
    wire N__15049;
    wire N__15048;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15033;
    wire N__15024;
    wire N__15023;
    wire N__15020;
    wire N__15019;
    wire N__15018;
    wire N__15017;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15009;
    wire N__15008;
    wire N__15005;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14985;
    wire N__14980;
    wire N__14967;
    wire N__14966;
    wire N__14965;
    wire N__14962;
    wire N__14961;
    wire N__14960;
    wire N__14959;
    wire N__14958;
    wire N__14957;
    wire N__14956;
    wire N__14953;
    wire N__14946;
    wire N__14943;
    wire N__14940;
    wire N__14937;
    wire N__14934;
    wire N__14931;
    wire N__14930;
    wire N__14929;
    wire N__14926;
    wire N__14921;
    wire N__14920;
    wire N__14919;
    wire N__14916;
    wire N__14909;
    wire N__14906;
    wire N__14905;
    wire N__14902;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14849;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14829;
    wire N__14826;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14807;
    wire N__14806;
    wire N__14805;
    wire N__14802;
    wire N__14795;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14783;
    wire N__14782;
    wire N__14779;
    wire N__14774;
    wire N__14769;
    wire N__14766;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14747;
    wire N__14746;
    wire N__14745;
    wire N__14744;
    wire N__14741;
    wire N__14736;
    wire N__14733;
    wire N__14732;
    wire N__14729;
    wire N__14724;
    wire N__14721;
    wire N__14718;
    wire N__14709;
    wire N__14708;
    wire N__14707;
    wire N__14704;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14689;
    wire N__14682;
    wire N__14679;
    wire N__14678;
    wire N__14673;
    wire N__14670;
    wire N__14667;
    wire N__14664;
    wire N__14663;
    wire N__14662;
    wire N__14661;
    wire N__14660;
    wire N__14659;
    wire N__14658;
    wire N__14655;
    wire N__14650;
    wire N__14647;
    wire N__14640;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14621;
    wire N__14620;
    wire N__14619;
    wire N__14618;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14599;
    wire N__14594;
    wire N__14591;
    wire N__14580;
    wire N__14579;
    wire N__14578;
    wire N__14573;
    wire N__14572;
    wire N__14571;
    wire N__14570;
    wire N__14569;
    wire N__14568;
    wire N__14565;
    wire N__14562;
    wire N__14555;
    wire N__14550;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14508;
    wire N__14507;
    wire N__14506;
    wire N__14505;
    wire N__14502;
    wire N__14501;
    wire N__14500;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14484;
    wire N__14475;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14465;
    wire N__14464;
    wire N__14463;
    wire N__14462;
    wire N__14461;
    wire N__14460;
    wire N__14459;
    wire N__14456;
    wire N__14451;
    wire N__14450;
    wire N__14449;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14431;
    wire N__14426;
    wire N__14423;
    wire N__14416;
    wire N__14413;
    wire N__14412;
    wire N__14411;
    wire N__14410;
    wire N__14409;
    wire N__14408;
    wire N__14407;
    wire N__14406;
    wire N__14405;
    wire N__14404;
    wire N__14403;
    wire N__14402;
    wire N__14401;
    wire N__14400;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14379;
    wire N__14374;
    wire N__14367;
    wire N__14356;
    wire N__14343;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14313;
    wire N__14310;
    wire N__14309;
    wire N__14306;
    wire N__14303;
    wire N__14298;
    wire N__14297;
    wire N__14296;
    wire N__14295;
    wire N__14294;
    wire N__14293;
    wire N__14290;
    wire N__14289;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14278;
    wire N__14271;
    wire N__14270;
    wire N__14267;
    wire N__14266;
    wire N__14263;
    wire N__14262;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14254;
    wire N__14249;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14238;
    wire N__14237;
    wire N__14234;
    wire N__14229;
    wire N__14226;
    wire N__14221;
    wire N__14220;
    wire N__14219;
    wire N__14218;
    wire N__14217;
    wire N__14216;
    wire N__14215;
    wire N__14212;
    wire N__14211;
    wire N__14210;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14196;
    wire N__14189;
    wire N__14186;
    wire N__14181;
    wire N__14170;
    wire N__14161;
    wire N__14158;
    wire N__14139;
    wire N__14138;
    wire N__14137;
    wire N__14134;
    wire N__14133;
    wire N__14132;
    wire N__14129;
    wire N__14128;
    wire N__14127;
    wire N__14126;
    wire N__14125;
    wire N__14124;
    wire N__14123;
    wire N__14118;
    wire N__14115;
    wire N__14108;
    wire N__14105;
    wire N__14100;
    wire N__14095;
    wire N__14094;
    wire N__14091;
    wire N__14090;
    wire N__14089;
    wire N__14088;
    wire N__14087;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14060;
    wire N__14059;
    wire N__14058;
    wire N__14057;
    wire N__14056;
    wire N__14055;
    wire N__14054;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14031;
    wire N__14026;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__13992;
    wire N__13989;
    wire N__13986;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13950;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13923;
    wire N__13922;
    wire N__13921;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13909;
    wire N__13902;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13890;
    wire N__13887;
    wire N__13886;
    wire N__13885;
    wire N__13884;
    wire N__13881;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13870;
    wire N__13869;
    wire N__13868;
    wire N__13867;
    wire N__13864;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13848;
    wire N__13847;
    wire N__13846;
    wire N__13845;
    wire N__13844;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13832;
    wire N__13825;
    wire N__13816;
    wire N__13813;
    wire N__13800;
    wire N__13799;
    wire N__13798;
    wire N__13797;
    wire N__13796;
    wire N__13795;
    wire N__13794;
    wire N__13793;
    wire N__13792;
    wire N__13791;
    wire N__13788;
    wire N__13787;
    wire N__13786;
    wire N__13785;
    wire N__13784;
    wire N__13783;
    wire N__13778;
    wire N__13769;
    wire N__13768;
    wire N__13767;
    wire N__13758;
    wire N__13753;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13736;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13724;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13710;
    wire N__13705;
    wire N__13702;
    wire N__13697;
    wire N__13694;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13668;
    wire N__13667;
    wire N__13666;
    wire N__13661;
    wire N__13660;
    wire N__13659;
    wire N__13656;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13645;
    wire N__13644;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13632;
    wire N__13631;
    wire N__13630;
    wire N__13629;
    wire N__13628;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13616;
    wire N__13609;
    wire N__13606;
    wire N__13597;
    wire N__13584;
    wire N__13581;
    wire N__13580;
    wire N__13579;
    wire N__13574;
    wire N__13571;
    wire N__13570;
    wire N__13569;
    wire N__13568;
    wire N__13565;
    wire N__13564;
    wire N__13563;
    wire N__13562;
    wire N__13561;
    wire N__13560;
    wire N__13559;
    wire N__13556;
    wire N__13549;
    wire N__13546;
    wire N__13543;
    wire N__13542;
    wire N__13539;
    wire N__13536;
    wire N__13533;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13521;
    wire N__13516;
    wire N__13513;
    wire N__13504;
    wire N__13491;
    wire N__13488;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13473;
    wire N__13472;
    wire N__13471;
    wire N__13470;
    wire N__13467;
    wire N__13462;
    wire N__13459;
    wire N__13452;
    wire N__13451;
    wire N__13450;
    wire N__13449;
    wire N__13446;
    wire N__13445;
    wire N__13444;
    wire N__13443;
    wire N__13442;
    wire N__13441;
    wire N__13438;
    wire N__13437;
    wire N__13436;
    wire N__13435;
    wire N__13432;
    wire N__13429;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13417;
    wire N__13408;
    wire N__13401;
    wire N__13398;
    wire N__13383;
    wire N__13380;
    wire N__13379;
    wire N__13378;
    wire N__13377;
    wire N__13376;
    wire N__13375;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13367;
    wire N__13366;
    wire N__13365;
    wire N__13364;
    wire N__13363;
    wire N__13360;
    wire N__13359;
    wire N__13356;
    wire N__13353;
    wire N__13350;
    wire N__13347;
    wire N__13342;
    wire N__13335;
    wire N__13332;
    wire N__13329;
    wire N__13322;
    wire N__13319;
    wire N__13302;
    wire N__13299;
    wire N__13296;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13269;
    wire N__13266;
    wire N__13263;
    wire N__13260;
    wire N__13257;
    wire N__13254;
    wire N__13251;
    wire N__13248;
    wire N__13247;
    wire N__13242;
    wire N__13239;
    wire N__13236;
    wire N__13233;
    wire N__13230;
    wire N__13227;
    wire N__13224;
    wire N__13221;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13206;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13178;
    wire N__13173;
    wire N__13170;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13152;
    wire N__13151;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13138;
    wire N__13131;
    wire N__13130;
    wire N__13127;
    wire N__13126;
    wire N__13123;
    wire N__13120;
    wire N__13115;
    wire N__13110;
    wire N__13107;
    wire N__13106;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13088;
    wire N__13087;
    wire N__13086;
    wire N__13083;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13052;
    wire N__13051;
    wire N__13050;
    wire N__13049;
    wire N__13046;
    wire N__13045;
    wire N__13042;
    wire N__13041;
    wire N__13038;
    wire N__13037;
    wire N__13036;
    wire N__13033;
    wire N__13032;
    wire N__13031;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13008;
    wire N__12999;
    wire N__12984;
    wire N__12981;
    wire N__12980;
    wire N__12979;
    wire N__12976;
    wire N__12975;
    wire N__12974;
    wire N__12973;
    wire N__12970;
    wire N__12969;
    wire N__12968;
    wire N__12967;
    wire N__12966;
    wire N__12965;
    wire N__12962;
    wire N__12959;
    wire N__12956;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12936;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12848;
    wire N__12847;
    wire N__12844;
    wire N__12841;
    wire N__12836;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12785;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12681;
    wire N__12678;
    wire N__12677;
    wire N__12674;
    wire N__12673;
    wire N__12670;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12656;
    wire N__12655;
    wire N__12654;
    wire N__12653;
    wire N__12652;
    wire N__12651;
    wire N__12650;
    wire N__12649;
    wire N__12648;
    wire N__12647;
    wire N__12646;
    wire N__12641;
    wire N__12636;
    wire N__12631;
    wire N__12624;
    wire N__12619;
    wire N__12616;
    wire N__12609;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12573;
    wire N__12570;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12546;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12522;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12507;
    wire N__12504;
    wire N__12503;
    wire N__12502;
    wire N__12501;
    wire N__12500;
    wire N__12497;
    wire N__12490;
    wire N__12487;
    wire N__12480;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12468;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12456;
    wire N__12453;
    wire N__12450;
    wire N__12447;
    wire N__12444;
    wire N__12441;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12419;
    wire N__12418;
    wire N__12415;
    wire N__12410;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12353;
    wire N__12352;
    wire N__12351;
    wire N__12348;
    wire N__12343;
    wire N__12340;
    wire N__12333;
    wire N__12332;
    wire N__12329;
    wire N__12328;
    wire N__12325;
    wire N__12320;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12296;
    wire N__12295;
    wire N__12294;
    wire N__12293;
    wire N__12292;
    wire N__12289;
    wire N__12286;
    wire N__12285;
    wire N__12282;
    wire N__12277;
    wire N__12268;
    wire N__12261;
    wire N__12258;
    wire N__12255;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12243;
    wire N__12240;
    wire N__12239;
    wire N__12238;
    wire N__12237;
    wire N__12236;
    wire N__12235;
    wire N__12234;
    wire N__12233;
    wire N__12230;
    wire N__12221;
    wire N__12218;
    wire N__12213;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire N__12192;
    wire N__12189;
    wire N__12186;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12173;
    wire N__12168;
    wire N__12165;
    wire N__12162;
    wire N__12159;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12149;
    wire N__12148;
    wire N__12147;
    wire N__12146;
    wire N__12145;
    wire N__12142;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12127;
    wire N__12126;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12030;
    wire N__12029;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12014;
    wire N__12013;
    wire N__12012;
    wire N__12011;
    wire N__12010;
    wire N__12005;
    wire N__11996;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11943;
    wire N__11940;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11900;
    wire N__11897;
    wire N__11892;
    wire N__11891;
    wire N__11890;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11870;
    wire N__11867;
    wire N__11864;
    wire N__11863;
    wire N__11858;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11844;
    wire N__11839;
    wire N__11836;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11664;
    wire N__11661;
    wire N__11658;
    wire N__11655;
    wire N__11652;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11624;
    wire N__11623;
    wire N__11620;
    wire N__11619;
    wire N__11616;
    wire N__11609;
    wire N__11606;
    wire N__11605;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11593;
    wire N__11590;
    wire N__11583;
    wire N__11582;
    wire N__11581;
    wire N__11580;
    wire N__11579;
    wire N__11576;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11556;
    wire N__11553;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11426;
    wire N__11425;
    wire N__11418;
    wire N__11415;
    wire N__11414;
    wire N__11413;
    wire N__11410;
    wire N__11405;
    wire N__11400;
    wire N__11399;
    wire N__11398;
    wire N__11397;
    wire N__11396;
    wire N__11395;
    wire N__11392;
    wire N__11385;
    wire N__11380;
    wire N__11375;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11301;
    wire N__11298;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11283;
    wire N__11280;
    wire N__11277;
    wire N__11274;
    wire N__11271;
    wire N__11268;
    wire N__11267;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11214;
    wire N__11211;
    wire N__11208;
    wire N__11205;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11151;
    wire N__11148;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire VCCG0;
    wire GNDG0;
    wire port_data_rw_0_i;
    wire rgb_c_0;
    wire rgb_c_2;
    wire rgb_c_4;
    wire port_nmib_0_i;
    wire rgb_c_3;
    wire this_vga_signals_vvisibility_i;
    wire rgb_c_5;
    wire rgb_c_1;
    wire M_this_map_address_qZ0Z_0;
    wire bfn_7_24_0_;
    wire M_this_map_address_qZ0Z_1;
    wire un1_M_this_map_address_q_cry_0;
    wire M_this_map_address_qZ0Z_2;
    wire un1_M_this_map_address_q_cry_1;
    wire M_this_map_address_qZ0Z_3;
    wire un1_M_this_map_address_q_cry_2;
    wire M_this_map_address_qZ0Z_4;
    wire un1_M_this_map_address_q_cry_3;
    wire M_this_map_address_qZ0Z_5;
    wire un1_M_this_map_address_q_cry_4;
    wire M_this_map_address_qZ0Z_6;
    wire un1_M_this_map_address_q_cry_5;
    wire M_this_map_address_qZ0Z_7;
    wire un1_M_this_map_address_q_cry_6;
    wire un1_M_this_map_address_q_cry_7;
    wire M_this_map_address_qZ0Z_8;
    wire bfn_7_25_0_;
    wire un1_M_this_map_address_q_cry_8;
    wire M_this_map_address_qZ0Z_9;
    wire M_this_vga_signals_address_5;
    wire M_this_vga_signals_address_4;
    wire M_this_vga_signals_address_1;
    wire M_this_vga_signals_address_6;
    wire \this_vga_signals.mult1_un82_sum_c3 ;
    wire \this_vga_signals.N_219 ;
    wire M_this_vram_read_data_2;
    wire M_this_vram_read_data_0;
    wire M_this_vram_read_data_1;
    wire M_this_vram_read_data_3;
    wire \this_vga_signals.g1_1_0_0_0_cascade_ ;
    wire \this_vga_signals.g1_0_1_0_0_cascade_ ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_1_0 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_1 ;
    wire M_this_vga_signals_address_3;
    wire \this_vga_signals.mult1_un61_sum_axb1_cascade_ ;
    wire this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_cascade_;
    wire \this_vga_signals.if_i4_mux ;
    wire \this_vga_signals.if_i4_mux_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_cascade_ ;
    wire \this_vga_signals.g1_0_2 ;
    wire \this_vga_signals.g0_1 ;
    wire \this_vga_signals.g1_4_0 ;
    wire \this_vga_signals.mult1_un61_sum_axb1 ;
    wire \this_vga_signals.g1_7_cascade_ ;
    wire \this_vga_signals.N_6_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_ ;
    wire \this_vga_signals.g1_0_0 ;
    wire \this_vga_signals.N_3_2_0_1 ;
    wire \this_vga_signals.mult1_un61_sum_axb1_3_cascade_ ;
    wire \this_vga_signals.g1_1 ;
    wire \this_vga_signals.g0_0 ;
    wire \this_vga_signals.g0_5_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0_0_0_0 ;
    wire \this_vga_signals.g1_0_0_0 ;
    wire \this_vga_signals.g1_2_1 ;
    wire \this_vga_signals.mult1_un61_sum_axb1_2 ;
    wire \this_vga_ramdac.N_24_mux ;
    wire \this_vga_ramdac.N_2806_reto ;
    wire \this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ;
    wire \this_vga_signals.M_pcounter_q_3_0_cascade_ ;
    wire N_2_0_cascade_;
    wire \this_vga_ramdac.i2_mux_0 ;
    wire \this_vga_ramdac.N_2811_reto ;
    wire \this_vga_ramdac.m16 ;
    wire \this_vga_ramdac.N_2809_reto ;
    wire \this_vga_ramdac.i2_mux ;
    wire \this_vga_ramdac.N_2808_reto ;
    wire \this_vga_ramdac.m6 ;
    wire G_463_cascade_;
    wire \this_vga_ramdac.N_2807_reto ;
    wire N_2_0;
    wire M_this_vga_signals_pixel_clk_0_0;
    wire G_463;
    wire \this_vga_ramdac.m19 ;
    wire \this_vga_ramdac.N_2810_reto ;
    wire M_this_map_ram_write_data_0;
    wire M_this_map_ram_write_data_5;
    wire M_this_map_ram_write_data_6;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_0_cascade_ ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.g1 ;
    wire \this_vga_signals.if_m2_0 ;
    wire \this_vga_signals.if_m2_1 ;
    wire \this_vga_signals.if_m2_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ;
    wire M_this_vga_ramdac_en_0;
    wire M_this_vga_signals_address_2;
    wire \this_vga_signals.g0_i_x4_0_4 ;
    wire this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0;
    wire this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0;
    wire \this_vga_signals.d_N_3_1_i ;
    wire \this_vga_signals.M_hcounter_q_RNIO08E8Z0Z_3 ;
    wire this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3;
    wire \this_vga_signals.g1_0_1_cascade_ ;
    wire \this_vga_signals.g1_2_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_1_0_0_1 ;
    wire \this_vga_signals.mult1_un89_sum_c3_1_0_0_1 ;
    wire this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0;
    wire \this_vga_signals.N_4_2 ;
    wire \this_vga_signals.mult1_un68_sum_axb1 ;
    wire \this_vga_signals.g1_7 ;
    wire \this_vga_signals.g0_i_x4_3_0 ;
    wire \this_vga_signals.mult1_un61_sum_axb1_3_0_cascade_ ;
    wire \this_vga_signals.g1_1_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_1 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_1_cascade_ ;
    wire \this_vga_signals.g1_0_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_3_1 ;
    wire \this_vga_signals.N_6_1_0 ;
    wire \this_vga_signals.N_234 ;
    wire \this_vga_signals.SUM_3_cascade_ ;
    wire \this_vga_signals.g0_6_1 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb1_1 ;
    wire \this_vga_signals.g1_2_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0 ;
    wire \this_vga_signals.SUM_3_0_0 ;
    wire \this_vga_signals.M_pcounter_q_i_3_0 ;
    wire this_vga_signals_hsync_1_i;
    wire this_vga_signals_hvisibility_i;
    wire \this_vga_signals.g3_0_1_cascade_ ;
    wire \this_vga_signals.g3_0 ;
    wire \this_vga_signals.g3_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0_2 ;
    wire \this_vga_signals.g0_0_a2_0_0_cascade_ ;
    wire \this_vga_signals.g1_0_a2_1 ;
    wire \this_vga_signals.vaddress_1_5 ;
    wire \this_vga_signals.mult1_un47_sum_c3_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_x0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_ns ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_ns_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0 ;
    wire \this_vga_signals.g0_i_x4_1 ;
    wire \this_vga_signals.g0_i_x4_0_1 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_0 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_2 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_2_cascade_ ;
    wire \this_vga_signals.g1_0_3 ;
    wire \this_vga_signals.g0_2_0_a2 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c2_0 ;
    wire \this_vga_signals.g0_1_2 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_x1 ;
    wire \this_vga_signals.g1_0 ;
    wire \this_vga_signals.g0_i_x4_2_0_0_1_cascade_ ;
    wire \this_vga_signals.g0_i_x4_0_0 ;
    wire \this_vga_signals.N_3_cascade_ ;
    wire \this_vga_signals.N_4_0_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_c2_0_0_0 ;
    wire \this_vga_signals.g0_2_1 ;
    wire \this_vga_signals.N_5_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_a0_0 ;
    wire \this_vga_signals.SUM_3 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_2 ;
    wire \this_vga_signals.if_N_6_0 ;
    wire bfn_11_13_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_11_14_0_;
    wire \this_vga_signals.un4_hsynclt9 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_pcounter_q_3_1_cascade_ ;
    wire N_3_0;
    wire N_3_0_cascade_;
    wire \this_vga_signals.M_pcounter_q_i_3_1 ;
    wire \this_vga_signals.g1_2 ;
    wire \this_vga_signals.SUM_3_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb1_0 ;
    wire M_this_map_ram_write_data_4;
    wire \this_vga_signals.mult1_un40_sum_axb1_i_0 ;
    wire \this_vga_signals.N_18_cascade_ ;
    wire \this_vga_signals.g1_0_0_1 ;
    wire \this_vga_signals.vaddress_1_6 ;
    wire \this_vga_signals.N_6_cascade_ ;
    wire \this_vga_signals.g1_1_1 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_661_cascade_ ;
    wire \this_vga_signals.g0_2_0_a2_1 ;
    wire \this_vga_signals.if_N_5_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c3_cascade_ ;
    wire \this_vga_signals.N_4_0_1_0 ;
    wire \this_vga_signals.mult1_un47_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_0_cascade_ ;
    wire \this_vga_signals.g0_0_0_a2_0 ;
    wire \this_vga_signals.mult1_un47_sum_c3 ;
    wire \this_vga_signals.mult1_un61_sum_c3 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1_661 ;
    wire \this_vga_signals.g0_i_x4_0_a3_2 ;
    wire \this_vga_signals.vaddress_0_6 ;
    wire \this_vga_signals.g0_i_x4_0_a3_0 ;
    wire \this_vga_signals.vsync_1_3 ;
    wire \this_vga_signals.vsync_1_2_cascade_ ;
    wire this_vga_signals_vsync_1_i;
    wire \this_vga_signals.un2_vsynclt8 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d ;
    wire \this_vga_signals.mult1_un54_sum_0_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.un2_hsynclto3_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_d7lto7_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.M_hcounter_d7lt7_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.N_852_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire \this_vga_signals.un2_hsynclt6_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.un2_hsynclt7 ;
    wire \this_vga_signals.un2_hsynclto3_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.un4_hsynclto7_0 ;
    wire M_this_map_ram_write_data_1;
    wire \this_vga_signals.SUM_2_i_1_1_1_3 ;
    wire \this_vga_signals.N_1_3_1_cascade_ ;
    wire \this_vga_signals.SUM_2_i_1_2_3 ;
    wire \this_vga_signals.SUM_2_i_1_2_3_cascade_ ;
    wire \this_vga_signals.SUM_2_i_1_1_3 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_x0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_N_2L1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_x1 ;
    wire \this_vga_signals.vaddress_5 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1 ;
    wire \this_vga_signals.g2_0_a2_5Z0Z_1_cascade_ ;
    wire \this_vga_signals.g2_0_a2_2 ;
    wire \this_vga_signals.g2_0_a2_5 ;
    wire \this_vga_signals.g2 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire \this_vga_signals.g1_3 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.if_m2 ;
    wire \this_vga_signals.N_1098_1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_0_N_2L1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.vaddress_c3_0 ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_1 ;
    wire \this_vga_signals.M_vcounter_q_7_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.un6_vvisibilitylto8_0_cascade_ ;
    wire \this_vga_signals.un6_vvisibilitylt9_0_cascade_ ;
    wire this_vga_signals_vvisibility_1_cascade_;
    wire \this_vga_signals.vvisibility ;
    wire \this_vga_signals.vaddress_ac0_9_0_a0_0 ;
    wire \this_ppu.N_1195_0_1_cascade_ ;
    wire bfn_14_13_0_;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_6_s1 ;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire port_clk_c;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire bfn_15_9_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_15_10_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire \this_vga_signals.N_852_0 ;
    wire \this_vga_signals.N_1098_g ;
    wire \this_ppu.N_1195_0_cascade_ ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ;
    wire \this_ppu.N_1195_0_1 ;
    wire \this_ppu.M_count_qZ0Z_0 ;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_5 ;
    wire \this_ppu.M_count_qZ0Z_4 ;
    wire \this_ppu.M_count_qZ0Z_6 ;
    wire \this_ppu.M_count_qZ0Z_2 ;
    wire \this_ppu.M_count_qZ0Z_1 ;
    wire \this_ppu.M_count_d_1_sqmuxa_1_i_a2_4_cascade_ ;
    wire \this_ppu.M_count_d_1_sqmuxa_1_i_a2_3 ;
    wire \this_ppu.un16_0 ;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ;
    wire \this_ppu.N_1195_0 ;
    wire \this_ppu.M_count_qZ0Z_3 ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_7 ;
    wire \this_ppu.M_count_qZ0Z_7 ;
    wire \this_vga_signals.N_85_cascade_ ;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_5 ;
    wire \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0Z0Z_2_cascade_ ;
    wire M_this_substate_qZ0;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire M_this_map_ram_write_data_3;
    wire M_this_map_ram_write_data_2;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_vcounter_d7lto8_1 ;
    wire \this_vga_signals.M_vcounter_d7lt8_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire \this_vga_signals.line_clk_1_cascade_ ;
    wire M_this_vga_signals_line_clk_0_cascade_;
    wire \this_vga_signals.un4_lvisibility_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.line_clk_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.M_lcounter_qZ0Z_0 ;
    wire \this_vga_signals.CO0 ;
    wire this_pixel_clk_M_counter_q_i_1;
    wire this_pixel_clk_M_counter_q_0;
    wire \this_vga_signals.N_152_0_cascade_ ;
    wire \this_sprites_ram.mem_WE_6 ;
    wire \this_vga_signals.M_this_state_q_srsts_i_i_1Z0Z_10 ;
    wire \this_sprites_ram.mem_WE_10 ;
    wire this_vga_signals_M_this_state_q_srsts_0_1_i_a2_0_0_1;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_6 ;
    wire \this_vga_signals.N_85 ;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_4 ;
    wire \this_vga_signals.M_this_state_q_srsts_i_1Z0Z_11 ;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0Z0Z_3 ;
    wire M_this_state_d_0_sqmuxa_1;
    wire M_this_map_ram_write_data_7;
    wire GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO;
    wire G_425;
    wire \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ;
    wire \this_vga_signals.M_lcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_vcounter_d8 ;
    wire \this_vga_signals.M_hcounter_d7_0 ;
    wire \this_vga_signals.un1_M_hcounter_d7_1_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire \this_vga_signals.N_153_0_cascade_ ;
    wire N_686_i_cascade_;
    wire N_164;
    wire \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_8 ;
    wire \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_8_cascade_ ;
    wire \this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_8 ;
    wire \this_vga_signals.N_124_0 ;
    wire \this_vga_signals.N_154_cascade_ ;
    wire \this_vga_signals.N_97 ;
    wire \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_2_0 ;
    wire \this_vga_signals.N_154 ;
    wire \this_vga_signals.N_62_cascade_ ;
    wire \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0 ;
    wire M_this_map_ram_read_data_2;
    wire M_this_ppu_sprites_addr_8;
    wire M_this_map_ram_read_data_1;
    wire M_this_ppu_sprites_addr_7;
    wire port_address_in_7;
    wire led_c_1;
    wire N_84;
    wire port_address_in_1;
    wire port_address_in_4;
    wire port_address_in_0;
    wire N_36;
    wire port_dmab_c_i;
    wire \this_ppu.un1_M_oam_idx_q_1_c1_cascade_ ;
    wire \this_ppu.un1_M_oam_idx_q_1_c3_cascade_ ;
    wire \this_ppu.M_count_d_0_sqmuxa_1_7 ;
    wire \this_ppu.un1_M_oam_idx_q_1_c3 ;
    wire \this_ppu.un1_M_oam_idx_q_1_c1 ;
    wire \this_ppu.N_1156_0 ;
    wire M_this_ppu_oam_addr_2;
    wire M_this_ppu_oam_addr_1;
    wire \this_ppu.M_oam_idx_qZ0Z_4 ;
    wire M_this_ppu_oam_addr_0;
    wire \this_ppu.un1_M_haddress_q_3_c2_cascade_ ;
    wire \this_ppu.un1_M_haddress_q_3_c5 ;
    wire \this_sprites_ram.mem_out_bus7_0 ;
    wire \this_sprites_ram.mem_out_bus3_0 ;
    wire \this_ppu.un2_hscroll_axb_0_cascade_ ;
    wire M_this_ppu_sprites_addr_0;
    wire \this_ppu.un1_M_haddress_q_3_c2 ;
    wire \this_ppu.M_state_q_RNIGL6V4Z0Z_0 ;
    wire \this_sprites_ram.mem_out_bus4_3 ;
    wire \this_sprites_ram.mem_out_bus0_3 ;
    wire \this_sprites_ram.mem_WE_8 ;
    wire N_686_i;
    wire M_this_data_count_qlde_i_i;
    wire M_this_data_count_qZ0Z_0;
    wire bfn_18_15_0_;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_data_count_q_cry_0_THRU_CO;
    wire M_this_data_count_q_cry_0;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_q_cry_1_THRU_CO;
    wire M_this_data_count_q_cry_1;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_q_cry_2_THRU_CO;
    wire M_this_data_count_q_cry_2;
    wire M_this_data_count_q_cry_3_THRU_CO;
    wire M_this_data_count_q_cry_3;
    wire M_this_data_count_q_cry_4_THRU_CO;
    wire M_this_data_count_q_cry_4;
    wire M_this_data_count_qZ0Z_6;
    wire M_this_data_count_q_s_6;
    wire M_this_data_count_q_cry_5;
    wire M_this_data_count_qZ0Z_7;
    wire M_this_data_count_q_cry_6_THRU_CO;
    wire M_this_data_count_q_cry_6;
    wire M_this_data_count_q_cry_7;
    wire M_this_data_count_q_cry_7_THRU_CO;
    wire bfn_18_16_0_;
    wire M_this_data_count_q_cry_8_THRU_CO;
    wire M_this_data_count_q_cry_8;
    wire M_this_data_count_qZ0Z_10;
    wire M_this_data_count_q_s_10;
    wire M_this_data_count_q_cry_9;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_q_cry_10_THRU_CO;
    wire M_this_data_count_q_cry_10;
    wire M_this_data_count_qZ0Z_12;
    wire CONSTANT_ONE_NET;
    wire M_this_data_count_q_cry_11_THRU_CO;
    wire M_this_data_count_q_cry_11;
    wire M_this_data_count_qZ0Z_13;
    wire M_this_data_count_q_cry_12;
    wire M_this_data_count_q_s_13;
    wire N_49;
    wire this_vga_signals_vvisibility_1;
    wire \this_ppu.un1_M_vaddress_q_2_c2_cascade_ ;
    wire \this_ppu.un1_M_vaddress_q_2_c5 ;
    wire bfn_18_19_0_;
    wire \this_ppu.un1_M_haddress_q_2_cry_0 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_1 ;
    wire M_this_ppu_map_addr_0;
    wire \this_ppu.un1_M_haddress_q_2_cry_2 ;
    wire M_this_ppu_map_addr_1;
    wire \this_ppu.un1_M_haddress_q_2_cry_3 ;
    wire M_this_ppu_map_addr_2;
    wire \this_ppu.un1_M_haddress_q_2_cry_4 ;
    wire M_this_ppu_map_addr_3;
    wire \this_ppu.un1_M_haddress_q_2_cry_5 ;
    wire M_this_ppu_map_addr_4;
    wire \this_ppu.un1_M_haddress_q_2_cry_6 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_7 ;
    wire bfn_18_20_0_;
    wire \this_ppu.M_state_qZ0Z_3 ;
    wire \this_ppu.un1_M_haddress_q_2_4 ;
    wire \this_ppu.N_148 ;
    wire \this_ppu.vscroll8 ;
    wire \this_ppu.un1_M_haddress_q_2_5 ;
    wire \this_ppu.M_state_qZ0Z_4 ;
    wire M_this_ppu_oam_addr_3;
    wire \this_ppu.N_144_4 ;
    wire \this_ppu.M_state_qZ0Z_2 ;
    wire \this_ppu.N_144 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ;
    wire M_this_ppu_vram_data_0;
    wire M_this_ppu_vram_data_0_cascade_;
    wire \this_ppu.N_156_cascade_ ;
    wire M_this_ppu_vram_en_0;
    wire \this_sprites_ram.mem_out_bus6_3 ;
    wire \this_sprites_ram.mem_out_bus2_3 ;
    wire \this_sprites_ram.mem_out_bus4_0 ;
    wire \this_sprites_ram.mem_out_bus0_0 ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_ ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ;
    wire M_this_map_ram_read_data_7;
    wire \this_sprites_ram.mem_out_bus7_3 ;
    wire \this_sprites_ram.mem_out_bus3_3 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ;
    wire M_this_ppu_vram_data_3;
    wire \this_ppu.N_156 ;
    wire \this_ppu.N_150 ;
    wire \this_ppu.M_state_qZ0Z_5 ;
    wire \this_ppu.M_state_qZ0Z_1 ;
    wire \this_sprites_ram.mem_out_bus5_3 ;
    wire \this_sprites_ram.mem_out_bus1_3 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ;
    wire M_this_state_qZ0Z_10;
    wire M_this_state_q_RNIH92SZ0Z_10_cascade_;
    wire \this_vga_signals.N_83 ;
    wire \this_vga_signals.N_94_0 ;
    wire \this_vga_signals.N_94_0_cascade_ ;
    wire \this_vga_signals.M_this_state_q_srsts_i_i_0Z0Z_12 ;
    wire M_this_state_q_RNI373A1Z0Z_8;
    wire this_vga_signals_un21_i_a3_1_1_cascade_;
    wire port_dmab_c;
    wire M_this_data_count_qZ0Z_8;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_qZ0Z_9;
    wire M_this_data_count_qZ0Z_4;
    wire \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_8 ;
    wire \this_vga_signals.M_this_state_q_srsts_i_a3_0_7_cascade_ ;
    wire \this_vga_signals.M_this_state_q_srsts_i_0Z0Z_7_cascade_ ;
    wire M_this_state_q_RNI6Q0SZ0Z_5;
    wire M_this_state_qZ0Z_12;
    wire N_848;
    wire \this_vga_signals.N_93_0 ;
    wire \this_ppu.M_state_qZ0Z_0 ;
    wire M_this_vga_signals_line_clk_0;
    wire \this_ppu.M_last_q ;
    wire \this_ppu.N_132_0 ;
    wire \this_ppu.un1_M_vaddress_q_2_c2 ;
    wire \this_ppu.M_state_q_RNILG0GDZ0Z_0 ;
    wire bfn_19_17_0_;
    wire \this_ppu.un1_M_vaddress_q_3_cry_0 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_1 ;
    wire M_this_ppu_map_addr_5;
    wire \this_ppu.un1_M_vaddress_q_3_cry_2 ;
    wire M_this_ppu_map_addr_6;
    wire \this_ppu.un1_M_vaddress_q_3_cry_3 ;
    wire M_this_ppu_map_addr_7;
    wire \this_ppu.un1_M_vaddress_q_3_cry_4 ;
    wire M_this_ppu_map_addr_8;
    wire \this_ppu.un1_M_vaddress_q_3_cry_5 ;
    wire M_this_ppu_map_addr_9;
    wire \this_ppu.un1_M_vaddress_q_3_cry_6 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_7 ;
    wire bfn_19_18_0_;
    wire \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO ;
    wire \this_reset_cond.M_stage_qZ0Z_3 ;
    wire \this_ppu.M_this_ppu_vram_addr_i_0 ;
    wire bfn_19_19_0_;
    wire \this_ppu.M_this_ppu_vram_addr_i_1 ;
    wire \this_ppu.un1_M_haddress_q_cry_0 ;
    wire \this_ppu.M_this_ppu_vram_addr_i_2 ;
    wire \this_ppu.un1_M_haddress_q_cry_1 ;
    wire \this_ppu.M_this_ppu_map_addr_i_0 ;
    wire \this_ppu.un1_M_haddress_q_cry_2 ;
    wire \this_ppu.M_this_ppu_map_addr_i_1 ;
    wire \this_ppu.un1_M_haddress_q_cry_3 ;
    wire \this_ppu.M_this_ppu_map_addr_i_2 ;
    wire \this_ppu.un1_M_haddress_q_cry_4 ;
    wire \this_ppu.M_this_ppu_map_addr_i_3 ;
    wire \this_ppu.un1_M_haddress_q_cry_5 ;
    wire \this_ppu.M_this_ppu_map_addr_i_4 ;
    wire \this_ppu.un1_M_haddress_q_cry_6 ;
    wire \this_ppu.un1_M_haddress_q_cry_7 ;
    wire bfn_19_20_0_;
    wire \this_ppu.vscroll8_1 ;
    wire \this_ppu.un1_M_vaddress_q_3_4 ;
    wire \this_sprites_ram.mem_out_bus4_1 ;
    wire \this_sprites_ram.mem_out_bus0_1 ;
    wire \this_sprites_ram.mem_out_bus7_1 ;
    wire \this_sprites_ram.mem_out_bus3_1 ;
    wire M_this_map_ram_read_data_6;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ;
    wire M_this_ppu_vram_data_1;
    wire \this_sprites_ram.mem_out_bus7_2 ;
    wire \this_sprites_ram.mem_out_bus3_2 ;
    wire \this_sprites_ram.mem_out_bus4_2 ;
    wire \this_sprites_ram.mem_out_bus0_2 ;
    wire \this_sprites_ram.mem_radregZ0Z_12 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ;
    wire M_this_ppu_vram_data_2;
    wire M_this_map_ram_read_data_0;
    wire M_this_ppu_sprites_addr_6;
    wire \this_sprites_ram.mem_out_bus6_2 ;
    wire \this_sprites_ram.mem_out_bus2_2 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ;
    wire N_792;
    wire M_this_sprites_address_qc_0_0_0;
    wire N_795;
    wire N_773_0;
    wire N_773_0_cascade_;
    wire \this_vga_signals.N_485 ;
    wire N_17;
    wire N_126;
    wire M_this_state_qZ0Z_7;
    wire port_dmab_ac0_1_3_cascade_;
    wire port_dmab_ac0_1_4;
    wire N_15;
    wire N_809_cascade_;
    wire M_this_state_qZ0Z_5;
    wire M_this_state_qZ0Z_8;
    wire M_this_state_qZ0Z_1;
    wire N_775_0;
    wire N_775_0_cascade_;
    wire port_address_in_5;
    wire \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0Z0Z_0 ;
    wire N_87_0_cascade_;
    wire M_this_state_qZ0Z_6;
    wire port_enb_c;
    wire this_start_data_delay_M_last_q;
    wire \this_reset_cond.M_stage_qZ0Z_4 ;
    wire M_this_state_qZ0Z_11;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire M_this_delay_clk_out_0;
    wire \this_ppu.M_this_ppu_vram_addr_i_7 ;
    wire bfn_20_19_0_;
    wire \this_ppu.M_vaddress_q_i_1 ;
    wire \this_ppu.un1_M_vaddress_q_cry_0 ;
    wire \this_ppu.M_vaddress_q_i_2 ;
    wire \this_ppu.un1_M_vaddress_q_cry_1 ;
    wire \this_ppu.M_this_ppu_map_addr_i_5 ;
    wire \this_ppu.un1_M_vaddress_q_cry_2 ;
    wire \this_ppu.M_this_ppu_map_addr_i_6 ;
    wire \this_ppu.un1_M_vaddress_q_cry_3 ;
    wire \this_ppu.M_this_ppu_map_addr_i_7 ;
    wire \this_ppu.un1_M_vaddress_q_cry_4 ;
    wire \this_ppu.M_this_ppu_map_addr_i_8 ;
    wire \this_ppu.un1_M_vaddress_q_cry_5 ;
    wire \this_ppu.M_this_ppu_map_addr_i_9 ;
    wire \this_ppu.un1_M_vaddress_q_cry_6 ;
    wire \this_ppu.un1_M_vaddress_q_cry_7 ;
    wire bfn_20_20_0_;
    wire \this_ppu.un1_M_vaddress_q_cry_7_THRU_CO ;
    wire M_this_map_ram_read_data_5;
    wire \this_sprites_ram.mem_radregZ0Z_11 ;
    wire M_this_state_qZ0Z_13;
    wire \this_sprites_ram.mem_out_bus6_1 ;
    wire \this_sprites_ram.mem_out_bus2_1 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus5_2 ;
    wire \this_sprites_ram.mem_out_bus1_2 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ;
    wire \this_sprites_ram.mem_out_bus5_0 ;
    wire \this_sprites_ram.mem_out_bus1_0 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ;
    wire M_this_sprites_address_qc_0_0;
    wire \this_sprites_ram.mem_WE_14 ;
    wire M_this_sprites_address_qZ0Z_0;
    wire N_443_i;
    wire M_this_sprites_address_q_RNO_0Z0Z_0;
    wire bfn_21_13_0_;
    wire un1_M_this_sprites_address_q_cry_0;
    wire un1_M_this_sprites_address_q_cry_1;
    wire un1_M_this_sprites_address_q_cry_2;
    wire un1_M_this_sprites_address_q_cry_3;
    wire un1_M_this_sprites_address_q_cry_4;
    wire un1_M_this_sprites_address_q_cry_5;
    wire un1_M_this_sprites_address_q_cry_6;
    wire un1_M_this_sprites_address_q_cry_7;
    wire bfn_21_14_0_;
    wire un1_M_this_sprites_address_q_cry_8;
    wire M_this_sprites_address_qZ0Z_10;
    wire M_this_sprites_address_q_RNO_1Z0Z_10;
    wire un1_M_this_sprites_address_q_cry_9;
    wire M_this_sprites_address_q_RNO_1Z0Z_11;
    wire un1_M_this_sprites_address_q_cry_10;
    wire un1_M_this_sprites_address_q_cry_11;
    wire M_this_sprites_address_qc_2_1;
    wire un1_M_this_sprites_address_q_cry_12;
    wire M_this_sprites_address_q_RNO_0Z0Z_12;
    wire N_807_cascade_;
    wire M_this_sprites_address_q_RNO_1Z0Z_7;
    wire M_this_sprites_address_q_RNO_1Z0Z_8;
    wire N_803_cascade_;
    wire M_this_sprites_address_qc_10_0;
    wire M_this_sprites_address_qZ0Z_8;
    wire N_602;
    wire M_this_state_qZ0Z_9;
    wire M_this_state_qZ0Z_3;
    wire M_this_sprites_address_qZ0Z_7;
    wire M_this_sprites_address_qc_9_0;
    wire M_this_oam_ram_read_data_i_19;
    wire M_this_oam_ram_read_data_i_11;
    wire M_this_oam_ram_read_data_15;
    wire \this_ppu.un1_M_haddress_q_2_7 ;
    wire M_this_oam_address_qZ0Z_4;
    wire un1_M_this_oam_address_q_c4;
    wire M_this_oam_address_qZ0Z_5;
    wire M_this_oam_address_qZ0Z_3;
    wire M_this_data_tmp_qZ0Z_2;
    wire N_746_0;
    wire M_this_oam_ram_write_data_28;
    wire M_this_state_qZ0Z_4;
    wire un1_M_this_sprites_address_q_cry_0_THRU_CO;
    wire M_this_sprites_address_q_RNO_0Z0Z_2;
    wire N_813;
    wire N_799;
    wire M_this_sprites_address_qc_11_0_cascade_;
    wire M_this_sprites_address_q_RNO_1Z0Z_9;
    wire M_this_sprites_address_qZ0Z_9;
    wire M_this_sprites_address_q_RNO_0Z0Z_3;
    wire M_this_sprites_address_qZ0Z_3;
    wire N_50;
    wire M_this_ppu_sprites_addr_3;
    wire M_this_sprites_address_qZ0Z_2;
    wire N_103;
    wire M_this_sprites_ram_write_data_iv_i_i_1;
    wire port_address_in_3;
    wire port_address_in_2;
    wire port_rw_in;
    wire port_address_in_6;
    wire \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_4_0 ;
    wire N_54_0;
    wire \this_ppu.un1_oam_data_1_c2 ;
    wire N_163;
    wire un1_M_this_oam_address_q_c2;
    wire M_this_oam_address_qZ0Z_2;
    wire N_1190_0;
    wire M_this_data_tmp_qZ0Z_6;
    wire N_742_0;
    wire N_34_0;
    wire M_this_data_tmp_qZ0Z_4;
    wire N_744_0;
    wire M_this_data_tmp_qZ0Z_7;
    wire N_56_0;
    wire M_this_data_tmp_qZ0Z_16;
    wire N_738_0;
    wire M_this_data_tmp_qZ0Z_22;
    wire N_40_0;
    wire \this_sprites_ram.mem_out_bus6_0 ;
    wire \this_sprites_ram.mem_out_bus2_0 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ;
    wire N_102;
    wire M_this_sprites_address_q_RNO_0Z0Z_4;
    wire M_this_sprites_address_qZ0Z_4;
    wire N_101_cascade_;
    wire M_this_sprites_address_q_RNO_0Z0Z_6;
    wire M_this_sprites_address_qZ0Z_6;
    wire \this_vga_signals.M_this_sprites_address_q_3_bmZ0Z_1 ;
    wire M_this_sprites_address_qZ0Z_1;
    wire M_this_state_qZ0Z_2;
    wire N_87_0;
    wire \this_vga_signals.M_this_sprites_address_q_3_amZ0Z_1 ;
    wire \this_vga_signals.un1_M_this_state_q_3_0_i_0_0 ;
    wire \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2 ;
    wire M_this_sprites_ram_write_data_iv_i_i_3;
    wire \this_ppu.un2_vscroll_axb_0 ;
    wire M_this_ppu_sprites_addr_1;
    wire M_this_data_tmp_qZ0Z_8;
    wire N_1182_0;
    wire M_this_data_tmp_qZ0Z_3;
    wire N_745_0;
    wire M_this_data_tmp_qZ0Z_14;
    wire N_739_0;
    wire M_this_data_tmp_qZ0Z_5;
    wire N_743_0;
    wire N_32_0;
    wire M_this_data_tmp_qZ0Z_11;
    wire M_this_oam_ram_write_data_11;
    wire M_this_data_tmp_qZ0Z_0;
    wire N_748_0;
    wire N_44_0;
    wire M_this_data_tmp_qZ0Z_17;
    wire N_1174_0;
    wire M_this_data_tmp_qZ0Z_23;
    wire M_this_oam_ram_write_data_23;
    wire M_this_data_tmp_qZ0Z_20;
    wire N_42_0;
    wire M_this_oam_ram_write_data_30;
    wire \this_sprites_ram.mem_out_bus5_1 ;
    wire \this_sprites_ram.mem_out_bus1_1 ;
    wire \this_sprites_ram.mem_radregZ0Z_13 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ;
    wire M_this_ppu_sprites_addr_2;
    wire \this_sprites_ram.mem_WE_4 ;
    wire \this_sprites_ram.mem_WE_12 ;
    wire M_this_ppu_sprites_addr_5;
    wire N_809;
    wire M_this_sprites_address_q_RNO_0Z0Z_5;
    wire N_595;
    wire N_383_0;
    wire M_this_sprites_address_qZ0Z_5;
    wire N_515_g;
    wire \this_sprites_ram.mem_WE_0 ;
    wire M_this_ppu_sprites_addr_4;
    wire M_this_ppu_vram_addr_7;
    wire M_this_oam_ram_read_data_16;
    wire \this_ppu.M_this_oam_ram_read_data_i_16 ;
    wire bfn_24_16_0_;
    wire \this_ppu.M_vaddress_qZ0Z_1 ;
    wire \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0 ;
    wire \this_ppu.un2_vscroll_cry_0 ;
    wire \this_ppu.M_vaddress_qZ0Z_2 ;
    wire M_this_oam_ram_read_data_18;
    wire \this_ppu.un2_vscroll_cry_1 ;
    wire \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0 ;
    wire M_this_map_ram_read_data_4;
    wire M_this_ppu_sprites_addr_10;
    wire M_this_sprites_address_qZ0Z_11;
    wire M_this_sprites_address_qZ0Z_12;
    wire M_this_sprites_address_qZ0Z_13;
    wire N_23_0;
    wire \this_sprites_ram.mem_WE_2 ;
    wire M_this_ppu_vram_addr_0;
    wire M_this_oam_ram_read_data_8;
    wire \this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ;
    wire bfn_24_19_0_;
    wire M_this_ppu_vram_addr_1;
    wire \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0 ;
    wire \this_ppu.un2_hscroll_cry_0 ;
    wire M_this_ppu_vram_addr_2;
    wire M_this_oam_ram_read_data_10;
    wire \this_ppu.un2_hscroll_cry_1 ;
    wire \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0 ;
    wire M_this_oam_ram_read_data_9;
    wire M_this_oam_ram_read_data_i_9;
    wire M_this_data_tmp_qZ0Z_1;
    wire N_747_0;
    wire M_this_data_tmp_qZ0Z_10;
    wire M_this_oam_ram_write_data_10;
    wire M_this_map_ram_read_data_3;
    wire \this_ppu.M_state_qZ0Z_6 ;
    wire \this_ppu.M_state_qZ0Z_7 ;
    wire M_this_ppu_sprites_addr_9;
    wire M_this_data_tmp_qZ0Z_12;
    wire N_740_0;
    wire M_this_oam_ram_read_data_13;
    wire M_this_oam_ram_read_data_12;
    wire M_this_oam_ram_read_data_14;
    wire M_this_oam_ram_read_data_11;
    wire \this_ppu.un1_M_haddress_q_2_6 ;
    wire M_this_data_tmp_qZ0Z_19;
    wire M_this_oam_ram_write_data_19;
    wire M_this_oam_ram_read_data_6;
    wire M_this_oam_ram_read_data_5;
    wire M_this_oam_ram_read_data_7;
    wire M_this_oam_ram_read_data_4;
    wire \this_ppu.un9lto7Z0Z_4 ;
    wire M_this_data_tmp_qZ0Z_9;
    wire N_741_0;
    wire M_this_oam_ram_read_data_23;
    wire \this_ppu.un1_oam_data_c2_cascade_ ;
    wire \this_ppu.un1_M_vaddress_q_3_7 ;
    wire M_this_data_tmp_qZ0Z_13;
    wire M_this_oam_ram_write_data_13;
    wire M_this_data_tmp_qZ0Z_15;
    wire M_this_oam_ram_write_data_15;
    wire N_123_0;
    wire M_this_oam_ram_read_data_2;
    wire M_this_oam_ram_read_data_1;
    wire M_this_oam_ram_read_data_3;
    wire M_this_oam_ram_read_data_0;
    wire \this_ppu.un9lto7Z0Z_5 ;
    wire M_this_oam_ram_read_data_17;
    wire M_this_oam_ram_read_data_i_17;
    wire M_this_data_tmp_qZ0Z_18;
    wire M_this_oam_ram_write_data_18;
    wire \this_ppu.un1_M_vaddress_q_3_5 ;
    wire N_38_0;
    wire M_this_oam_ram_write_data_31;
    wire N_736_0;
    wire N_737_0;
    wire M_this_oam_ram_read_data_21;
    wire M_this_oam_ram_read_data_20;
    wire M_this_oam_ram_read_data_22;
    wire M_this_oam_ram_read_data_19;
    wire \this_ppu.un1_M_vaddress_q_3_6 ;
    wire M_this_oam_address_qZ0Z_0;
    wire M_this_oam_address_qZ0Z_1;
    wire M_this_data_tmp_qZ0Z_21;
    wire N_122_0;
    wire M_this_oam_ram_write_data_21;
    wire \this_reset_cond.M_stage_qZ0Z_5 ;
    wire \this_reset_cond.M_stage_qZ0Z_6 ;
    wire \this_reset_cond.M_stage_qZ0Z_7 ;
    wire un1_M_this_state_q_9_0_i;
    wire M_this_external_address_qZ0Z_0;
    wire bfn_28_21_0_;
    wire M_this_external_address_qZ0Z_1;
    wire un1_M_this_external_address_q_cry_0;
    wire M_this_external_address_qZ0Z_2;
    wire un1_M_this_external_address_q_cry_1;
    wire M_this_external_address_qZ0Z_3;
    wire un1_M_this_external_address_q_cry_2;
    wire M_this_external_address_qZ0Z_4;
    wire un1_M_this_external_address_q_cry_3;
    wire M_this_external_address_qZ0Z_5;
    wire un1_M_this_external_address_q_cry_4;
    wire M_this_external_address_qZ0Z_6;
    wire un1_M_this_external_address_q_cry_5;
    wire M_this_external_address_qZ0Z_7;
    wire un1_M_this_external_address_q_cry_6;
    wire un1_M_this_external_address_q_cry_7;
    wire port_data_c_0;
    wire M_this_external_address_qZ0Z_8;
    wire bfn_28_22_0_;
    wire port_data_c_1;
    wire M_this_external_address_qZ0Z_9;
    wire un1_M_this_external_address_q_cry_8;
    wire port_data_c_2;
    wire M_this_external_address_qZ0Z_10;
    wire un1_M_this_external_address_q_cry_9;
    wire port_data_c_3;
    wire M_this_external_address_qZ0Z_11;
    wire un1_M_this_external_address_q_cry_10;
    wire port_data_c_4;
    wire M_this_external_address_qZ0Z_12;
    wire un1_M_this_external_address_q_cry_11;
    wire port_data_c_5;
    wire M_this_external_address_qZ0Z_13;
    wire un1_M_this_external_address_q_cry_12;
    wire port_data_c_6;
    wire M_this_external_address_qZ0Z_14;
    wire un1_M_this_external_address_q_cry_13;
    wire N_749_0;
    wire port_data_c_7;
    wire un1_M_this_external_address_q_cry_14;
    wire M_this_external_address_qZ0Z_15;
    wire M_this_reset_cond_out_g_0;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_8 ;
    wire M_this_reset_cond_out_0;
    wire clk_0_c_g;
    wire _gnd_net_;

    defparam \this_map_ram.mem_mem_0_0_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_0_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,M_this_map_ram_read_data_3,dangling_wire_2,dangling_wire_3,dangling_wire_4,M_this_map_ram_read_data_2,dangling_wire_5,dangling_wire_6,dangling_wire_7,M_this_map_ram_read_data_1,dangling_wire_8,dangling_wire_9,dangling_wire_10,M_this_map_ram_read_data_0,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__22140,N__21819,N__21867,N__21906,N__21957,N__20424,N__20490,N__20568,N__20631,N__20271}),
            .WADDR({dangling_wire_13,N__11217,N__11250,N__11280,N__11310,N__11340,N__11370,N__11022,N__11052,N__11082,N__11109}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__16197,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__16185,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__13986,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__11958,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__34633),
            .RE(N__19658),
            .WCLKE(N__17434),
            .WCLK(N__34634),
            .WE(N__19667));
    defparam \this_map_ram.mem_mem_0_1_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_1_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_42,dangling_wire_43,M_this_map_ram_read_data_7,dangling_wire_44,dangling_wire_45,dangling_wire_46,M_this_map_ram_read_data_6,dangling_wire_47,dangling_wire_48,dangling_wire_49,M_this_map_ram_read_data_5,dangling_wire_50,dangling_wire_51,dangling_wire_52,M_this_map_ram_read_data_4,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__22134,N__21813,N__21861,N__21900,N__21951,N__20418,N__20484,N__20562,N__20625,N__20265}),
            .WADDR({dangling_wire_55,N__11211,N__11244,N__11274,N__11304,N__11334,N__11364,N__11016,N__11046,N__11076,N__11103}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__17331,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__11940,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__11952,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__13215,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__34640),
            .RE(N__19581),
            .WCLKE(N__17435),
            .WCLK(N__34641),
            .WE(N__19617));
    defparam \this_oam_ram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_0_physical  (
            .RDATA({M_this_oam_ram_read_data_15,M_this_oam_ram_read_data_14,M_this_oam_ram_read_data_13,M_this_oam_ram_read_data_12,M_this_oam_ram_read_data_11,M_this_oam_ram_read_data_10,M_this_oam_ram_read_data_9,M_this_oam_ram_read_data_8,M_this_oam_ram_read_data_7,M_this_oam_ram_read_data_6,M_this_oam_ram_read_data_5,M_this_oam_ram_read_data_4,M_this_oam_ram_read_data_3,M_this_oam_ram_read_data_2,M_this_oam_ram_read_data_1,M_this_oam_ram_read_data_0}),
            .RADDR({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,N__20862,N__19056,N__19011,N__18954}),
            .WADDR({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__24822,N__24876,N__24789,N__26421}),
            .MASK({dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113}),
            .WDATA({N__32043,N__28149,N__32067,N__31074,N__28383,N__31713,N__32130,N__26517,N__26931,N__26343,N__28125,N__26952,N__28173,N__25278,N__31734,N__28362}),
            .RCLKE(),
            .RCLK(N__34629),
            .RE(N__19822),
            .WCLKE(N__32033),
            .WCLK(N__34630),
            .WE(N__19746));
    defparam \this_oam_ram.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,M_this_oam_ram_read_data_23,M_this_oam_ram_read_data_22,M_this_oam_ram_read_data_21,M_this_oam_ram_read_data_20,M_this_oam_ram_read_data_19,M_this_oam_ram_read_data_18,M_this_oam_ram_read_data_17,M_this_oam_ram_read_data_16}),
            .RADDR({dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__20856,N__19050,N__19005,N__18948}),
            .WADDR({dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,N__24816,N__24870,N__24783,N__26415}),
            .MASK({dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151}),
            .WDATA({N__33093,N__29685,N__33087,N__25263,N__28407,N__26331,N__33081,N__33102,N__28260,N__26889,N__32265,N__28239,N__30867,N__33132,N__28350,N__26910}),
            .RCLKE(),
            .RCLK(N__34635),
            .RE(N__19744),
            .WCLKE(N__32037),
            .WCLK(N__34636),
            .WE(N__19745));
    defparam \this_sprites_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,\this_sprites_ram.mem_out_bus0_1 ,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,\this_sprites_ram.mem_out_bus0_0 ,dangling_wire_163,dangling_wire_164,dangling_wire_165}),
            .RADDR({N__30493,N__31334,N__18325,N__18096,N__22535,N__29315,N__28591,N__25785,N__29522,N__27180,N__18858}),
            .WADDR({N__24366,N__26227,N__24711,N__25169,N__28101,N__28859,N__26821,N__26000,N__25544,N__27891,N__23988}),
            .MASK({dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181}),
            .WDATA({dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,N__25370,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,N__22818,dangling_wire_193,dangling_wire_194,dangling_wire_195}),
            .RCLKE(),
            .RCLK(N__34518),
            .RE(N__20100),
            .WCLKE(N__24018),
            .WCLK(N__34519),
            .WE(N__20012));
    defparam \this_sprites_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,\this_sprites_ram.mem_out_bus0_3 ,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,\this_sprites_ram.mem_out_bus0_2 ,dangling_wire_207,dangling_wire_208,dangling_wire_209}),
            .RADDR({N__30475,N__31314,N__18313,N__18092,N__22487,N__29297,N__28592,N__25784,N__29521,N__27179,N__18854}),
            .WADDR({N__24365,N__26208,N__24707,N__25157,N__28100,N__28858,N__26820,N__26019,N__25590,N__27890,N__23987}),
            .MASK({dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225}),
            .WDATA({dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,N__27273,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,N__23100,dangling_wire_237,dangling_wire_238,dangling_wire_239}),
            .RCLKE(),
            .RCLK(N__34528),
            .RE(N__19887),
            .WCLKE(N__24017),
            .WCLK(N__34529),
            .WE(N__20092));
    defparam \this_sprites_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,\this_sprites_ram.mem_out_bus1_1 ,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,\this_sprites_ram.mem_out_bus1_0 ,dangling_wire_251,dangling_wire_252,dangling_wire_253}),
            .RADDR({N__30474,N__31325,N__18292,N__18085,N__22530,N__29299,N__28570,N__25776,N__29503,N__27172,N__18844}),
            .WADDR({N__24357,N__26207,N__24698,N__25170,N__28091,N__28838,N__26801,N__26004,N__25584,N__27877,N__23977}),
            .MASK({dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269}),
            .WDATA({dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,N__25362,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,N__22813,dangling_wire_281,dangling_wire_282,dangling_wire_283}),
            .RCLKE(),
            .RCLK(N__34542),
            .RE(N__20097),
            .WCLKE(N__29343),
            .WCLK(N__34543),
            .WE(N__20091));
    defparam \this_sprites_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,\this_sprites_ram.mem_out_bus1_3 ,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,\this_sprites_ram.mem_out_bus1_2 ,dangling_wire_295,dangling_wire_296,dangling_wire_297}),
            .RADDR({N__30453,N__31291,N__18327,N__18075,N__22506,N__29268,N__28574,N__25761,N__29499,N__27161,N__18843}),
            .WADDR({N__24343,N__26182,N__24679,N__25114,N__28090,N__28837,N__26800,N__25977,N__25569,N__27876,N__23976}),
            .MASK({dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313}),
            .WDATA({dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,N__27276,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,N__23095,dangling_wire_325,dangling_wire_326,dangling_wire_327}),
            .RCLKE(),
            .RCLK(N__34558),
            .RE(N__20096),
            .WCLKE(N__29342),
            .WCLK(N__34559),
            .WE(N__20057));
    defparam \this_sprites_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,\this_sprites_ram.mem_out_bus2_1 ,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,\this_sprites_ram.mem_out_bus2_0 ,dangling_wire_339,dangling_wire_340,dangling_wire_341}),
            .RADDR({N__30452,N__31307,N__18321,N__18063,N__22511,N__29277,N__28540,N__25739,N__29474,N__27144,N__18816}),
            .WADDR({N__24319,N__26181,N__24650,N__25155,N__28065,N__28806,N__26749,N__26005,N__25547,N__27842,N__23950}),
            .MASK({dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357}),
            .WDATA({dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,N__25349,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,N__22800,dangling_wire_369,dangling_wire_370,dangling_wire_371}),
            .RCLKE(),
            .RCLK(N__34573),
            .RE(N__20068),
            .WCLKE(N__16955),
            .WCLK(N__34572),
            .WE(N__20056));
    defparam \this_sprites_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,\this_sprites_ram.mem_out_bus2_3 ,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,\this_sprites_ram.mem_out_bus2_2 ,dangling_wire_383,dangling_wire_384,dangling_wire_385}),
            .RADDR({N__30519,N__31335,N__18326,N__18021,N__22527,N__29325,N__28608,N__25783,N__29547,N__27097,N__18832}),
            .WADDR({N__24356,N__26238,N__24706,N__25168,N__28099,N__28869,N__26822,N__26021,N__25589,N__27888,N__23985}),
            .MASK({dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,dangling_wire_401}),
            .WDATA({dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,N__27275,dangling_wire_406,dangling_wire_407,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,N__23099,dangling_wire_413,dangling_wire_414,dangling_wire_415}),
            .RCLKE(),
            .RCLK(N__34550),
            .RE(N__20080),
            .WCLKE(N__16962),
            .WCLK(N__34551),
            .WE(N__20076));
    defparam \this_sprites_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,\this_sprites_ram.mem_out_bus3_1 ,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,\this_sprites_ram.mem_out_bus3_0 ,dangling_wire_427,dangling_wire_428,dangling_wire_429}),
            .RADDR({N__30515,N__31261,N__18248,N__18020,N__22525,N__29324,N__28604,N__25772,N__29543,N__27160,N__18831}),
            .WADDR({N__24339,N__26237,N__24705,N__25158,N__28086,N__28868,N__26811,N__26020,N__25588,N__27887,N__23984}),
            .MASK({dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,dangling_wire_445}),
            .WDATA({dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,N__25371,dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,N__22817,dangling_wire_457,dangling_wire_458,dangling_wire_459}),
            .RCLKE(),
            .RCLK(N__34565),
            .RE(N__19809),
            .WCLKE(N__19080),
            .WCLK(N__34564),
            .WE(N__20075));
    defparam \this_sprites_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,\this_sprites_ram.mem_out_bus3_3 ,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,\this_sprites_ram.mem_out_bus3_2 ,dangling_wire_471,dangling_wire_472,dangling_wire_473}),
            .RADDR({N__30514,N__31330,N__18317,N__18019,N__22528,N__29316,N__28603,N__25771,N__29507,N__27159,N__18790}),
            .WADDR({N__24270,N__26230,N__24691,N__25176,N__28085,N__28861,N__26810,N__26008,N__25577,N__27886,N__23964}),
            .MASK({dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489}),
            .WDATA({dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,N__27274,dangling_wire_494,dangling_wire_495,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,N__23091,dangling_wire_501,dangling_wire_502,dangling_wire_503}),
            .RCLKE(),
            .RCLK(N__34578),
            .RE(N__20023),
            .WCLKE(N__19076),
            .WCLK(N__34579),
            .WE(N__19878));
    defparam \this_sprites_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,\this_sprites_ram.mem_out_bus4_1 ,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,\this_sprites_ram.mem_out_bus4_0 ,dangling_wire_515,dangling_wire_516,dangling_wire_517}),
            .RADDR({N__30507,N__31329,N__18299,N__18018,N__22524,N__29284,N__28593,N__25751,N__29535,N__27137,N__18829}),
            .WADDR({N__24337,N__26228,N__24690,N__25172,N__28083,N__28824,N__26808,N__26018,N__25531,N__27884,N__23963}),
            .MASK({dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,dangling_wire_533}),
            .WDATA({dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,N__25366,dangling_wire_538,dangling_wire_539,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,N__22807,dangling_wire_545,dangling_wire_546,dangling_wire_547}),
            .RCLKE(),
            .RCLK(N__34592),
            .RE(N__20013),
            .WCLKE(N__16995),
            .WCLK(N__34593),
            .WE(N__19877));
    defparam \this_sprites_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,\this_sprites_ram.mem_out_bus4_3 ,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,\this_sprites_ram.mem_out_bus4_2 ,dangling_wire_559,dangling_wire_560,dangling_wire_561}),
            .RADDR({N__30494,N__31315,N__18272,N__18017,N__22526,N__29323,N__28578,N__25701,N__29542,N__27171,N__18830}),
            .WADDR({N__24338,N__26229,N__24689,N__25171,N__28084,N__28860,N__26809,N__26022,N__25576,N__27885,N__23925}),
            .MASK({dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,dangling_wire_577}),
            .WDATA({dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,N__27262,dangling_wire_582,dangling_wire_583,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,N__23077,dangling_wire_589,dangling_wire_590,dangling_wire_591}),
            .RCLKE(),
            .RCLK(N__34603),
            .RE(N__19865),
            .WCLKE(N__16991),
            .WCLK(N__34604),
            .WE(N__19802));
    defparam \this_sprites_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,\this_sprites_ram.mem_out_bus5_1 ,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,\this_sprites_ram.mem_out_bus5_0 ,dangling_wire_603,dangling_wire_604,dangling_wire_605}),
            .RADDR({N__30428,N__31262,N__18306,N__18051,N__22464,N__29229,N__28547,N__25713,N__29419,N__27122,N__18789}),
            .WADDR({N__24215,N__26150,N__24616,N__25130,N__28064,N__28805,N__26750,N__25983,N__25519,N__27855,N__23949}),
            .MASK({dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,dangling_wire_621}),
            .WDATA({dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,N__25348,dangling_wire_626,dangling_wire_627,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,N__22811,dangling_wire_633,dangling_wire_634,dangling_wire_635}),
            .RCLKE(),
            .RCLK(N__34586),
            .RE(N__20067),
            .WCLKE(N__29354),
            .WCLK(N__34587),
            .WE(N__20085));
    defparam \this_sprites_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,\this_sprites_ram.mem_out_bus5_3 ,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,\this_sprites_ram.mem_out_bus5_2 ,dangling_wire_647,dangling_wire_648,dangling_wire_649}),
            .RADDR({N__30427,N__31281,N__18282,N__18038,N__22507,N__29191,N__28504,N__25682,N__29455,N__27098,N__18803}),
            .WADDR({N__24283,N__26141,N__24642,N__25129,N__28020,N__28730,N__26748,N__25984,N__25471,N__27831,N__23948}),
            .MASK({dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,dangling_wire_665}),
            .WDATA({dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,N__27251,dangling_wire_670,dangling_wire_671,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,N__23072,dangling_wire_677,dangling_wire_678,dangling_wire_679}),
            .RCLKE(),
            .RCLK(N__34599),
            .RE(N__20099),
            .WCLKE(N__29361),
            .WCLK(N__34600),
            .WE(N__19987));
    defparam \this_sprites_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,\this_sprites_ram.mem_out_bus6_1 ,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,\this_sprites_ram.mem_out_bus6_0 ,dangling_wire_691,dangling_wire_692,dangling_wire_693}),
            .RADDR({N__30394,N__31227,N__18249,N__18022,N__22480,N__29236,N__28469,N__25651,N__29491,N__27073,N__18833}),
            .WADDR({N__24297,N__26142,N__24603,N__25127,N__28039,N__28765,N__26790,N__25982,N__25511,N__27832,N__23938}),
            .MASK({dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,dangling_wire_709}),
            .WDATA({dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,N__25330,dangling_wire_714,dangling_wire_715,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,N__22793,dangling_wire_721,dangling_wire_722,dangling_wire_723}),
            .RCLKE(),
            .RCLK(N__34607),
            .RE(N__19913),
            .WCLKE(N__29985),
            .WCLK(N__34608),
            .WE(N__20087));
    defparam \this_sprites_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_724,dangling_wire_725,dangling_wire_726,dangling_wire_727,\this_sprites_ram.mem_out_bus6_3 ,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,\this_sprites_ram.mem_out_bus6_2 ,dangling_wire_735,dangling_wire_736,dangling_wire_737}),
            .RADDR({N__30367,N__31248,N__18180,N__17999,N__22529,N__29272,N__28514,N__25694,N__29492,N__27046,N__18851}),
            .WADDR({N__24332,N__26143,N__24643,N__25128,N__28078,N__28819,N__26815,N__25981,N__25512,N__27871,N__23971}),
            .MASK({dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741,dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,dangling_wire_753}),
            .WDATA({dangling_wire_754,dangling_wire_755,dangling_wire_756,dangling_wire_757,N__27252,dangling_wire_758,dangling_wire_759,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,N__23073,dangling_wire_765,dangling_wire_766,dangling_wire_767}),
            .RCLKE(),
            .RCLK(N__34613),
            .RE(N__20042),
            .WCLKE(N__29984),
            .WCLK(N__34614),
            .WE(N__20086));
    defparam \this_sprites_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_768,dangling_wire_769,dangling_wire_770,dangling_wire_771,\this_sprites_ram.mem_out_bus7_1 ,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,\this_sprites_ram.mem_out_bus7_0 ,dangling_wire_779,dangling_wire_780,dangling_wire_781}),
            .RADDR({N__30425,N__31190,N__18261,N__18034,N__22531,N__29273,N__28554,N__25725,N__29519,N__27020,N__18852}),
            .WADDR({N__24333,N__26179,N__24677,N__25113,N__28079,N__28820,N__26816,N__26006,N__25545,N__27872,N__23972}),
            .MASK({dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785,dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,dangling_wire_797}),
            .WDATA({dangling_wire_798,dangling_wire_799,dangling_wire_800,dangling_wire_801,N__25342,dangling_wire_802,dangling_wire_803,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,N__22812,dangling_wire_809,dangling_wire_810,dangling_wire_811}),
            .RCLKE(),
            .RCLK(N__34620),
            .RE(N__20046),
            .WCLKE(N__28625),
            .WCLK(N__34621),
            .WE(N__19986));
    defparam \this_sprites_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_812,dangling_wire_813,dangling_wire_814,dangling_wire_815,\this_sprites_ram.mem_out_bus7_3 ,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,\this_sprites_ram.mem_out_bus7_2 ,dangling_wire_823,dangling_wire_824,dangling_wire_825}),
            .RADDR({N__30426,N__31133,N__18262,N__18050,N__22536,N__29298,N__28555,N__25726,N__29520,N__27061,N__18853}),
            .WADDR({N__24364,N__26180,N__24678,N__25156,N__28098,N__28845,N__26823,N__26007,N__25546,N__27889,N__23986}),
            .MASK({dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829,dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,dangling_wire_841}),
            .WDATA({dangling_wire_842,dangling_wire_843,dangling_wire_844,dangling_wire_845,N__27269,dangling_wire_846,dangling_wire_847,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,N__23090,dangling_wire_853,dangling_wire_854,dangling_wire_855}),
            .RCLKE(),
            .RCLK(N__34626),
            .RE(N__19968),
            .WCLKE(N__28626),
            .WCLK(N__34627),
            .WE(N__19975));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_856,dangling_wire_857,dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_868,dangling_wire_869,dangling_wire_870,N__12195,N__11457,N__11190,N__11181,N__11499,N__12084,N__11469,N__11529}),
            .WADDR({dangling_wire_871,dangling_wire_872,dangling_wire_873,N__30855,N__20480,N__20561,N__20618,N__20264,N__29757,N__29836,N__29969}),
            .MASK({dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,dangling_wire_885,dangling_wire_886,dangling_wire_887,dangling_wire_888,dangling_wire_889}),
            .WDATA({dangling_wire_890,dangling_wire_891,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,dangling_wire_899,dangling_wire_900,dangling_wire_901,N__21138,N__22581,N__22713,N__20763}),
            .RCLKE(),
            .RCLK(N__34534),
            .RE(N__20098),
            .WCLKE(N__20736),
            .WCLK(N__34535),
            .WE(N__19964));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__35920),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__35922),
            .DIN(N__35921),
            .DOUT(N__35920),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__35922),
            .PADOUT(N__35921),
            .PADIN(N__35920),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__35911),
            .DIN(N__35910),
            .DOUT(N__35909),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__35911),
            .PADOUT(N__35910),
            .PADIN(N__35909),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__35902),
            .DIN(N__35901),
            .DOUT(N__35900),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__35902),
            .PADOUT(N__35901),
            .PADIN(N__35900),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__35893),
            .DIN(N__35892),
            .DOUT(N__35891),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__35893),
            .PADOUT(N__35892),
            .PADIN(N__35891),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12537),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__35884),
            .DIN(N__35883),
            .DOUT(N__35882),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__35884),
            .PADOUT(N__35883),
            .PADIN(N__35882),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12558),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__35875),
            .DIN(N__35874),
            .DOUT(N__35873),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__35875),
            .PADOUT(N__35874),
            .PADIN(N__35873),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__20041),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__35866),
            .DIN(N__35865),
            .DOUT(N__35864),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__35866),
            .PADOUT(N__35865),
            .PADIN(N__35864),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__17889),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__35857),
            .DIN(N__35856),
            .DOUT(N__35855),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__35857),
            .PADOUT(N__35856),
            .PADIN(N__35855),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__35848),
            .DIN(N__35847),
            .DOUT(N__35846),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__35848),
            .PADOUT(N__35847),
            .PADIN(N__35846),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__35839),
            .DIN(N__35838),
            .DOUT(N__35837),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__35839),
            .PADOUT(N__35838),
            .PADIN(N__35837),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__35830),
            .DIN(N__35829),
            .DOUT(N__35828),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__35830),
            .PADOUT(N__35829),
            .PADIN(N__35828),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__35821),
            .DIN(N__35820),
            .DOUT(N__35819),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__35821),
            .PADOUT(N__35820),
            .PADIN(N__35819),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__35812),
            .DIN(N__35811),
            .DOUT(N__35810),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__35812),
            .PADOUT(N__35811),
            .PADIN(N__35810),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__35803),
            .DIN(N__35802),
            .DOUT(N__35801),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__35803),
            .PADOUT(N__35802),
            .PADIN(N__35801),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__33282),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18556));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__35794),
            .DIN(N__35793),
            .DOUT(N__35792),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__35794),
            .PADOUT(N__35793),
            .PADIN(N__35792),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__33258),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18643));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__35785),
            .DIN(N__35784),
            .DOUT(N__35783),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__35785),
            .PADOUT(N__35784),
            .PADIN(N__35783),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__33231),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18626));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__35776),
            .DIN(N__35775),
            .DOUT(N__35774),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__35776),
            .PADOUT(N__35775),
            .PADIN(N__35774),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__33210),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18647));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__35767),
            .DIN(N__35766),
            .DOUT(N__35765),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__35767),
            .PADOUT(N__35766),
            .PADIN(N__35765),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__33186),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18613));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__35758),
            .DIN(N__35757),
            .DOUT(N__35756),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__35758),
            .PADOUT(N__35757),
            .PADIN(N__35756),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__33165),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18611));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__35749),
            .DIN(N__35748),
            .DOUT(N__35747),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__35749),
            .PADOUT(N__35748),
            .PADIN(N__35747),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__34251),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18609));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__35740),
            .DIN(N__35739),
            .DOUT(N__35738),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__35740),
            .PADOUT(N__35739),
            .PADIN(N__35738),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__34227),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18641));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__35731),
            .DIN(N__35730),
            .DOUT(N__35729),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__35731),
            .PADOUT(N__35730),
            .PADIN(N__35729),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__33786),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18597));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__35722),
            .DIN(N__35721),
            .DOUT(N__35720),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__35722),
            .PADOUT(N__35721),
            .PADIN(N__35720),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__33639),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18648));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__35713),
            .DIN(N__35712),
            .DOUT(N__35711),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__35713),
            .PADOUT(N__35712),
            .PADIN(N__35711),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__33492),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18636));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__35704),
            .DIN(N__35703),
            .DOUT(N__35702),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__35704),
            .PADOUT(N__35703),
            .PADIN(N__35702),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__33348),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18612));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__35695),
            .DIN(N__35694),
            .DOUT(N__35693),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__35695),
            .PADOUT(N__35694),
            .PADIN(N__35693),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35337),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18610));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__35686),
            .DIN(N__35685),
            .DOUT(N__35684),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__35686),
            .PADOUT(N__35685),
            .PADIN(N__35684),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35124),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18640));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__35677),
            .DIN(N__35676),
            .DOUT(N__35675),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__35677),
            .PADOUT(N__35676),
            .PADIN(N__35675),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__34083),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18596));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__35668),
            .DIN(N__35667),
            .DOUT(N__35666),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__35668),
            .PADOUT(N__35667),
            .PADIN(N__35666),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__33939),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18642));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__35659),
            .DIN(N__35658),
            .DOUT(N__35657),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__35659),
            .PADOUT(N__35658),
            .PADIN(N__35657),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__35650),
            .DIN(N__35649),
            .DOUT(N__35648),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__35650),
            .PADOUT(N__35649),
            .PADIN(N__35648),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__35641),
            .DIN(N__35640),
            .DOUT(N__35639),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__35641),
            .PADOUT(N__35640),
            .PADIN(N__35639),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__35632),
            .DIN(N__35631),
            .DOUT(N__35630),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__35632),
            .PADOUT(N__35631),
            .PADIN(N__35630),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__35623),
            .DIN(N__35622),
            .DOUT(N__35621),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__35623),
            .PADOUT(N__35622),
            .PADIN(N__35621),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__35614),
            .DIN(N__35613),
            .DOUT(N__35612),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__35614),
            .PADOUT(N__35613),
            .PADIN(N__35612),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__35605),
            .DIN(N__35604),
            .DOUT(N__35603),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__35605),
            .PADOUT(N__35604),
            .PADIN(N__35603),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__35596),
            .DIN(N__35595),
            .DOUT(N__35594),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__35596),
            .PADOUT(N__35595),
            .PADIN(N__35594),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__35587),
            .DIN(N__35586),
            .DOUT(N__35585),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__35587),
            .PADOUT(N__35586),
            .PADIN(N__35585),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__35578),
            .DIN(N__35577),
            .DOUT(N__35576),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__35578),
            .PADOUT(N__35577),
            .PADIN(N__35576),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10992),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__35569),
            .DIN(N__35568),
            .DOUT(N__35567),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__35569),
            .PADOUT(N__35568),
            .PADIN(N__35567),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21400),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__35560),
            .DIN(N__35559),
            .DOUT(N__35558),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__35560),
            .PADOUT(N__35559),
            .PADIN(N__35558),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__35551),
            .DIN(N__35550),
            .DOUT(N__35549),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__35551),
            .PADOUT(N__35550),
            .PADIN(N__35549),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10932),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__35542),
            .DIN(N__35541),
            .DOUT(N__35540),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__35542),
            .PADOUT(N__35541),
            .PADIN(N__35540),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__19729),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18590));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__35533),
            .DIN(N__35532),
            .DOUT(N__35531),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__35533),
            .PADOUT(N__35532),
            .PADIN(N__35531),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10977),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__35524),
            .DIN(N__35523),
            .DOUT(N__35522),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__35524),
            .PADOUT(N__35523),
            .PADIN(N__35522),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11124),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__35515),
            .DIN(N__35514),
            .DOUT(N__35513),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__35515),
            .PADOUT(N__35514),
            .PADIN(N__35513),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10962),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__35506),
            .DIN(N__35505),
            .DOUT(N__35504),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__35506),
            .PADOUT(N__35505),
            .PADIN(N__35504),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11172),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__35497),
            .DIN(N__35496),
            .DOUT(N__35495),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__35497),
            .PADOUT(N__35496),
            .PADIN(N__35495),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10950),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__35488),
            .DIN(N__35487),
            .DOUT(N__35486),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__35488),
            .PADOUT(N__35487),
            .PADIN(N__35486),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11145),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__35479),
            .DIN(N__35478),
            .DOUT(N__35477),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__35479),
            .PADOUT(N__35478),
            .PADIN(N__35477),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__35470),
            .DIN(N__35469),
            .DOUT(N__35468),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__35470),
            .PADOUT(N__35469),
            .PADIN(N__35468),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11154),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__35461),
            .DIN(N__35460),
            .DOUT(N__35459),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__35461),
            .PADOUT(N__35460),
            .PADIN(N__35459),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13956),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__8978 (
            .O(N__35442),
            .I(un1_M_this_external_address_q_cry_12));
    InMux I__8977 (
            .O(N__35439),
            .I(N__35434));
    InMux I__8976 (
            .O(N__35438),
            .I(N__35431));
    InMux I__8975 (
            .O(N__35437),
            .I(N__35428));
    LocalMux I__8974 (
            .O(N__35434),
            .I(N__35422));
    LocalMux I__8973 (
            .O(N__35431),
            .I(N__35417));
    LocalMux I__8972 (
            .O(N__35428),
            .I(N__35417));
    InMux I__8971 (
            .O(N__35427),
            .I(N__35414));
    InMux I__8970 (
            .O(N__35426),
            .I(N__35411));
    CascadeMux I__8969 (
            .O(N__35425),
            .I(N__35407));
    Span4Mux_v I__8968 (
            .O(N__35422),
            .I(N__35403));
    Span4Mux_v I__8967 (
            .O(N__35417),
            .I(N__35396));
    LocalMux I__8966 (
            .O(N__35414),
            .I(N__35396));
    LocalMux I__8965 (
            .O(N__35411),
            .I(N__35396));
    InMux I__8964 (
            .O(N__35410),
            .I(N__35393));
    InMux I__8963 (
            .O(N__35407),
            .I(N__35390));
    CascadeMux I__8962 (
            .O(N__35406),
            .I(N__35387));
    Sp12to4 I__8961 (
            .O(N__35403),
            .I(N__35384));
    Span4Mux_v I__8960 (
            .O(N__35396),
            .I(N__35380));
    LocalMux I__8959 (
            .O(N__35393),
            .I(N__35375));
    LocalMux I__8958 (
            .O(N__35390),
            .I(N__35375));
    InMux I__8957 (
            .O(N__35387),
            .I(N__35372));
    Span12Mux_h I__8956 (
            .O(N__35384),
            .I(N__35369));
    InMux I__8955 (
            .O(N__35383),
            .I(N__35366));
    Span4Mux_v I__8954 (
            .O(N__35380),
            .I(N__35359));
    Span4Mux_h I__8953 (
            .O(N__35375),
            .I(N__35359));
    LocalMux I__8952 (
            .O(N__35372),
            .I(N__35359));
    Span12Mux_v I__8951 (
            .O(N__35369),
            .I(N__35356));
    LocalMux I__8950 (
            .O(N__35366),
            .I(N__35353));
    Span4Mux_v I__8949 (
            .O(N__35359),
            .I(N__35350));
    Span12Mux_h I__8948 (
            .O(N__35356),
            .I(N__35345));
    Span12Mux_v I__8947 (
            .O(N__35353),
            .I(N__35345));
    Sp12to4 I__8946 (
            .O(N__35350),
            .I(N__35342));
    Odrv12 I__8945 (
            .O(N__35345),
            .I(port_data_c_6));
    Odrv12 I__8944 (
            .O(N__35342),
            .I(port_data_c_6));
    IoInMux I__8943 (
            .O(N__35337),
            .I(N__35334));
    LocalMux I__8942 (
            .O(N__35334),
            .I(N__35330));
    CascadeMux I__8941 (
            .O(N__35333),
            .I(N__35327));
    Span12Mux_s4_h I__8940 (
            .O(N__35330),
            .I(N__35324));
    InMux I__8939 (
            .O(N__35327),
            .I(N__35321));
    Odrv12 I__8938 (
            .O(N__35324),
            .I(M_this_external_address_qZ0Z_14));
    LocalMux I__8937 (
            .O(N__35321),
            .I(M_this_external_address_qZ0Z_14));
    InMux I__8936 (
            .O(N__35316),
            .I(un1_M_this_external_address_q_cry_13));
    InMux I__8935 (
            .O(N__35313),
            .I(N__35289));
    InMux I__8934 (
            .O(N__35312),
            .I(N__35289));
    InMux I__8933 (
            .O(N__35311),
            .I(N__35289));
    InMux I__8932 (
            .O(N__35310),
            .I(N__35289));
    InMux I__8931 (
            .O(N__35309),
            .I(N__35280));
    InMux I__8930 (
            .O(N__35308),
            .I(N__35280));
    InMux I__8929 (
            .O(N__35307),
            .I(N__35280));
    InMux I__8928 (
            .O(N__35306),
            .I(N__35280));
    InMux I__8927 (
            .O(N__35305),
            .I(N__35271));
    InMux I__8926 (
            .O(N__35304),
            .I(N__35271));
    InMux I__8925 (
            .O(N__35303),
            .I(N__35271));
    InMux I__8924 (
            .O(N__35302),
            .I(N__35271));
    InMux I__8923 (
            .O(N__35301),
            .I(N__35262));
    InMux I__8922 (
            .O(N__35300),
            .I(N__35262));
    InMux I__8921 (
            .O(N__35299),
            .I(N__35262));
    InMux I__8920 (
            .O(N__35298),
            .I(N__35262));
    LocalMux I__8919 (
            .O(N__35289),
            .I(N__35256));
    LocalMux I__8918 (
            .O(N__35280),
            .I(N__35256));
    LocalMux I__8917 (
            .O(N__35271),
            .I(N__35251));
    LocalMux I__8916 (
            .O(N__35262),
            .I(N__35251));
    InMux I__8915 (
            .O(N__35261),
            .I(N__35248));
    Span4Mux_v I__8914 (
            .O(N__35256),
            .I(N__35243));
    Span4Mux_v I__8913 (
            .O(N__35251),
            .I(N__35243));
    LocalMux I__8912 (
            .O(N__35248),
            .I(N__35240));
    Span4Mux_h I__8911 (
            .O(N__35243),
            .I(N__35237));
    Span4Mux_v I__8910 (
            .O(N__35240),
            .I(N__35234));
    Span4Mux_h I__8909 (
            .O(N__35237),
            .I(N__35231));
    Odrv4 I__8908 (
            .O(N__35234),
            .I(N_749_0));
    Odrv4 I__8907 (
            .O(N__35231),
            .I(N_749_0));
    InMux I__8906 (
            .O(N__35226),
            .I(N__35223));
    LocalMux I__8905 (
            .O(N__35223),
            .I(N__35218));
    InMux I__8904 (
            .O(N__35222),
            .I(N__35215));
    CascadeMux I__8903 (
            .O(N__35221),
            .I(N__35212));
    Span4Mux_v I__8902 (
            .O(N__35218),
            .I(N__35208));
    LocalMux I__8901 (
            .O(N__35215),
            .I(N__35205));
    InMux I__8900 (
            .O(N__35212),
            .I(N__35202));
    CascadeMux I__8899 (
            .O(N__35211),
            .I(N__35197));
    Span4Mux_h I__8898 (
            .O(N__35208),
            .I(N__35192));
    Span4Mux_v I__8897 (
            .O(N__35205),
            .I(N__35192));
    LocalMux I__8896 (
            .O(N__35202),
            .I(N__35189));
    CascadeMux I__8895 (
            .O(N__35201),
            .I(N__35186));
    InMux I__8894 (
            .O(N__35200),
            .I(N__35183));
    InMux I__8893 (
            .O(N__35197),
            .I(N__35180));
    Span4Mux_h I__8892 (
            .O(N__35192),
            .I(N__35175));
    Span4Mux_v I__8891 (
            .O(N__35189),
            .I(N__35175));
    InMux I__8890 (
            .O(N__35186),
            .I(N__35172));
    LocalMux I__8889 (
            .O(N__35183),
            .I(N__35169));
    LocalMux I__8888 (
            .O(N__35180),
            .I(N__35165));
    Sp12to4 I__8887 (
            .O(N__35175),
            .I(N__35160));
    LocalMux I__8886 (
            .O(N__35172),
            .I(N__35160));
    Span4Mux_v I__8885 (
            .O(N__35169),
            .I(N__35157));
    InMux I__8884 (
            .O(N__35168),
            .I(N__35154));
    Span4Mux_v I__8883 (
            .O(N__35165),
            .I(N__35151));
    Span12Mux_s6_h I__8882 (
            .O(N__35160),
            .I(N__35148));
    Sp12to4 I__8881 (
            .O(N__35157),
            .I(N__35143));
    LocalMux I__8880 (
            .O(N__35154),
            .I(N__35143));
    Span4Mux_v I__8879 (
            .O(N__35151),
            .I(N__35140));
    Span12Mux_v I__8878 (
            .O(N__35148),
            .I(N__35137));
    Span12Mux_v I__8877 (
            .O(N__35143),
            .I(N__35132));
    Sp12to4 I__8876 (
            .O(N__35140),
            .I(N__35132));
    Odrv12 I__8875 (
            .O(N__35137),
            .I(port_data_c_7));
    Odrv12 I__8874 (
            .O(N__35132),
            .I(port_data_c_7));
    InMux I__8873 (
            .O(N__35127),
            .I(un1_M_this_external_address_q_cry_14));
    IoInMux I__8872 (
            .O(N__35124),
            .I(N__35121));
    LocalMux I__8871 (
            .O(N__35121),
            .I(N__35118));
    Span4Mux_s0_h I__8870 (
            .O(N__35118),
            .I(N__35115));
    Span4Mux_h I__8869 (
            .O(N__35115),
            .I(N__35112));
    Sp12to4 I__8868 (
            .O(N__35112),
            .I(N__35109));
    Span12Mux_v I__8867 (
            .O(N__35109),
            .I(N__35105));
    InMux I__8866 (
            .O(N__35108),
            .I(N__35102));
    Odrv12 I__8865 (
            .O(N__35105),
            .I(M_this_external_address_qZ0Z_15));
    LocalMux I__8864 (
            .O(N__35102),
            .I(M_this_external_address_qZ0Z_15));
    InMux I__8863 (
            .O(N__35097),
            .I(N__35065));
    InMux I__8862 (
            .O(N__35096),
            .I(N__35065));
    InMux I__8861 (
            .O(N__35095),
            .I(N__35058));
    InMux I__8860 (
            .O(N__35094),
            .I(N__35058));
    InMux I__8859 (
            .O(N__35093),
            .I(N__35058));
    InMux I__8858 (
            .O(N__35092),
            .I(N__35055));
    InMux I__8857 (
            .O(N__35091),
            .I(N__35050));
    InMux I__8856 (
            .O(N__35090),
            .I(N__35050));
    InMux I__8855 (
            .O(N__35089),
            .I(N__35047));
    InMux I__8854 (
            .O(N__35088),
            .I(N__35044));
    InMux I__8853 (
            .O(N__35087),
            .I(N__35041));
    InMux I__8852 (
            .O(N__35086),
            .I(N__35038));
    InMux I__8851 (
            .O(N__35085),
            .I(N__35033));
    InMux I__8850 (
            .O(N__35084),
            .I(N__35033));
    InMux I__8849 (
            .O(N__35083),
            .I(N__35030));
    InMux I__8848 (
            .O(N__35082),
            .I(N__35027));
    InMux I__8847 (
            .O(N__35081),
            .I(N__35024));
    InMux I__8846 (
            .O(N__35080),
            .I(N__35019));
    InMux I__8845 (
            .O(N__35079),
            .I(N__35019));
    InMux I__8844 (
            .O(N__35078),
            .I(N__35014));
    InMux I__8843 (
            .O(N__35077),
            .I(N__35014));
    InMux I__8842 (
            .O(N__35076),
            .I(N__35011));
    InMux I__8841 (
            .O(N__35075),
            .I(N__35008));
    InMux I__8840 (
            .O(N__35074),
            .I(N__35001));
    InMux I__8839 (
            .O(N__35073),
            .I(N__35001));
    InMux I__8838 (
            .O(N__35072),
            .I(N__35001));
    InMux I__8837 (
            .O(N__35071),
            .I(N__34996));
    InMux I__8836 (
            .O(N__35070),
            .I(N__34996));
    LocalMux I__8835 (
            .O(N__35065),
            .I(N__34978));
    LocalMux I__8834 (
            .O(N__35058),
            .I(N__34975));
    LocalMux I__8833 (
            .O(N__35055),
            .I(N__34972));
    LocalMux I__8832 (
            .O(N__35050),
            .I(N__34969));
    LocalMux I__8831 (
            .O(N__35047),
            .I(N__34966));
    LocalMux I__8830 (
            .O(N__35044),
            .I(N__34963));
    LocalMux I__8829 (
            .O(N__35041),
            .I(N__34960));
    LocalMux I__8828 (
            .O(N__35038),
            .I(N__34957));
    LocalMux I__8827 (
            .O(N__35033),
            .I(N__34954));
    LocalMux I__8826 (
            .O(N__35030),
            .I(N__34951));
    LocalMux I__8825 (
            .O(N__35027),
            .I(N__34948));
    LocalMux I__8824 (
            .O(N__35024),
            .I(N__34945));
    LocalMux I__8823 (
            .O(N__35019),
            .I(N__34942));
    LocalMux I__8822 (
            .O(N__35014),
            .I(N__34939));
    LocalMux I__8821 (
            .O(N__35011),
            .I(N__34936));
    LocalMux I__8820 (
            .O(N__35008),
            .I(N__34933));
    LocalMux I__8819 (
            .O(N__35001),
            .I(N__34930));
    LocalMux I__8818 (
            .O(N__34996),
            .I(N__34927));
    SRMux I__8817 (
            .O(N__34995),
            .I(N__34860));
    SRMux I__8816 (
            .O(N__34994),
            .I(N__34860));
    SRMux I__8815 (
            .O(N__34993),
            .I(N__34860));
    SRMux I__8814 (
            .O(N__34992),
            .I(N__34860));
    SRMux I__8813 (
            .O(N__34991),
            .I(N__34860));
    SRMux I__8812 (
            .O(N__34990),
            .I(N__34860));
    SRMux I__8811 (
            .O(N__34989),
            .I(N__34860));
    SRMux I__8810 (
            .O(N__34988),
            .I(N__34860));
    SRMux I__8809 (
            .O(N__34987),
            .I(N__34860));
    SRMux I__8808 (
            .O(N__34986),
            .I(N__34860));
    SRMux I__8807 (
            .O(N__34985),
            .I(N__34860));
    SRMux I__8806 (
            .O(N__34984),
            .I(N__34860));
    SRMux I__8805 (
            .O(N__34983),
            .I(N__34860));
    SRMux I__8804 (
            .O(N__34982),
            .I(N__34860));
    SRMux I__8803 (
            .O(N__34981),
            .I(N__34860));
    Glb2LocalMux I__8802 (
            .O(N__34978),
            .I(N__34860));
    Glb2LocalMux I__8801 (
            .O(N__34975),
            .I(N__34860));
    Glb2LocalMux I__8800 (
            .O(N__34972),
            .I(N__34860));
    Glb2LocalMux I__8799 (
            .O(N__34969),
            .I(N__34860));
    Glb2LocalMux I__8798 (
            .O(N__34966),
            .I(N__34860));
    Glb2LocalMux I__8797 (
            .O(N__34963),
            .I(N__34860));
    Glb2LocalMux I__8796 (
            .O(N__34960),
            .I(N__34860));
    Glb2LocalMux I__8795 (
            .O(N__34957),
            .I(N__34860));
    Glb2LocalMux I__8794 (
            .O(N__34954),
            .I(N__34860));
    Glb2LocalMux I__8793 (
            .O(N__34951),
            .I(N__34860));
    Glb2LocalMux I__8792 (
            .O(N__34948),
            .I(N__34860));
    Glb2LocalMux I__8791 (
            .O(N__34945),
            .I(N__34860));
    Glb2LocalMux I__8790 (
            .O(N__34942),
            .I(N__34860));
    Glb2LocalMux I__8789 (
            .O(N__34939),
            .I(N__34860));
    Glb2LocalMux I__8788 (
            .O(N__34936),
            .I(N__34860));
    Glb2LocalMux I__8787 (
            .O(N__34933),
            .I(N__34860));
    Glb2LocalMux I__8786 (
            .O(N__34930),
            .I(N__34860));
    Glb2LocalMux I__8785 (
            .O(N__34927),
            .I(N__34860));
    GlobalMux I__8784 (
            .O(N__34860),
            .I(N__34857));
    gio2CtrlBuf I__8783 (
            .O(N__34857),
            .I(M_this_reset_cond_out_g_0));
    InMux I__8782 (
            .O(N__34854),
            .I(N__34851));
    LocalMux I__8781 (
            .O(N__34851),
            .I(N__34845));
    InMux I__8780 (
            .O(N__34850),
            .I(N__34838));
    InMux I__8779 (
            .O(N__34849),
            .I(N__34838));
    InMux I__8778 (
            .O(N__34848),
            .I(N__34838));
    Span4Mux_s3_h I__8777 (
            .O(N__34845),
            .I(N__34832));
    LocalMux I__8776 (
            .O(N__34838),
            .I(N__34832));
    InMux I__8775 (
            .O(N__34837),
            .I(N__34826));
    Span4Mux_h I__8774 (
            .O(N__34832),
            .I(N__34823));
    InMux I__8773 (
            .O(N__34831),
            .I(N__34820));
    InMux I__8772 (
            .O(N__34830),
            .I(N__34817));
    InMux I__8771 (
            .O(N__34829),
            .I(N__34813));
    LocalMux I__8770 (
            .O(N__34826),
            .I(N__34810));
    Span4Mux_h I__8769 (
            .O(N__34823),
            .I(N__34803));
    LocalMux I__8768 (
            .O(N__34820),
            .I(N__34803));
    LocalMux I__8767 (
            .O(N__34817),
            .I(N__34803));
    InMux I__8766 (
            .O(N__34816),
            .I(N__34800));
    LocalMux I__8765 (
            .O(N__34813),
            .I(N__34797));
    Span4Mux_h I__8764 (
            .O(N__34810),
            .I(N__34792));
    Span4Mux_h I__8763 (
            .O(N__34803),
            .I(N__34792));
    LocalMux I__8762 (
            .O(N__34800),
            .I(N__34789));
    Span4Mux_h I__8761 (
            .O(N__34797),
            .I(N__34786));
    Span4Mux_v I__8760 (
            .O(N__34792),
            .I(N__34781));
    Span4Mux_h I__8759 (
            .O(N__34789),
            .I(N__34781));
    Span4Mux_v I__8758 (
            .O(N__34786),
            .I(N__34777));
    Span4Mux_v I__8757 (
            .O(N__34781),
            .I(N__34774));
    InMux I__8756 (
            .O(N__34780),
            .I(N__34771));
    Span4Mux_v I__8755 (
            .O(N__34777),
            .I(N__34768));
    Span4Mux_v I__8754 (
            .O(N__34774),
            .I(N__34765));
    LocalMux I__8753 (
            .O(N__34771),
            .I(N__34762));
    Span4Mux_v I__8752 (
            .O(N__34768),
            .I(N__34759));
    Span4Mux_v I__8751 (
            .O(N__34765),
            .I(N__34756));
    Span12Mux_v I__8750 (
            .O(N__34762),
            .I(N__34753));
    Odrv4 I__8749 (
            .O(N__34759),
            .I(rst_n_c));
    Odrv4 I__8748 (
            .O(N__34756),
            .I(rst_n_c));
    Odrv12 I__8747 (
            .O(N__34753),
            .I(rst_n_c));
    InMux I__8746 (
            .O(N__34746),
            .I(N__34743));
    LocalMux I__8745 (
            .O(N__34743),
            .I(N__34740));
    Span4Mux_s2_h I__8744 (
            .O(N__34740),
            .I(N__34737));
    Odrv4 I__8743 (
            .O(N__34737),
            .I(\this_reset_cond.M_stage_qZ0Z_8 ));
    InMux I__8742 (
            .O(N__34734),
            .I(N__34730));
    InMux I__8741 (
            .O(N__34733),
            .I(N__34727));
    LocalMux I__8740 (
            .O(N__34730),
            .I(N__34716));
    LocalMux I__8739 (
            .O(N__34727),
            .I(N__34716));
    InMux I__8738 (
            .O(N__34726),
            .I(N__34705));
    InMux I__8737 (
            .O(N__34725),
            .I(N__34705));
    InMux I__8736 (
            .O(N__34724),
            .I(N__34705));
    InMux I__8735 (
            .O(N__34723),
            .I(N__34705));
    InMux I__8734 (
            .O(N__34722),
            .I(N__34705));
    InMux I__8733 (
            .O(N__34721),
            .I(N__34702));
    Span4Mux_h I__8732 (
            .O(N__34716),
            .I(N__34696));
    LocalMux I__8731 (
            .O(N__34705),
            .I(N__34696));
    LocalMux I__8730 (
            .O(N__34702),
            .I(N__34692));
    InMux I__8729 (
            .O(N__34701),
            .I(N__34689));
    Span4Mux_v I__8728 (
            .O(N__34696),
            .I(N__34686));
    InMux I__8727 (
            .O(N__34695),
            .I(N__34683));
    Span4Mux_h I__8726 (
            .O(N__34692),
            .I(N__34678));
    LocalMux I__8725 (
            .O(N__34689),
            .I(N__34678));
    Span4Mux_h I__8724 (
            .O(N__34686),
            .I(N__34675));
    LocalMux I__8723 (
            .O(N__34683),
            .I(N__34672));
    Sp12to4 I__8722 (
            .O(N__34678),
            .I(N__34669));
    Span4Mux_h I__8721 (
            .O(N__34675),
            .I(N__34664));
    Span4Mux_v I__8720 (
            .O(N__34672),
            .I(N__34664));
    Span12Mux_v I__8719 (
            .O(N__34669),
            .I(N__34661));
    Sp12to4 I__8718 (
            .O(N__34664),
            .I(N__34658));
    Span12Mux_h I__8717 (
            .O(N__34661),
            .I(N__34654));
    Span12Mux_h I__8716 (
            .O(N__34658),
            .I(N__34651));
    IoInMux I__8715 (
            .O(N__34657),
            .I(N__34648));
    Odrv12 I__8714 (
            .O(N__34654),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__8713 (
            .O(N__34651),
            .I(M_this_reset_cond_out_0));
    LocalMux I__8712 (
            .O(N__34648),
            .I(M_this_reset_cond_out_0));
    ClkMux I__8711 (
            .O(N__34641),
            .I(N__34257));
    ClkMux I__8710 (
            .O(N__34640),
            .I(N__34257));
    ClkMux I__8709 (
            .O(N__34639),
            .I(N__34257));
    ClkMux I__8708 (
            .O(N__34638),
            .I(N__34257));
    ClkMux I__8707 (
            .O(N__34637),
            .I(N__34257));
    ClkMux I__8706 (
            .O(N__34636),
            .I(N__34257));
    ClkMux I__8705 (
            .O(N__34635),
            .I(N__34257));
    ClkMux I__8704 (
            .O(N__34634),
            .I(N__34257));
    ClkMux I__8703 (
            .O(N__34633),
            .I(N__34257));
    ClkMux I__8702 (
            .O(N__34632),
            .I(N__34257));
    ClkMux I__8701 (
            .O(N__34631),
            .I(N__34257));
    ClkMux I__8700 (
            .O(N__34630),
            .I(N__34257));
    ClkMux I__8699 (
            .O(N__34629),
            .I(N__34257));
    ClkMux I__8698 (
            .O(N__34628),
            .I(N__34257));
    ClkMux I__8697 (
            .O(N__34627),
            .I(N__34257));
    ClkMux I__8696 (
            .O(N__34626),
            .I(N__34257));
    ClkMux I__8695 (
            .O(N__34625),
            .I(N__34257));
    ClkMux I__8694 (
            .O(N__34624),
            .I(N__34257));
    ClkMux I__8693 (
            .O(N__34623),
            .I(N__34257));
    ClkMux I__8692 (
            .O(N__34622),
            .I(N__34257));
    ClkMux I__8691 (
            .O(N__34621),
            .I(N__34257));
    ClkMux I__8690 (
            .O(N__34620),
            .I(N__34257));
    ClkMux I__8689 (
            .O(N__34619),
            .I(N__34257));
    ClkMux I__8688 (
            .O(N__34618),
            .I(N__34257));
    ClkMux I__8687 (
            .O(N__34617),
            .I(N__34257));
    ClkMux I__8686 (
            .O(N__34616),
            .I(N__34257));
    ClkMux I__8685 (
            .O(N__34615),
            .I(N__34257));
    ClkMux I__8684 (
            .O(N__34614),
            .I(N__34257));
    ClkMux I__8683 (
            .O(N__34613),
            .I(N__34257));
    ClkMux I__8682 (
            .O(N__34612),
            .I(N__34257));
    ClkMux I__8681 (
            .O(N__34611),
            .I(N__34257));
    ClkMux I__8680 (
            .O(N__34610),
            .I(N__34257));
    ClkMux I__8679 (
            .O(N__34609),
            .I(N__34257));
    ClkMux I__8678 (
            .O(N__34608),
            .I(N__34257));
    ClkMux I__8677 (
            .O(N__34607),
            .I(N__34257));
    ClkMux I__8676 (
            .O(N__34606),
            .I(N__34257));
    ClkMux I__8675 (
            .O(N__34605),
            .I(N__34257));
    ClkMux I__8674 (
            .O(N__34604),
            .I(N__34257));
    ClkMux I__8673 (
            .O(N__34603),
            .I(N__34257));
    ClkMux I__8672 (
            .O(N__34602),
            .I(N__34257));
    ClkMux I__8671 (
            .O(N__34601),
            .I(N__34257));
    ClkMux I__8670 (
            .O(N__34600),
            .I(N__34257));
    ClkMux I__8669 (
            .O(N__34599),
            .I(N__34257));
    ClkMux I__8668 (
            .O(N__34598),
            .I(N__34257));
    ClkMux I__8667 (
            .O(N__34597),
            .I(N__34257));
    ClkMux I__8666 (
            .O(N__34596),
            .I(N__34257));
    ClkMux I__8665 (
            .O(N__34595),
            .I(N__34257));
    ClkMux I__8664 (
            .O(N__34594),
            .I(N__34257));
    ClkMux I__8663 (
            .O(N__34593),
            .I(N__34257));
    ClkMux I__8662 (
            .O(N__34592),
            .I(N__34257));
    ClkMux I__8661 (
            .O(N__34591),
            .I(N__34257));
    ClkMux I__8660 (
            .O(N__34590),
            .I(N__34257));
    ClkMux I__8659 (
            .O(N__34589),
            .I(N__34257));
    ClkMux I__8658 (
            .O(N__34588),
            .I(N__34257));
    ClkMux I__8657 (
            .O(N__34587),
            .I(N__34257));
    ClkMux I__8656 (
            .O(N__34586),
            .I(N__34257));
    ClkMux I__8655 (
            .O(N__34585),
            .I(N__34257));
    ClkMux I__8654 (
            .O(N__34584),
            .I(N__34257));
    ClkMux I__8653 (
            .O(N__34583),
            .I(N__34257));
    ClkMux I__8652 (
            .O(N__34582),
            .I(N__34257));
    ClkMux I__8651 (
            .O(N__34581),
            .I(N__34257));
    ClkMux I__8650 (
            .O(N__34580),
            .I(N__34257));
    ClkMux I__8649 (
            .O(N__34579),
            .I(N__34257));
    ClkMux I__8648 (
            .O(N__34578),
            .I(N__34257));
    ClkMux I__8647 (
            .O(N__34577),
            .I(N__34257));
    ClkMux I__8646 (
            .O(N__34576),
            .I(N__34257));
    ClkMux I__8645 (
            .O(N__34575),
            .I(N__34257));
    ClkMux I__8644 (
            .O(N__34574),
            .I(N__34257));
    ClkMux I__8643 (
            .O(N__34573),
            .I(N__34257));
    ClkMux I__8642 (
            .O(N__34572),
            .I(N__34257));
    ClkMux I__8641 (
            .O(N__34571),
            .I(N__34257));
    ClkMux I__8640 (
            .O(N__34570),
            .I(N__34257));
    ClkMux I__8639 (
            .O(N__34569),
            .I(N__34257));
    ClkMux I__8638 (
            .O(N__34568),
            .I(N__34257));
    ClkMux I__8637 (
            .O(N__34567),
            .I(N__34257));
    ClkMux I__8636 (
            .O(N__34566),
            .I(N__34257));
    ClkMux I__8635 (
            .O(N__34565),
            .I(N__34257));
    ClkMux I__8634 (
            .O(N__34564),
            .I(N__34257));
    ClkMux I__8633 (
            .O(N__34563),
            .I(N__34257));
    ClkMux I__8632 (
            .O(N__34562),
            .I(N__34257));
    ClkMux I__8631 (
            .O(N__34561),
            .I(N__34257));
    ClkMux I__8630 (
            .O(N__34560),
            .I(N__34257));
    ClkMux I__8629 (
            .O(N__34559),
            .I(N__34257));
    ClkMux I__8628 (
            .O(N__34558),
            .I(N__34257));
    ClkMux I__8627 (
            .O(N__34557),
            .I(N__34257));
    ClkMux I__8626 (
            .O(N__34556),
            .I(N__34257));
    ClkMux I__8625 (
            .O(N__34555),
            .I(N__34257));
    ClkMux I__8624 (
            .O(N__34554),
            .I(N__34257));
    ClkMux I__8623 (
            .O(N__34553),
            .I(N__34257));
    ClkMux I__8622 (
            .O(N__34552),
            .I(N__34257));
    ClkMux I__8621 (
            .O(N__34551),
            .I(N__34257));
    ClkMux I__8620 (
            .O(N__34550),
            .I(N__34257));
    ClkMux I__8619 (
            .O(N__34549),
            .I(N__34257));
    ClkMux I__8618 (
            .O(N__34548),
            .I(N__34257));
    ClkMux I__8617 (
            .O(N__34547),
            .I(N__34257));
    ClkMux I__8616 (
            .O(N__34546),
            .I(N__34257));
    ClkMux I__8615 (
            .O(N__34545),
            .I(N__34257));
    ClkMux I__8614 (
            .O(N__34544),
            .I(N__34257));
    ClkMux I__8613 (
            .O(N__34543),
            .I(N__34257));
    ClkMux I__8612 (
            .O(N__34542),
            .I(N__34257));
    ClkMux I__8611 (
            .O(N__34541),
            .I(N__34257));
    ClkMux I__8610 (
            .O(N__34540),
            .I(N__34257));
    ClkMux I__8609 (
            .O(N__34539),
            .I(N__34257));
    ClkMux I__8608 (
            .O(N__34538),
            .I(N__34257));
    ClkMux I__8607 (
            .O(N__34537),
            .I(N__34257));
    ClkMux I__8606 (
            .O(N__34536),
            .I(N__34257));
    ClkMux I__8605 (
            .O(N__34535),
            .I(N__34257));
    ClkMux I__8604 (
            .O(N__34534),
            .I(N__34257));
    ClkMux I__8603 (
            .O(N__34533),
            .I(N__34257));
    ClkMux I__8602 (
            .O(N__34532),
            .I(N__34257));
    ClkMux I__8601 (
            .O(N__34531),
            .I(N__34257));
    ClkMux I__8600 (
            .O(N__34530),
            .I(N__34257));
    ClkMux I__8599 (
            .O(N__34529),
            .I(N__34257));
    ClkMux I__8598 (
            .O(N__34528),
            .I(N__34257));
    ClkMux I__8597 (
            .O(N__34527),
            .I(N__34257));
    ClkMux I__8596 (
            .O(N__34526),
            .I(N__34257));
    ClkMux I__8595 (
            .O(N__34525),
            .I(N__34257));
    ClkMux I__8594 (
            .O(N__34524),
            .I(N__34257));
    ClkMux I__8593 (
            .O(N__34523),
            .I(N__34257));
    ClkMux I__8592 (
            .O(N__34522),
            .I(N__34257));
    ClkMux I__8591 (
            .O(N__34521),
            .I(N__34257));
    ClkMux I__8590 (
            .O(N__34520),
            .I(N__34257));
    ClkMux I__8589 (
            .O(N__34519),
            .I(N__34257));
    ClkMux I__8588 (
            .O(N__34518),
            .I(N__34257));
    ClkMux I__8587 (
            .O(N__34517),
            .I(N__34257));
    ClkMux I__8586 (
            .O(N__34516),
            .I(N__34257));
    ClkMux I__8585 (
            .O(N__34515),
            .I(N__34257));
    ClkMux I__8584 (
            .O(N__34514),
            .I(N__34257));
    GlobalMux I__8583 (
            .O(N__34257),
            .I(N__34254));
    gio2CtrlBuf I__8582 (
            .O(N__34254),
            .I(clk_0_c_g));
    IoInMux I__8581 (
            .O(N__34251),
            .I(N__34248));
    LocalMux I__8580 (
            .O(N__34248),
            .I(N__34245));
    Span4Mux_s1_h I__8579 (
            .O(N__34245),
            .I(N__34242));
    Span4Mux_v I__8578 (
            .O(N__34242),
            .I(N__34238));
    InMux I__8577 (
            .O(N__34241),
            .I(N__34235));
    Odrv4 I__8576 (
            .O(N__34238),
            .I(M_this_external_address_qZ0Z_6));
    LocalMux I__8575 (
            .O(N__34235),
            .I(M_this_external_address_qZ0Z_6));
    InMux I__8574 (
            .O(N__34230),
            .I(un1_M_this_external_address_q_cry_5));
    IoInMux I__8573 (
            .O(N__34227),
            .I(N__34224));
    LocalMux I__8572 (
            .O(N__34224),
            .I(N__34221));
    Span4Mux_s0_h I__8571 (
            .O(N__34221),
            .I(N__34218));
    Span4Mux_h I__8570 (
            .O(N__34218),
            .I(N__34215));
    Sp12to4 I__8569 (
            .O(N__34215),
            .I(N__34212));
    Span12Mux_v I__8568 (
            .O(N__34212),
            .I(N__34208));
    InMux I__8567 (
            .O(N__34211),
            .I(N__34205));
    Odrv12 I__8566 (
            .O(N__34208),
            .I(M_this_external_address_qZ0Z_7));
    LocalMux I__8565 (
            .O(N__34205),
            .I(M_this_external_address_qZ0Z_7));
    InMux I__8564 (
            .O(N__34200),
            .I(un1_M_this_external_address_q_cry_6));
    CascadeMux I__8563 (
            .O(N__34197),
            .I(N__34194));
    InMux I__8562 (
            .O(N__34194),
            .I(N__34188));
    InMux I__8561 (
            .O(N__34193),
            .I(N__34185));
    InMux I__8560 (
            .O(N__34192),
            .I(N__34182));
    CascadeMux I__8559 (
            .O(N__34191),
            .I(N__34179));
    LocalMux I__8558 (
            .O(N__34188),
            .I(N__34174));
    LocalMux I__8557 (
            .O(N__34185),
            .I(N__34174));
    LocalMux I__8556 (
            .O(N__34182),
            .I(N__34170));
    InMux I__8555 (
            .O(N__34179),
            .I(N__34167));
    Span4Mux_h I__8554 (
            .O(N__34174),
            .I(N__34163));
    InMux I__8553 (
            .O(N__34173),
            .I(N__34160));
    Span4Mux_v I__8552 (
            .O(N__34170),
            .I(N__34155));
    LocalMux I__8551 (
            .O(N__34167),
            .I(N__34152));
    InMux I__8550 (
            .O(N__34166),
            .I(N__34149));
    Span4Mux_h I__8549 (
            .O(N__34163),
            .I(N__34144));
    LocalMux I__8548 (
            .O(N__34160),
            .I(N__34144));
    InMux I__8547 (
            .O(N__34159),
            .I(N__34141));
    InMux I__8546 (
            .O(N__34158),
            .I(N__34138));
    Span4Mux_h I__8545 (
            .O(N__34155),
            .I(N__34133));
    Span4Mux_v I__8544 (
            .O(N__34152),
            .I(N__34133));
    LocalMux I__8543 (
            .O(N__34149),
            .I(N__34130));
    Span4Mux_v I__8542 (
            .O(N__34144),
            .I(N__34127));
    LocalMux I__8541 (
            .O(N__34141),
            .I(N__34124));
    LocalMux I__8540 (
            .O(N__34138),
            .I(N__34120));
    Span4Mux_h I__8539 (
            .O(N__34133),
            .I(N__34117));
    Span4Mux_v I__8538 (
            .O(N__34130),
            .I(N__34110));
    Span4Mux_v I__8537 (
            .O(N__34127),
            .I(N__34110));
    Span4Mux_v I__8536 (
            .O(N__34124),
            .I(N__34110));
    InMux I__8535 (
            .O(N__34123),
            .I(N__34107));
    Span4Mux_v I__8534 (
            .O(N__34120),
            .I(N__34104));
    Sp12to4 I__8533 (
            .O(N__34117),
            .I(N__34097));
    Sp12to4 I__8532 (
            .O(N__34110),
            .I(N__34097));
    LocalMux I__8531 (
            .O(N__34107),
            .I(N__34097));
    Span4Mux_v I__8530 (
            .O(N__34104),
            .I(N__34094));
    Span12Mux_h I__8529 (
            .O(N__34097),
            .I(N__34091));
    Span4Mux_h I__8528 (
            .O(N__34094),
            .I(N__34088));
    Odrv12 I__8527 (
            .O(N__34091),
            .I(port_data_c_0));
    Odrv4 I__8526 (
            .O(N__34088),
            .I(port_data_c_0));
    IoInMux I__8525 (
            .O(N__34083),
            .I(N__34080));
    LocalMux I__8524 (
            .O(N__34080),
            .I(N__34077));
    Span4Mux_s2_v I__8523 (
            .O(N__34077),
            .I(N__34074));
    Sp12to4 I__8522 (
            .O(N__34074),
            .I(N__34071));
    Span12Mux_v I__8521 (
            .O(N__34071),
            .I(N__34067));
    CascadeMux I__8520 (
            .O(N__34070),
            .I(N__34064));
    Span12Mux_h I__8519 (
            .O(N__34067),
            .I(N__34061));
    InMux I__8518 (
            .O(N__34064),
            .I(N__34058));
    Odrv12 I__8517 (
            .O(N__34061),
            .I(M_this_external_address_qZ0Z_8));
    LocalMux I__8516 (
            .O(N__34058),
            .I(M_this_external_address_qZ0Z_8));
    InMux I__8515 (
            .O(N__34053),
            .I(bfn_28_22_0_));
    CascadeMux I__8514 (
            .O(N__34050),
            .I(N__34047));
    InMux I__8513 (
            .O(N__34047),
            .I(N__34043));
    InMux I__8512 (
            .O(N__34046),
            .I(N__34038));
    LocalMux I__8511 (
            .O(N__34043),
            .I(N__34033));
    InMux I__8510 (
            .O(N__34042),
            .I(N__34030));
    CascadeMux I__8509 (
            .O(N__34041),
            .I(N__34027));
    LocalMux I__8508 (
            .O(N__34038),
            .I(N__34024));
    InMux I__8507 (
            .O(N__34037),
            .I(N__34021));
    CascadeMux I__8506 (
            .O(N__34036),
            .I(N__34017));
    Span4Mux_v I__8505 (
            .O(N__34033),
            .I(N__34011));
    LocalMux I__8504 (
            .O(N__34030),
            .I(N__34011));
    InMux I__8503 (
            .O(N__34027),
            .I(N__34008));
    Span4Mux_v I__8502 (
            .O(N__34024),
            .I(N__34005));
    LocalMux I__8501 (
            .O(N__34021),
            .I(N__34002));
    InMux I__8500 (
            .O(N__34020),
            .I(N__33999));
    InMux I__8499 (
            .O(N__34017),
            .I(N__33996));
    InMux I__8498 (
            .O(N__34016),
            .I(N__33993));
    Span4Mux_v I__8497 (
            .O(N__34011),
            .I(N__33990));
    LocalMux I__8496 (
            .O(N__34008),
            .I(N__33987));
    Span4Mux_h I__8495 (
            .O(N__34005),
            .I(N__33980));
    Span4Mux_v I__8494 (
            .O(N__34002),
            .I(N__33980));
    LocalMux I__8493 (
            .O(N__33999),
            .I(N__33980));
    LocalMux I__8492 (
            .O(N__33996),
            .I(N__33974));
    LocalMux I__8491 (
            .O(N__33993),
            .I(N__33974));
    Span4Mux_v I__8490 (
            .O(N__33990),
            .I(N__33971));
    Span4Mux_v I__8489 (
            .O(N__33987),
            .I(N__33966));
    Span4Mux_v I__8488 (
            .O(N__33980),
            .I(N__33966));
    InMux I__8487 (
            .O(N__33979),
            .I(N__33963));
    Span12Mux_h I__8486 (
            .O(N__33974),
            .I(N__33960));
    Sp12to4 I__8485 (
            .O(N__33971),
            .I(N__33955));
    Sp12to4 I__8484 (
            .O(N__33966),
            .I(N__33955));
    LocalMux I__8483 (
            .O(N__33963),
            .I(N__33952));
    Span12Mux_v I__8482 (
            .O(N__33960),
            .I(N__33947));
    Span12Mux_h I__8481 (
            .O(N__33955),
            .I(N__33947));
    Sp12to4 I__8480 (
            .O(N__33952),
            .I(N__33944));
    Odrv12 I__8479 (
            .O(N__33947),
            .I(port_data_c_1));
    Odrv12 I__8478 (
            .O(N__33944),
            .I(port_data_c_1));
    IoInMux I__8477 (
            .O(N__33939),
            .I(N__33936));
    LocalMux I__8476 (
            .O(N__33936),
            .I(N__33933));
    IoSpan4Mux I__8475 (
            .O(N__33933),
            .I(N__33930));
    Span4Mux_s2_v I__8474 (
            .O(N__33930),
            .I(N__33926));
    CascadeMux I__8473 (
            .O(N__33929),
            .I(N__33923));
    Sp12to4 I__8472 (
            .O(N__33926),
            .I(N__33920));
    InMux I__8471 (
            .O(N__33923),
            .I(N__33917));
    Odrv12 I__8470 (
            .O(N__33920),
            .I(M_this_external_address_qZ0Z_9));
    LocalMux I__8469 (
            .O(N__33917),
            .I(M_this_external_address_qZ0Z_9));
    InMux I__8468 (
            .O(N__33912),
            .I(un1_M_this_external_address_q_cry_8));
    CascadeMux I__8467 (
            .O(N__33909),
            .I(N__33905));
    CascadeMux I__8466 (
            .O(N__33908),
            .I(N__33901));
    InMux I__8465 (
            .O(N__33905),
            .I(N__33898));
    InMux I__8464 (
            .O(N__33904),
            .I(N__33893));
    InMux I__8463 (
            .O(N__33901),
            .I(N__33889));
    LocalMux I__8462 (
            .O(N__33898),
            .I(N__33886));
    InMux I__8461 (
            .O(N__33897),
            .I(N__33883));
    CascadeMux I__8460 (
            .O(N__33896),
            .I(N__33880));
    LocalMux I__8459 (
            .O(N__33893),
            .I(N__33876));
    InMux I__8458 (
            .O(N__33892),
            .I(N__33873));
    LocalMux I__8457 (
            .O(N__33889),
            .I(N__33870));
    Span4Mux_v I__8456 (
            .O(N__33886),
            .I(N__33865));
    LocalMux I__8455 (
            .O(N__33883),
            .I(N__33865));
    InMux I__8454 (
            .O(N__33880),
            .I(N__33862));
    InMux I__8453 (
            .O(N__33879),
            .I(N__33859));
    Span4Mux_v I__8452 (
            .O(N__33876),
            .I(N__33854));
    LocalMux I__8451 (
            .O(N__33873),
            .I(N__33854));
    Span4Mux_h I__8450 (
            .O(N__33870),
            .I(N__33851));
    Span4Mux_v I__8449 (
            .O(N__33865),
            .I(N__33846));
    LocalMux I__8448 (
            .O(N__33862),
            .I(N__33846));
    LocalMux I__8447 (
            .O(N__33859),
            .I(N__33841));
    Span4Mux_v I__8446 (
            .O(N__33854),
            .I(N__33838));
    Span4Mux_h I__8445 (
            .O(N__33851),
            .I(N__33835));
    Span4Mux_v I__8444 (
            .O(N__33846),
            .I(N__33832));
    InMux I__8443 (
            .O(N__33845),
            .I(N__33829));
    InMux I__8442 (
            .O(N__33844),
            .I(N__33826));
    Span4Mux_v I__8441 (
            .O(N__33841),
            .I(N__33823));
    Sp12to4 I__8440 (
            .O(N__33838),
            .I(N__33820));
    Sp12to4 I__8439 (
            .O(N__33835),
            .I(N__33817));
    Span4Mux_h I__8438 (
            .O(N__33832),
            .I(N__33814));
    LocalMux I__8437 (
            .O(N__33829),
            .I(N__33809));
    LocalMux I__8436 (
            .O(N__33826),
            .I(N__33809));
    Span4Mux_v I__8435 (
            .O(N__33823),
            .I(N__33806));
    Span12Mux_h I__8434 (
            .O(N__33820),
            .I(N__33803));
    Span12Mux_v I__8433 (
            .O(N__33817),
            .I(N__33796));
    Sp12to4 I__8432 (
            .O(N__33814),
            .I(N__33796));
    Span12Mux_h I__8431 (
            .O(N__33809),
            .I(N__33796));
    IoSpan4Mux I__8430 (
            .O(N__33806),
            .I(N__33793));
    Odrv12 I__8429 (
            .O(N__33803),
            .I(port_data_c_2));
    Odrv12 I__8428 (
            .O(N__33796),
            .I(port_data_c_2));
    Odrv4 I__8427 (
            .O(N__33793),
            .I(port_data_c_2));
    IoInMux I__8426 (
            .O(N__33786),
            .I(N__33783));
    LocalMux I__8425 (
            .O(N__33783),
            .I(N__33780));
    Span4Mux_s3_v I__8424 (
            .O(N__33780),
            .I(N__33777));
    Span4Mux_h I__8423 (
            .O(N__33777),
            .I(N__33774));
    Span4Mux_h I__8422 (
            .O(N__33774),
            .I(N__33770));
    CascadeMux I__8421 (
            .O(N__33773),
            .I(N__33767));
    Span4Mux_v I__8420 (
            .O(N__33770),
            .I(N__33764));
    InMux I__8419 (
            .O(N__33767),
            .I(N__33761));
    Odrv4 I__8418 (
            .O(N__33764),
            .I(M_this_external_address_qZ0Z_10));
    LocalMux I__8417 (
            .O(N__33761),
            .I(M_this_external_address_qZ0Z_10));
    InMux I__8416 (
            .O(N__33756),
            .I(un1_M_this_external_address_q_cry_9));
    CascadeMux I__8415 (
            .O(N__33753),
            .I(N__33750));
    InMux I__8414 (
            .O(N__33750),
            .I(N__33746));
    CascadeMux I__8413 (
            .O(N__33749),
            .I(N__33743));
    LocalMux I__8412 (
            .O(N__33746),
            .I(N__33739));
    InMux I__8411 (
            .O(N__33743),
            .I(N__33736));
    InMux I__8410 (
            .O(N__33742),
            .I(N__33733));
    Span4Mux_v I__8409 (
            .O(N__33739),
            .I(N__33725));
    LocalMux I__8408 (
            .O(N__33736),
            .I(N__33725));
    LocalMux I__8407 (
            .O(N__33733),
            .I(N__33722));
    InMux I__8406 (
            .O(N__33732),
            .I(N__33719));
    InMux I__8405 (
            .O(N__33731),
            .I(N__33715));
    InMux I__8404 (
            .O(N__33730),
            .I(N__33712));
    Span4Mux_h I__8403 (
            .O(N__33725),
            .I(N__33705));
    Span4Mux_v I__8402 (
            .O(N__33722),
            .I(N__33705));
    LocalMux I__8401 (
            .O(N__33719),
            .I(N__33705));
    InMux I__8400 (
            .O(N__33718),
            .I(N__33702));
    LocalMux I__8399 (
            .O(N__33715),
            .I(N__33698));
    LocalMux I__8398 (
            .O(N__33712),
            .I(N__33694));
    Span4Mux_v I__8397 (
            .O(N__33705),
            .I(N__33691));
    LocalMux I__8396 (
            .O(N__33702),
            .I(N__33688));
    CascadeMux I__8395 (
            .O(N__33701),
            .I(N__33685));
    Span4Mux_h I__8394 (
            .O(N__33698),
            .I(N__33682));
    InMux I__8393 (
            .O(N__33697),
            .I(N__33679));
    Span4Mux_v I__8392 (
            .O(N__33694),
            .I(N__33676));
    Span4Mux_v I__8391 (
            .O(N__33691),
            .I(N__33673));
    Span4Mux_v I__8390 (
            .O(N__33688),
            .I(N__33670));
    InMux I__8389 (
            .O(N__33685),
            .I(N__33667));
    Span4Mux_h I__8388 (
            .O(N__33682),
            .I(N__33662));
    LocalMux I__8387 (
            .O(N__33679),
            .I(N__33662));
    Sp12to4 I__8386 (
            .O(N__33676),
            .I(N__33653));
    Sp12to4 I__8385 (
            .O(N__33673),
            .I(N__33653));
    Sp12to4 I__8384 (
            .O(N__33670),
            .I(N__33653));
    LocalMux I__8383 (
            .O(N__33667),
            .I(N__33653));
    Span4Mux_v I__8382 (
            .O(N__33662),
            .I(N__33650));
    Span12Mux_h I__8381 (
            .O(N__33653),
            .I(N__33647));
    Span4Mux_v I__8380 (
            .O(N__33650),
            .I(N__33644));
    Odrv12 I__8379 (
            .O(N__33647),
            .I(port_data_c_3));
    Odrv4 I__8378 (
            .O(N__33644),
            .I(port_data_c_3));
    IoInMux I__8377 (
            .O(N__33639),
            .I(N__33636));
    LocalMux I__8376 (
            .O(N__33636),
            .I(N__33633));
    IoSpan4Mux I__8375 (
            .O(N__33633),
            .I(N__33630));
    Span4Mux_s3_v I__8374 (
            .O(N__33630),
            .I(N__33626));
    CascadeMux I__8373 (
            .O(N__33629),
            .I(N__33623));
    Span4Mux_v I__8372 (
            .O(N__33626),
            .I(N__33620));
    InMux I__8371 (
            .O(N__33623),
            .I(N__33617));
    Odrv4 I__8370 (
            .O(N__33620),
            .I(M_this_external_address_qZ0Z_11));
    LocalMux I__8369 (
            .O(N__33617),
            .I(M_this_external_address_qZ0Z_11));
    InMux I__8368 (
            .O(N__33612),
            .I(un1_M_this_external_address_q_cry_10));
    CascadeMux I__8367 (
            .O(N__33609),
            .I(N__33601));
    InMux I__8366 (
            .O(N__33608),
            .I(N__33598));
    CascadeMux I__8365 (
            .O(N__33607),
            .I(N__33595));
    CascadeMux I__8364 (
            .O(N__33606),
            .I(N__33592));
    InMux I__8363 (
            .O(N__33605),
            .I(N__33589));
    InMux I__8362 (
            .O(N__33604),
            .I(N__33586));
    InMux I__8361 (
            .O(N__33601),
            .I(N__33581));
    LocalMux I__8360 (
            .O(N__33598),
            .I(N__33578));
    InMux I__8359 (
            .O(N__33595),
            .I(N__33575));
    InMux I__8358 (
            .O(N__33592),
            .I(N__33571));
    LocalMux I__8357 (
            .O(N__33589),
            .I(N__33568));
    LocalMux I__8356 (
            .O(N__33586),
            .I(N__33565));
    InMux I__8355 (
            .O(N__33585),
            .I(N__33562));
    InMux I__8354 (
            .O(N__33584),
            .I(N__33559));
    LocalMux I__8353 (
            .O(N__33581),
            .I(N__33556));
    Span4Mux_h I__8352 (
            .O(N__33578),
            .I(N__33553));
    LocalMux I__8351 (
            .O(N__33575),
            .I(N__33550));
    InMux I__8350 (
            .O(N__33574),
            .I(N__33547));
    LocalMux I__8349 (
            .O(N__33571),
            .I(N__33544));
    Span4Mux_v I__8348 (
            .O(N__33568),
            .I(N__33537));
    Span4Mux_h I__8347 (
            .O(N__33565),
            .I(N__33537));
    LocalMux I__8346 (
            .O(N__33562),
            .I(N__33537));
    LocalMux I__8345 (
            .O(N__33559),
            .I(N__33534));
    Span12Mux_h I__8344 (
            .O(N__33556),
            .I(N__33531));
    Sp12to4 I__8343 (
            .O(N__33553),
            .I(N__33526));
    Span12Mux_v I__8342 (
            .O(N__33550),
            .I(N__33526));
    LocalMux I__8341 (
            .O(N__33547),
            .I(N__33523));
    Span4Mux_v I__8340 (
            .O(N__33544),
            .I(N__33520));
    Span4Mux_v I__8339 (
            .O(N__33537),
            .I(N__33517));
    Span4Mux_v I__8338 (
            .O(N__33534),
            .I(N__33514));
    Span12Mux_v I__8337 (
            .O(N__33531),
            .I(N__33511));
    Span12Mux_v I__8336 (
            .O(N__33526),
            .I(N__33502));
    Span12Mux_h I__8335 (
            .O(N__33523),
            .I(N__33502));
    Sp12to4 I__8334 (
            .O(N__33520),
            .I(N__33502));
    Sp12to4 I__8333 (
            .O(N__33517),
            .I(N__33502));
    Span4Mux_v I__8332 (
            .O(N__33514),
            .I(N__33499));
    Odrv12 I__8331 (
            .O(N__33511),
            .I(port_data_c_4));
    Odrv12 I__8330 (
            .O(N__33502),
            .I(port_data_c_4));
    Odrv4 I__8329 (
            .O(N__33499),
            .I(port_data_c_4));
    IoInMux I__8328 (
            .O(N__33492),
            .I(N__33489));
    LocalMux I__8327 (
            .O(N__33489),
            .I(N__33485));
    CascadeMux I__8326 (
            .O(N__33488),
            .I(N__33482));
    Span4Mux_s3_h I__8325 (
            .O(N__33485),
            .I(N__33479));
    InMux I__8324 (
            .O(N__33482),
            .I(N__33476));
    Odrv4 I__8323 (
            .O(N__33479),
            .I(M_this_external_address_qZ0Z_12));
    LocalMux I__8322 (
            .O(N__33476),
            .I(M_this_external_address_qZ0Z_12));
    InMux I__8321 (
            .O(N__33471),
            .I(un1_M_this_external_address_q_cry_11));
    CascadeMux I__8320 (
            .O(N__33468),
            .I(N__33464));
    CascadeMux I__8319 (
            .O(N__33467),
            .I(N__33460));
    InMux I__8318 (
            .O(N__33464),
            .I(N__33454));
    InMux I__8317 (
            .O(N__33463),
            .I(N__33451));
    InMux I__8316 (
            .O(N__33460),
            .I(N__33448));
    InMux I__8315 (
            .O(N__33459),
            .I(N__33444));
    InMux I__8314 (
            .O(N__33458),
            .I(N__33441));
    CascadeMux I__8313 (
            .O(N__33457),
            .I(N__33438));
    LocalMux I__8312 (
            .O(N__33454),
            .I(N__33435));
    LocalMux I__8311 (
            .O(N__33451),
            .I(N__33432));
    LocalMux I__8310 (
            .O(N__33448),
            .I(N__33429));
    InMux I__8309 (
            .O(N__33447),
            .I(N__33426));
    LocalMux I__8308 (
            .O(N__33444),
            .I(N__33423));
    LocalMux I__8307 (
            .O(N__33441),
            .I(N__33420));
    InMux I__8306 (
            .O(N__33438),
            .I(N__33417));
    Span4Mux_v I__8305 (
            .O(N__33435),
            .I(N__33413));
    Span4Mux_h I__8304 (
            .O(N__33432),
            .I(N__33406));
    Span4Mux_v I__8303 (
            .O(N__33429),
            .I(N__33406));
    LocalMux I__8302 (
            .O(N__33426),
            .I(N__33406));
    Sp12to4 I__8301 (
            .O(N__33423),
            .I(N__33402));
    Span4Mux_v I__8300 (
            .O(N__33420),
            .I(N__33399));
    LocalMux I__8299 (
            .O(N__33417),
            .I(N__33396));
    InMux I__8298 (
            .O(N__33416),
            .I(N__33393));
    Span4Mux_v I__8297 (
            .O(N__33413),
            .I(N__33388));
    Span4Mux_v I__8296 (
            .O(N__33406),
            .I(N__33388));
    InMux I__8295 (
            .O(N__33405),
            .I(N__33385));
    Span12Mux_v I__8294 (
            .O(N__33402),
            .I(N__33382));
    Span4Mux_v I__8293 (
            .O(N__33399),
            .I(N__33377));
    Span4Mux_v I__8292 (
            .O(N__33396),
            .I(N__33377));
    LocalMux I__8291 (
            .O(N__33393),
            .I(N__33374));
    Span4Mux_h I__8290 (
            .O(N__33388),
            .I(N__33371));
    LocalMux I__8289 (
            .O(N__33385),
            .I(N__33368));
    Span12Mux_h I__8288 (
            .O(N__33382),
            .I(N__33361));
    Sp12to4 I__8287 (
            .O(N__33377),
            .I(N__33361));
    Span12Mux_v I__8286 (
            .O(N__33374),
            .I(N__33361));
    Span4Mux_h I__8285 (
            .O(N__33371),
            .I(N__33358));
    Span4Mux_v I__8284 (
            .O(N__33368),
            .I(N__33355));
    Odrv12 I__8283 (
            .O(N__33361),
            .I(port_data_c_5));
    Odrv4 I__8282 (
            .O(N__33358),
            .I(port_data_c_5));
    Odrv4 I__8281 (
            .O(N__33355),
            .I(port_data_c_5));
    IoInMux I__8280 (
            .O(N__33348),
            .I(N__33345));
    LocalMux I__8279 (
            .O(N__33345),
            .I(N__33341));
    CascadeMux I__8278 (
            .O(N__33344),
            .I(N__33338));
    Span4Mux_s3_h I__8277 (
            .O(N__33341),
            .I(N__33335));
    InMux I__8276 (
            .O(N__33338),
            .I(N__33332));
    Odrv4 I__8275 (
            .O(N__33335),
            .I(M_this_external_address_qZ0Z_13));
    LocalMux I__8274 (
            .O(N__33332),
            .I(M_this_external_address_qZ0Z_13));
    InMux I__8273 (
            .O(N__33327),
            .I(N__33324));
    LocalMux I__8272 (
            .O(N__33324),
            .I(N__33321));
    Odrv12 I__8271 (
            .O(N__33321),
            .I(\this_reset_cond.M_stage_qZ0Z_5 ));
    InMux I__8270 (
            .O(N__33318),
            .I(N__33315));
    LocalMux I__8269 (
            .O(N__33315),
            .I(\this_reset_cond.M_stage_qZ0Z_6 ));
    InMux I__8268 (
            .O(N__33312),
            .I(N__33309));
    LocalMux I__8267 (
            .O(N__33309),
            .I(\this_reset_cond.M_stage_qZ0Z_7 ));
    CascadeMux I__8266 (
            .O(N__33306),
            .I(N__33302));
    InMux I__8265 (
            .O(N__33305),
            .I(N__33299));
    InMux I__8264 (
            .O(N__33302),
            .I(N__33296));
    LocalMux I__8263 (
            .O(N__33299),
            .I(N__33291));
    LocalMux I__8262 (
            .O(N__33296),
            .I(N__33291));
    Span4Mux_h I__8261 (
            .O(N__33291),
            .I(N__33288));
    Span4Mux_h I__8260 (
            .O(N__33288),
            .I(N__33285));
    Odrv4 I__8259 (
            .O(N__33285),
            .I(un1_M_this_state_q_9_0_i));
    IoInMux I__8258 (
            .O(N__33282),
            .I(N__33279));
    LocalMux I__8257 (
            .O(N__33279),
            .I(N__33276));
    Span4Mux_s3_v I__8256 (
            .O(N__33276),
            .I(N__33273));
    Sp12to4 I__8255 (
            .O(N__33273),
            .I(N__33270));
    Span12Mux_h I__8254 (
            .O(N__33270),
            .I(N__33266));
    InMux I__8253 (
            .O(N__33269),
            .I(N__33263));
    Odrv12 I__8252 (
            .O(N__33266),
            .I(M_this_external_address_qZ0Z_0));
    LocalMux I__8251 (
            .O(N__33263),
            .I(M_this_external_address_qZ0Z_0));
    IoInMux I__8250 (
            .O(N__33258),
            .I(N__33255));
    LocalMux I__8249 (
            .O(N__33255),
            .I(N__33252));
    Span4Mux_s3_v I__8248 (
            .O(N__33252),
            .I(N__33249));
    Span4Mux_v I__8247 (
            .O(N__33249),
            .I(N__33246));
    Span4Mux_v I__8246 (
            .O(N__33246),
            .I(N__33242));
    InMux I__8245 (
            .O(N__33245),
            .I(N__33239));
    Odrv4 I__8244 (
            .O(N__33242),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__8243 (
            .O(N__33239),
            .I(M_this_external_address_qZ0Z_1));
    InMux I__8242 (
            .O(N__33234),
            .I(un1_M_this_external_address_q_cry_0));
    IoInMux I__8241 (
            .O(N__33231),
            .I(N__33228));
    LocalMux I__8240 (
            .O(N__33228),
            .I(N__33225));
    Span12Mux_s11_v I__8239 (
            .O(N__33225),
            .I(N__33221));
    InMux I__8238 (
            .O(N__33224),
            .I(N__33218));
    Odrv12 I__8237 (
            .O(N__33221),
            .I(M_this_external_address_qZ0Z_2));
    LocalMux I__8236 (
            .O(N__33218),
            .I(M_this_external_address_qZ0Z_2));
    InMux I__8235 (
            .O(N__33213),
            .I(un1_M_this_external_address_q_cry_1));
    IoInMux I__8234 (
            .O(N__33210),
            .I(N__33207));
    LocalMux I__8233 (
            .O(N__33207),
            .I(N__33204));
    Span4Mux_s3_h I__8232 (
            .O(N__33204),
            .I(N__33201));
    Span4Mux_v I__8231 (
            .O(N__33201),
            .I(N__33197));
    InMux I__8230 (
            .O(N__33200),
            .I(N__33194));
    Odrv4 I__8229 (
            .O(N__33197),
            .I(M_this_external_address_qZ0Z_3));
    LocalMux I__8228 (
            .O(N__33194),
            .I(M_this_external_address_qZ0Z_3));
    InMux I__8227 (
            .O(N__33189),
            .I(un1_M_this_external_address_q_cry_2));
    IoInMux I__8226 (
            .O(N__33186),
            .I(N__33183));
    LocalMux I__8225 (
            .O(N__33183),
            .I(N__33180));
    Span4Mux_s3_h I__8224 (
            .O(N__33180),
            .I(N__33176));
    InMux I__8223 (
            .O(N__33179),
            .I(N__33173));
    Odrv4 I__8222 (
            .O(N__33176),
            .I(M_this_external_address_qZ0Z_4));
    LocalMux I__8221 (
            .O(N__33173),
            .I(M_this_external_address_qZ0Z_4));
    InMux I__8220 (
            .O(N__33168),
            .I(un1_M_this_external_address_q_cry_3));
    IoInMux I__8219 (
            .O(N__33165),
            .I(N__33162));
    LocalMux I__8218 (
            .O(N__33162),
            .I(N__33158));
    InMux I__8217 (
            .O(N__33161),
            .I(N__33155));
    Odrv12 I__8216 (
            .O(N__33158),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__8215 (
            .O(N__33155),
            .I(M_this_external_address_qZ0Z_5));
    InMux I__8214 (
            .O(N__33150),
            .I(un1_M_this_external_address_q_cry_4));
    CascadeMux I__8213 (
            .O(N__33147),
            .I(N__33144));
    InMux I__8212 (
            .O(N__33144),
            .I(N__33141));
    LocalMux I__8211 (
            .O(N__33141),
            .I(N__33138));
    Span4Mux_h I__8210 (
            .O(N__33138),
            .I(N__33135));
    Odrv4 I__8209 (
            .O(N__33135),
            .I(M_this_data_tmp_qZ0Z_18));
    InMux I__8208 (
            .O(N__33132),
            .I(N__33129));
    LocalMux I__8207 (
            .O(N__33129),
            .I(N__33126));
    Odrv4 I__8206 (
            .O(N__33126),
            .I(M_this_oam_ram_write_data_18));
    CascadeMux I__8205 (
            .O(N__33123),
            .I(N__33120));
    InMux I__8204 (
            .O(N__33120),
            .I(N__33117));
    LocalMux I__8203 (
            .O(N__33117),
            .I(N__33114));
    Span4Mux_v I__8202 (
            .O(N__33114),
            .I(N__33111));
    Span4Mux_v I__8201 (
            .O(N__33111),
            .I(N__33108));
    Span4Mux_h I__8200 (
            .O(N__33108),
            .I(N__33105));
    Odrv4 I__8199 (
            .O(N__33105),
            .I(\this_ppu.un1_M_vaddress_q_3_5 ));
    InMux I__8198 (
            .O(N__33102),
            .I(N__33099));
    LocalMux I__8197 (
            .O(N__33099),
            .I(N__33096));
    Odrv4 I__8196 (
            .O(N__33096),
            .I(N_38_0));
    InMux I__8195 (
            .O(N__33093),
            .I(N__33090));
    LocalMux I__8194 (
            .O(N__33090),
            .I(M_this_oam_ram_write_data_31));
    InMux I__8193 (
            .O(N__33087),
            .I(N__33084));
    LocalMux I__8192 (
            .O(N__33084),
            .I(N_736_0));
    InMux I__8191 (
            .O(N__33081),
            .I(N__33078));
    LocalMux I__8190 (
            .O(N__33078),
            .I(N_737_0));
    InMux I__8189 (
            .O(N__33075),
            .I(N__33072));
    LocalMux I__8188 (
            .O(N__33072),
            .I(N__33068));
    InMux I__8187 (
            .O(N__33071),
            .I(N__33063));
    Span4Mux_v I__8186 (
            .O(N__33068),
            .I(N__33060));
    InMux I__8185 (
            .O(N__33067),
            .I(N__33057));
    InMux I__8184 (
            .O(N__33066),
            .I(N__33054));
    LocalMux I__8183 (
            .O(N__33063),
            .I(N__33047));
    Span4Mux_h I__8182 (
            .O(N__33060),
            .I(N__33047));
    LocalMux I__8181 (
            .O(N__33057),
            .I(N__33047));
    LocalMux I__8180 (
            .O(N__33054),
            .I(M_this_oam_ram_read_data_21));
    Odrv4 I__8179 (
            .O(N__33047),
            .I(M_this_oam_ram_read_data_21));
    InMux I__8178 (
            .O(N__33042),
            .I(N__33038));
    InMux I__8177 (
            .O(N__33041),
            .I(N__33035));
    LocalMux I__8176 (
            .O(N__33038),
            .I(N__33031));
    LocalMux I__8175 (
            .O(N__33035),
            .I(N__33026));
    InMux I__8174 (
            .O(N__33034),
            .I(N__33023));
    Span4Mux_v I__8173 (
            .O(N__33031),
            .I(N__33020));
    InMux I__8172 (
            .O(N__33030),
            .I(N__33017));
    InMux I__8171 (
            .O(N__33029),
            .I(N__33014));
    Span12Mux_h I__8170 (
            .O(N__33026),
            .I(N__33011));
    LocalMux I__8169 (
            .O(N__33023),
            .I(N__33004));
    Span4Mux_h I__8168 (
            .O(N__33020),
            .I(N__33004));
    LocalMux I__8167 (
            .O(N__33017),
            .I(N__33004));
    LocalMux I__8166 (
            .O(N__33014),
            .I(M_this_oam_ram_read_data_20));
    Odrv12 I__8165 (
            .O(N__33011),
            .I(M_this_oam_ram_read_data_20));
    Odrv4 I__8164 (
            .O(N__33004),
            .I(M_this_oam_ram_read_data_20));
    InMux I__8163 (
            .O(N__32997),
            .I(N__32992));
    InMux I__8162 (
            .O(N__32996),
            .I(N__32989));
    CascadeMux I__8161 (
            .O(N__32995),
            .I(N__32986));
    LocalMux I__8160 (
            .O(N__32992),
            .I(N__32983));
    LocalMux I__8159 (
            .O(N__32989),
            .I(N__32980));
    InMux I__8158 (
            .O(N__32986),
            .I(N__32977));
    Span12Mux_v I__8157 (
            .O(N__32983),
            .I(N__32974));
    Odrv4 I__8156 (
            .O(N__32980),
            .I(M_this_oam_ram_read_data_22));
    LocalMux I__8155 (
            .O(N__32977),
            .I(M_this_oam_ram_read_data_22));
    Odrv12 I__8154 (
            .O(N__32974),
            .I(M_this_oam_ram_read_data_22));
    InMux I__8153 (
            .O(N__32967),
            .I(N__32962));
    InMux I__8152 (
            .O(N__32966),
            .I(N__32959));
    InMux I__8151 (
            .O(N__32965),
            .I(N__32956));
    LocalMux I__8150 (
            .O(N__32962),
            .I(N__32953));
    LocalMux I__8149 (
            .O(N__32959),
            .I(N__32950));
    LocalMux I__8148 (
            .O(N__32956),
            .I(N__32944));
    Span4Mux_v I__8147 (
            .O(N__32953),
            .I(N__32944));
    Span4Mux_h I__8146 (
            .O(N__32950),
            .I(N__32939));
    InMux I__8145 (
            .O(N__32949),
            .I(N__32936));
    Span4Mux_v I__8144 (
            .O(N__32944),
            .I(N__32933));
    InMux I__8143 (
            .O(N__32943),
            .I(N__32930));
    InMux I__8142 (
            .O(N__32942),
            .I(N__32927));
    Span4Mux_h I__8141 (
            .O(N__32939),
            .I(N__32924));
    LocalMux I__8140 (
            .O(N__32936),
            .I(N__32917));
    Span4Mux_h I__8139 (
            .O(N__32933),
            .I(N__32917));
    LocalMux I__8138 (
            .O(N__32930),
            .I(N__32917));
    LocalMux I__8137 (
            .O(N__32927),
            .I(M_this_oam_ram_read_data_19));
    Odrv4 I__8136 (
            .O(N__32924),
            .I(M_this_oam_ram_read_data_19));
    Odrv4 I__8135 (
            .O(N__32917),
            .I(M_this_oam_ram_read_data_19));
    CascadeMux I__8134 (
            .O(N__32910),
            .I(N__32907));
    InMux I__8133 (
            .O(N__32907),
            .I(N__32904));
    LocalMux I__8132 (
            .O(N__32904),
            .I(N__32901));
    Span12Mux_h I__8131 (
            .O(N__32901),
            .I(N__32898));
    Odrv12 I__8130 (
            .O(N__32898),
            .I(\this_ppu.un1_M_vaddress_q_3_6 ));
    InMux I__8129 (
            .O(N__32895),
            .I(N__32887));
    InMux I__8128 (
            .O(N__32894),
            .I(N__32887));
    InMux I__8127 (
            .O(N__32893),
            .I(N__32882));
    InMux I__8126 (
            .O(N__32892),
            .I(N__32882));
    LocalMux I__8125 (
            .O(N__32887),
            .I(N__32871));
    LocalMux I__8124 (
            .O(N__32882),
            .I(N__32871));
    InMux I__8123 (
            .O(N__32881),
            .I(N__32866));
    InMux I__8122 (
            .O(N__32880),
            .I(N__32866));
    InMux I__8121 (
            .O(N__32879),
            .I(N__32837));
    InMux I__8120 (
            .O(N__32878),
            .I(N__32837));
    InMux I__8119 (
            .O(N__32877),
            .I(N__32832));
    InMux I__8118 (
            .O(N__32876),
            .I(N__32832));
    Span4Mux_v I__8117 (
            .O(N__32871),
            .I(N__32827));
    LocalMux I__8116 (
            .O(N__32866),
            .I(N__32827));
    InMux I__8115 (
            .O(N__32865),
            .I(N__32820));
    InMux I__8114 (
            .O(N__32864),
            .I(N__32820));
    InMux I__8113 (
            .O(N__32863),
            .I(N__32820));
    InMux I__8112 (
            .O(N__32862),
            .I(N__32817));
    InMux I__8111 (
            .O(N__32861),
            .I(N__32808));
    InMux I__8110 (
            .O(N__32860),
            .I(N__32808));
    InMux I__8109 (
            .O(N__32859),
            .I(N__32808));
    InMux I__8108 (
            .O(N__32858),
            .I(N__32808));
    InMux I__8107 (
            .O(N__32857),
            .I(N__32803));
    InMux I__8106 (
            .O(N__32856),
            .I(N__32803));
    InMux I__8105 (
            .O(N__32855),
            .I(N__32798));
    InMux I__8104 (
            .O(N__32854),
            .I(N__32798));
    InMux I__8103 (
            .O(N__32853),
            .I(N__32789));
    InMux I__8102 (
            .O(N__32852),
            .I(N__32789));
    InMux I__8101 (
            .O(N__32851),
            .I(N__32789));
    InMux I__8100 (
            .O(N__32850),
            .I(N__32789));
    InMux I__8099 (
            .O(N__32849),
            .I(N__32780));
    InMux I__8098 (
            .O(N__32848),
            .I(N__32780));
    InMux I__8097 (
            .O(N__32847),
            .I(N__32780));
    InMux I__8096 (
            .O(N__32846),
            .I(N__32780));
    InMux I__8095 (
            .O(N__32845),
            .I(N__32775));
    CascadeMux I__8094 (
            .O(N__32844),
            .I(N__32770));
    InMux I__8093 (
            .O(N__32843),
            .I(N__32766));
    InMux I__8092 (
            .O(N__32842),
            .I(N__32763));
    LocalMux I__8091 (
            .O(N__32837),
            .I(N__32754));
    LocalMux I__8090 (
            .O(N__32832),
            .I(N__32754));
    Span4Mux_h I__8089 (
            .O(N__32827),
            .I(N__32754));
    LocalMux I__8088 (
            .O(N__32820),
            .I(N__32754));
    LocalMux I__8087 (
            .O(N__32817),
            .I(N__32747));
    LocalMux I__8086 (
            .O(N__32808),
            .I(N__32747));
    LocalMux I__8085 (
            .O(N__32803),
            .I(N__32747));
    LocalMux I__8084 (
            .O(N__32798),
            .I(N__32744));
    LocalMux I__8083 (
            .O(N__32789),
            .I(N__32739));
    LocalMux I__8082 (
            .O(N__32780),
            .I(N__32739));
    InMux I__8081 (
            .O(N__32779),
            .I(N__32736));
    InMux I__8080 (
            .O(N__32778),
            .I(N__32733));
    LocalMux I__8079 (
            .O(N__32775),
            .I(N__32730));
    InMux I__8078 (
            .O(N__32774),
            .I(N__32721));
    InMux I__8077 (
            .O(N__32773),
            .I(N__32721));
    InMux I__8076 (
            .O(N__32770),
            .I(N__32721));
    InMux I__8075 (
            .O(N__32769),
            .I(N__32721));
    LocalMux I__8074 (
            .O(N__32766),
            .I(N__32710));
    LocalMux I__8073 (
            .O(N__32763),
            .I(N__32710));
    Span4Mux_v I__8072 (
            .O(N__32754),
            .I(N__32710));
    Span4Mux_v I__8071 (
            .O(N__32747),
            .I(N__32710));
    Span4Mux_v I__8070 (
            .O(N__32744),
            .I(N__32710));
    Span4Mux_h I__8069 (
            .O(N__32739),
            .I(N__32707));
    LocalMux I__8068 (
            .O(N__32736),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__8067 (
            .O(N__32733),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv12 I__8066 (
            .O(N__32730),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__8065 (
            .O(N__32721),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__8064 (
            .O(N__32710),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__8063 (
            .O(N__32707),
            .I(M_this_oam_address_qZ0Z_0));
    CascadeMux I__8062 (
            .O(N__32694),
            .I(N__32673));
    CascadeMux I__8061 (
            .O(N__32693),
            .I(N__32670));
    CascadeMux I__8060 (
            .O(N__32692),
            .I(N__32661));
    CascadeMux I__8059 (
            .O(N__32691),
            .I(N__32658));
    CascadeMux I__8058 (
            .O(N__32690),
            .I(N__32649));
    InMux I__8057 (
            .O(N__32689),
            .I(N__32646));
    InMux I__8056 (
            .O(N__32688),
            .I(N__32641));
    InMux I__8055 (
            .O(N__32687),
            .I(N__32641));
    InMux I__8054 (
            .O(N__32686),
            .I(N__32638));
    InMux I__8053 (
            .O(N__32685),
            .I(N__32633));
    InMux I__8052 (
            .O(N__32684),
            .I(N__32633));
    InMux I__8051 (
            .O(N__32683),
            .I(N__32628));
    InMux I__8050 (
            .O(N__32682),
            .I(N__32628));
    InMux I__8049 (
            .O(N__32681),
            .I(N__32623));
    InMux I__8048 (
            .O(N__32680),
            .I(N__32623));
    InMux I__8047 (
            .O(N__32679),
            .I(N__32618));
    InMux I__8046 (
            .O(N__32678),
            .I(N__32618));
    InMux I__8045 (
            .O(N__32677),
            .I(N__32613));
    InMux I__8044 (
            .O(N__32676),
            .I(N__32613));
    InMux I__8043 (
            .O(N__32673),
            .I(N__32606));
    InMux I__8042 (
            .O(N__32670),
            .I(N__32606));
    InMux I__8041 (
            .O(N__32669),
            .I(N__32606));
    InMux I__8040 (
            .O(N__32668),
            .I(N__32601));
    InMux I__8039 (
            .O(N__32667),
            .I(N__32601));
    InMux I__8038 (
            .O(N__32666),
            .I(N__32598));
    InMux I__8037 (
            .O(N__32665),
            .I(N__32591));
    InMux I__8036 (
            .O(N__32664),
            .I(N__32591));
    InMux I__8035 (
            .O(N__32661),
            .I(N__32591));
    InMux I__8034 (
            .O(N__32658),
            .I(N__32588));
    CascadeMux I__8033 (
            .O(N__32657),
            .I(N__32583));
    InMux I__8032 (
            .O(N__32656),
            .I(N__32575));
    InMux I__8031 (
            .O(N__32655),
            .I(N__32575));
    InMux I__8030 (
            .O(N__32654),
            .I(N__32575));
    InMux I__8029 (
            .O(N__32653),
            .I(N__32566));
    InMux I__8028 (
            .O(N__32652),
            .I(N__32566));
    InMux I__8027 (
            .O(N__32649),
            .I(N__32563));
    LocalMux I__8026 (
            .O(N__32646),
            .I(N__32560));
    LocalMux I__8025 (
            .O(N__32641),
            .I(N__32557));
    LocalMux I__8024 (
            .O(N__32638),
            .I(N__32538));
    LocalMux I__8023 (
            .O(N__32633),
            .I(N__32538));
    LocalMux I__8022 (
            .O(N__32628),
            .I(N__32538));
    LocalMux I__8021 (
            .O(N__32623),
            .I(N__32538));
    LocalMux I__8020 (
            .O(N__32618),
            .I(N__32538));
    LocalMux I__8019 (
            .O(N__32613),
            .I(N__32538));
    LocalMux I__8018 (
            .O(N__32606),
            .I(N__32538));
    LocalMux I__8017 (
            .O(N__32601),
            .I(N__32538));
    LocalMux I__8016 (
            .O(N__32598),
            .I(N__32538));
    LocalMux I__8015 (
            .O(N__32591),
            .I(N__32533));
    LocalMux I__8014 (
            .O(N__32588),
            .I(N__32533));
    InMux I__8013 (
            .O(N__32587),
            .I(N__32524));
    InMux I__8012 (
            .O(N__32586),
            .I(N__32524));
    InMux I__8011 (
            .O(N__32583),
            .I(N__32524));
    InMux I__8010 (
            .O(N__32582),
            .I(N__32524));
    LocalMux I__8009 (
            .O(N__32575),
            .I(N__32521));
    InMux I__8008 (
            .O(N__32574),
            .I(N__32516));
    InMux I__8007 (
            .O(N__32573),
            .I(N__32516));
    InMux I__8006 (
            .O(N__32572),
            .I(N__32513));
    InMux I__8005 (
            .O(N__32571),
            .I(N__32510));
    LocalMux I__8004 (
            .O(N__32566),
            .I(N__32507));
    LocalMux I__8003 (
            .O(N__32563),
            .I(N__32502));
    Span4Mux_v I__8002 (
            .O(N__32560),
            .I(N__32502));
    Span4Mux_v I__8001 (
            .O(N__32557),
            .I(N__32495));
    Span4Mux_v I__8000 (
            .O(N__32538),
            .I(N__32495));
    Span4Mux_v I__7999 (
            .O(N__32533),
            .I(N__32495));
    LocalMux I__7998 (
            .O(N__32524),
            .I(N__32490));
    Span4Mux_h I__7997 (
            .O(N__32521),
            .I(N__32490));
    LocalMux I__7996 (
            .O(N__32516),
            .I(M_this_oam_address_qZ0Z_1));
    LocalMux I__7995 (
            .O(N__32513),
            .I(M_this_oam_address_qZ0Z_1));
    LocalMux I__7994 (
            .O(N__32510),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv12 I__7993 (
            .O(N__32507),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__7992 (
            .O(N__32502),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__7991 (
            .O(N__32495),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__7990 (
            .O(N__32490),
            .I(M_this_oam_address_qZ0Z_1));
    CascadeMux I__7989 (
            .O(N__32475),
            .I(N__32472));
    InMux I__7988 (
            .O(N__32472),
            .I(N__32469));
    LocalMux I__7987 (
            .O(N__32469),
            .I(N__32466));
    Odrv4 I__7986 (
            .O(N__32466),
            .I(M_this_data_tmp_qZ0Z_21));
    InMux I__7985 (
            .O(N__32463),
            .I(N__32444));
    InMux I__7984 (
            .O(N__32462),
            .I(N__32444));
    InMux I__7983 (
            .O(N__32461),
            .I(N__32444));
    InMux I__7982 (
            .O(N__32460),
            .I(N__32444));
    InMux I__7981 (
            .O(N__32459),
            .I(N__32421));
    InMux I__7980 (
            .O(N__32458),
            .I(N__32421));
    InMux I__7979 (
            .O(N__32457),
            .I(N__32414));
    InMux I__7978 (
            .O(N__32456),
            .I(N__32414));
    InMux I__7977 (
            .O(N__32455),
            .I(N__32414));
    InMux I__7976 (
            .O(N__32454),
            .I(N__32409));
    InMux I__7975 (
            .O(N__32453),
            .I(N__32409));
    LocalMux I__7974 (
            .O(N__32444),
            .I(N__32406));
    InMux I__7973 (
            .O(N__32443),
            .I(N__32403));
    InMux I__7972 (
            .O(N__32442),
            .I(N__32394));
    InMux I__7971 (
            .O(N__32441),
            .I(N__32394));
    InMux I__7970 (
            .O(N__32440),
            .I(N__32394));
    InMux I__7969 (
            .O(N__32439),
            .I(N__32394));
    InMux I__7968 (
            .O(N__32438),
            .I(N__32385));
    InMux I__7967 (
            .O(N__32437),
            .I(N__32385));
    InMux I__7966 (
            .O(N__32436),
            .I(N__32385));
    InMux I__7965 (
            .O(N__32435),
            .I(N__32385));
    InMux I__7964 (
            .O(N__32434),
            .I(N__32378));
    InMux I__7963 (
            .O(N__32433),
            .I(N__32378));
    InMux I__7962 (
            .O(N__32432),
            .I(N__32368));
    InMux I__7961 (
            .O(N__32431),
            .I(N__32368));
    InMux I__7960 (
            .O(N__32430),
            .I(N__32359));
    InMux I__7959 (
            .O(N__32429),
            .I(N__32359));
    InMux I__7958 (
            .O(N__32428),
            .I(N__32359));
    InMux I__7957 (
            .O(N__32427),
            .I(N__32359));
    InMux I__7956 (
            .O(N__32426),
            .I(N__32356));
    LocalMux I__7955 (
            .O(N__32421),
            .I(N__32349));
    LocalMux I__7954 (
            .O(N__32414),
            .I(N__32349));
    LocalMux I__7953 (
            .O(N__32409),
            .I(N__32349));
    Span4Mux_h I__7952 (
            .O(N__32406),
            .I(N__32340));
    LocalMux I__7951 (
            .O(N__32403),
            .I(N__32340));
    LocalMux I__7950 (
            .O(N__32394),
            .I(N__32340));
    LocalMux I__7949 (
            .O(N__32385),
            .I(N__32340));
    CascadeMux I__7948 (
            .O(N__32384),
            .I(N__32337));
    InMux I__7947 (
            .O(N__32383),
            .I(N__32332));
    LocalMux I__7946 (
            .O(N__32378),
            .I(N__32329));
    InMux I__7945 (
            .O(N__32377),
            .I(N__32326));
    InMux I__7944 (
            .O(N__32376),
            .I(N__32323));
    InMux I__7943 (
            .O(N__32375),
            .I(N__32320));
    InMux I__7942 (
            .O(N__32374),
            .I(N__32315));
    InMux I__7941 (
            .O(N__32373),
            .I(N__32315));
    LocalMux I__7940 (
            .O(N__32368),
            .I(N__32310));
    LocalMux I__7939 (
            .O(N__32359),
            .I(N__32310));
    LocalMux I__7938 (
            .O(N__32356),
            .I(N__32303));
    Span4Mux_v I__7937 (
            .O(N__32349),
            .I(N__32303));
    Span4Mux_v I__7936 (
            .O(N__32340),
            .I(N__32303));
    InMux I__7935 (
            .O(N__32337),
            .I(N__32296));
    InMux I__7934 (
            .O(N__32336),
            .I(N__32296));
    InMux I__7933 (
            .O(N__32335),
            .I(N__32296));
    LocalMux I__7932 (
            .O(N__32332),
            .I(N__32287));
    Span4Mux_h I__7931 (
            .O(N__32329),
            .I(N__32287));
    LocalMux I__7930 (
            .O(N__32326),
            .I(N__32287));
    LocalMux I__7929 (
            .O(N__32323),
            .I(N__32287));
    LocalMux I__7928 (
            .O(N__32320),
            .I(N__32280));
    LocalMux I__7927 (
            .O(N__32315),
            .I(N__32280));
    Span4Mux_v I__7926 (
            .O(N__32310),
            .I(N__32280));
    Span4Mux_v I__7925 (
            .O(N__32303),
            .I(N__32277));
    LocalMux I__7924 (
            .O(N__32296),
            .I(N__32270));
    Span4Mux_v I__7923 (
            .O(N__32287),
            .I(N__32270));
    Span4Mux_h I__7922 (
            .O(N__32280),
            .I(N__32270));
    Odrv4 I__7921 (
            .O(N__32277),
            .I(N_122_0));
    Odrv4 I__7920 (
            .O(N__32270),
            .I(N_122_0));
    InMux I__7919 (
            .O(N__32265),
            .I(N__32262));
    LocalMux I__7918 (
            .O(N__32262),
            .I(M_this_oam_ram_write_data_21));
    InMux I__7917 (
            .O(N__32259),
            .I(N__32256));
    LocalMux I__7916 (
            .O(N__32256),
            .I(N__32252));
    InMux I__7915 (
            .O(N__32255),
            .I(N__32249));
    Span12Mux_s11_v I__7914 (
            .O(N__32252),
            .I(N__32246));
    LocalMux I__7913 (
            .O(N__32249),
            .I(N__32243));
    Span12Mux_v I__7912 (
            .O(N__32246),
            .I(N__32240));
    Span4Mux_h I__7911 (
            .O(N__32243),
            .I(N__32237));
    Odrv12 I__7910 (
            .O(N__32240),
            .I(M_this_oam_ram_read_data_6));
    Odrv4 I__7909 (
            .O(N__32237),
            .I(M_this_oam_ram_read_data_6));
    InMux I__7908 (
            .O(N__32232),
            .I(N__32229));
    LocalMux I__7907 (
            .O(N__32229),
            .I(N__32226));
    Span4Mux_h I__7906 (
            .O(N__32226),
            .I(N__32222));
    InMux I__7905 (
            .O(N__32225),
            .I(N__32219));
    Span4Mux_h I__7904 (
            .O(N__32222),
            .I(N__32214));
    LocalMux I__7903 (
            .O(N__32219),
            .I(N__32214));
    Odrv4 I__7902 (
            .O(N__32214),
            .I(M_this_oam_ram_read_data_5));
    InMux I__7901 (
            .O(N__32211),
            .I(N__32208));
    LocalMux I__7900 (
            .O(N__32208),
            .I(N__32205));
    Span4Mux_v I__7899 (
            .O(N__32205),
            .I(N__32202));
    Sp12to4 I__7898 (
            .O(N__32202),
            .I(N__32198));
    CascadeMux I__7897 (
            .O(N__32201),
            .I(N__32195));
    Span12Mux_h I__7896 (
            .O(N__32198),
            .I(N__32192));
    InMux I__7895 (
            .O(N__32195),
            .I(N__32189));
    Span12Mux_v I__7894 (
            .O(N__32192),
            .I(N__32186));
    LocalMux I__7893 (
            .O(N__32189),
            .I(N__32183));
    Odrv12 I__7892 (
            .O(N__32186),
            .I(M_this_oam_ram_read_data_7));
    Odrv4 I__7891 (
            .O(N__32183),
            .I(M_this_oam_ram_read_data_7));
    InMux I__7890 (
            .O(N__32178),
            .I(N__32175));
    LocalMux I__7889 (
            .O(N__32175),
            .I(N__32171));
    InMux I__7888 (
            .O(N__32174),
            .I(N__32168));
    Span4Mux_v I__7887 (
            .O(N__32171),
            .I(N__32165));
    LocalMux I__7886 (
            .O(N__32168),
            .I(N__32162));
    Odrv4 I__7885 (
            .O(N__32165),
            .I(M_this_oam_ram_read_data_4));
    Odrv4 I__7884 (
            .O(N__32162),
            .I(M_this_oam_ram_read_data_4));
    InMux I__7883 (
            .O(N__32157),
            .I(N__32154));
    LocalMux I__7882 (
            .O(N__32154),
            .I(N__32151));
    Span4Mux_h I__7881 (
            .O(N__32151),
            .I(N__32148));
    Span4Mux_h I__7880 (
            .O(N__32148),
            .I(N__32145));
    Odrv4 I__7879 (
            .O(N__32145),
            .I(\this_ppu.un9lto7Z0Z_4 ));
    CascadeMux I__7878 (
            .O(N__32142),
            .I(N__32139));
    InMux I__7877 (
            .O(N__32139),
            .I(N__32136));
    LocalMux I__7876 (
            .O(N__32136),
            .I(N__32133));
    Odrv4 I__7875 (
            .O(N__32133),
            .I(M_this_data_tmp_qZ0Z_9));
    InMux I__7874 (
            .O(N__32130),
            .I(N__32127));
    LocalMux I__7873 (
            .O(N__32127),
            .I(N_741_0));
    CascadeMux I__7872 (
            .O(N__32124),
            .I(N__32121));
    InMux I__7871 (
            .O(N__32121),
            .I(N__32118));
    LocalMux I__7870 (
            .O(N__32118),
            .I(N__32115));
    Span4Mux_v I__7869 (
            .O(N__32115),
            .I(N__32112));
    Span4Mux_h I__7868 (
            .O(N__32112),
            .I(N__32108));
    InMux I__7867 (
            .O(N__32111),
            .I(N__32105));
    Span4Mux_h I__7866 (
            .O(N__32108),
            .I(N__32100));
    LocalMux I__7865 (
            .O(N__32105),
            .I(N__32100));
    Odrv4 I__7864 (
            .O(N__32100),
            .I(M_this_oam_ram_read_data_23));
    CascadeMux I__7863 (
            .O(N__32097),
            .I(\this_ppu.un1_oam_data_c2_cascade_ ));
    InMux I__7862 (
            .O(N__32094),
            .I(N__32091));
    LocalMux I__7861 (
            .O(N__32091),
            .I(N__32088));
    Span4Mux_v I__7860 (
            .O(N__32088),
            .I(N__32085));
    Span4Mux_h I__7859 (
            .O(N__32085),
            .I(N__32082));
    Odrv4 I__7858 (
            .O(N__32082),
            .I(\this_ppu.un1_M_vaddress_q_3_7 ));
    CascadeMux I__7857 (
            .O(N__32079),
            .I(N__32076));
    InMux I__7856 (
            .O(N__32076),
            .I(N__32073));
    LocalMux I__7855 (
            .O(N__32073),
            .I(N__32070));
    Odrv4 I__7854 (
            .O(N__32070),
            .I(M_this_data_tmp_qZ0Z_13));
    InMux I__7853 (
            .O(N__32067),
            .I(N__32064));
    LocalMux I__7852 (
            .O(N__32064),
            .I(M_this_oam_ram_write_data_13));
    CascadeMux I__7851 (
            .O(N__32061),
            .I(N__32058));
    InMux I__7850 (
            .O(N__32058),
            .I(N__32055));
    LocalMux I__7849 (
            .O(N__32055),
            .I(N__32052));
    Span4Mux_v I__7848 (
            .O(N__32052),
            .I(N__32049));
    Span4Mux_h I__7847 (
            .O(N__32049),
            .I(N__32046));
    Odrv4 I__7846 (
            .O(N__32046),
            .I(M_this_data_tmp_qZ0Z_15));
    InMux I__7845 (
            .O(N__32043),
            .I(N__32040));
    LocalMux I__7844 (
            .O(N__32040),
            .I(M_this_oam_ram_write_data_15));
    CEMux I__7843 (
            .O(N__32037),
            .I(N__32034));
    LocalMux I__7842 (
            .O(N__32034),
            .I(N__32030));
    CEMux I__7841 (
            .O(N__32033),
            .I(N__32027));
    Span4Mux_v I__7840 (
            .O(N__32030),
            .I(N__32024));
    LocalMux I__7839 (
            .O(N__32027),
            .I(N__32021));
    Span4Mux_h I__7838 (
            .O(N__32024),
            .I(N__32018));
    Span4Mux_h I__7837 (
            .O(N__32021),
            .I(N__32015));
    Odrv4 I__7836 (
            .O(N__32018),
            .I(N_123_0));
    Odrv4 I__7835 (
            .O(N__32015),
            .I(N_123_0));
    InMux I__7834 (
            .O(N__32010),
            .I(N__32006));
    InMux I__7833 (
            .O(N__32009),
            .I(N__32003));
    LocalMux I__7832 (
            .O(N__32006),
            .I(N__32000));
    LocalMux I__7831 (
            .O(N__32003),
            .I(N__31997));
    Span12Mux_h I__7830 (
            .O(N__32000),
            .I(N__31994));
    Span4Mux_h I__7829 (
            .O(N__31997),
            .I(N__31991));
    Odrv12 I__7828 (
            .O(N__31994),
            .I(M_this_oam_ram_read_data_2));
    Odrv4 I__7827 (
            .O(N__31991),
            .I(M_this_oam_ram_read_data_2));
    CascadeMux I__7826 (
            .O(N__31986),
            .I(N__31983));
    InMux I__7825 (
            .O(N__31983),
            .I(N__31980));
    LocalMux I__7824 (
            .O(N__31980),
            .I(N__31977));
    Span4Mux_h I__7823 (
            .O(N__31977),
            .I(N__31974));
    Span4Mux_v I__7822 (
            .O(N__31974),
            .I(N__31970));
    InMux I__7821 (
            .O(N__31973),
            .I(N__31967));
    Span4Mux_h I__7820 (
            .O(N__31970),
            .I(N__31964));
    LocalMux I__7819 (
            .O(N__31967),
            .I(M_this_oam_ram_read_data_1));
    Odrv4 I__7818 (
            .O(N__31964),
            .I(M_this_oam_ram_read_data_1));
    InMux I__7817 (
            .O(N__31959),
            .I(N__31955));
    CascadeMux I__7816 (
            .O(N__31958),
            .I(N__31952));
    LocalMux I__7815 (
            .O(N__31955),
            .I(N__31949));
    InMux I__7814 (
            .O(N__31952),
            .I(N__31946));
    Odrv4 I__7813 (
            .O(N__31949),
            .I(M_this_oam_ram_read_data_3));
    LocalMux I__7812 (
            .O(N__31946),
            .I(M_this_oam_ram_read_data_3));
    InMux I__7811 (
            .O(N__31941),
            .I(N__31938));
    LocalMux I__7810 (
            .O(N__31938),
            .I(N__31935));
    Span4Mux_v I__7809 (
            .O(N__31935),
            .I(N__31932));
    Span4Mux_v I__7808 (
            .O(N__31932),
            .I(N__31929));
    Span4Mux_v I__7807 (
            .O(N__31929),
            .I(N__31926));
    Span4Mux_h I__7806 (
            .O(N__31926),
            .I(N__31922));
    InMux I__7805 (
            .O(N__31925),
            .I(N__31919));
    Odrv4 I__7804 (
            .O(N__31922),
            .I(M_this_oam_ram_read_data_0));
    LocalMux I__7803 (
            .O(N__31919),
            .I(M_this_oam_ram_read_data_0));
    InMux I__7802 (
            .O(N__31914),
            .I(N__31911));
    LocalMux I__7801 (
            .O(N__31911),
            .I(N__31908));
    Span4Mux_h I__7800 (
            .O(N__31908),
            .I(N__31905));
    Span4Mux_h I__7799 (
            .O(N__31905),
            .I(N__31902));
    Odrv4 I__7798 (
            .O(N__31902),
            .I(\this_ppu.un9lto7Z0Z_5 ));
    CascadeMux I__7797 (
            .O(N__31899),
            .I(N__31896));
    InMux I__7796 (
            .O(N__31896),
            .I(N__31892));
    CascadeMux I__7795 (
            .O(N__31895),
            .I(N__31889));
    LocalMux I__7794 (
            .O(N__31892),
            .I(N__31886));
    InMux I__7793 (
            .O(N__31889),
            .I(N__31883));
    Span4Mux_h I__7792 (
            .O(N__31886),
            .I(N__31880));
    LocalMux I__7791 (
            .O(N__31883),
            .I(N__31877));
    Span4Mux_v I__7790 (
            .O(N__31880),
            .I(N__31874));
    Span4Mux_h I__7789 (
            .O(N__31877),
            .I(N__31870));
    Span4Mux_v I__7788 (
            .O(N__31874),
            .I(N__31867));
    InMux I__7787 (
            .O(N__31873),
            .I(N__31864));
    Span4Mux_v I__7786 (
            .O(N__31870),
            .I(N__31861));
    Span4Mux_h I__7785 (
            .O(N__31867),
            .I(N__31858));
    LocalMux I__7784 (
            .O(N__31864),
            .I(N__31853));
    Span4Mux_h I__7783 (
            .O(N__31861),
            .I(N__31853));
    Odrv4 I__7782 (
            .O(N__31858),
            .I(M_this_oam_ram_read_data_17));
    Odrv4 I__7781 (
            .O(N__31853),
            .I(M_this_oam_ram_read_data_17));
    CascadeMux I__7780 (
            .O(N__31848),
            .I(N__31845));
    InMux I__7779 (
            .O(N__31845),
            .I(N__31842));
    LocalMux I__7778 (
            .O(N__31842),
            .I(N__31839));
    Odrv12 I__7777 (
            .O(N__31839),
            .I(M_this_oam_ram_read_data_i_17));
    CascadeMux I__7776 (
            .O(N__31836),
            .I(N__31832));
    InMux I__7775 (
            .O(N__31835),
            .I(N__31829));
    InMux I__7774 (
            .O(N__31832),
            .I(N__31826));
    LocalMux I__7773 (
            .O(N__31829),
            .I(N__31820));
    LocalMux I__7772 (
            .O(N__31826),
            .I(N__31820));
    InMux I__7771 (
            .O(N__31825),
            .I(N__31817));
    Span4Mux_h I__7770 (
            .O(N__31820),
            .I(N__31812));
    LocalMux I__7769 (
            .O(N__31817),
            .I(N__31812));
    Span4Mux_h I__7768 (
            .O(N__31812),
            .I(N__31809));
    Odrv4 I__7767 (
            .O(N__31809),
            .I(M_this_oam_ram_read_data_10));
    InMux I__7766 (
            .O(N__31806),
            .I(\this_ppu.un2_hscroll_cry_1 ));
    InMux I__7765 (
            .O(N__31803),
            .I(N__31800));
    LocalMux I__7764 (
            .O(N__31800),
            .I(N__31797));
    Odrv12 I__7763 (
            .O(N__31797),
            .I(\this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0 ));
    CascadeMux I__7762 (
            .O(N__31794),
            .I(N__31791));
    InMux I__7761 (
            .O(N__31791),
            .I(N__31786));
    CascadeMux I__7760 (
            .O(N__31790),
            .I(N__31783));
    InMux I__7759 (
            .O(N__31789),
            .I(N__31780));
    LocalMux I__7758 (
            .O(N__31786),
            .I(N__31777));
    InMux I__7757 (
            .O(N__31783),
            .I(N__31774));
    LocalMux I__7756 (
            .O(N__31780),
            .I(N__31771));
    Span4Mux_h I__7755 (
            .O(N__31777),
            .I(N__31766));
    LocalMux I__7754 (
            .O(N__31774),
            .I(N__31766));
    Span4Mux_h I__7753 (
            .O(N__31771),
            .I(N__31761));
    Span4Mux_h I__7752 (
            .O(N__31766),
            .I(N__31761));
    Span4Mux_v I__7751 (
            .O(N__31761),
            .I(N__31758));
    Odrv4 I__7750 (
            .O(N__31758),
            .I(M_this_oam_ram_read_data_9));
    CascadeMux I__7749 (
            .O(N__31755),
            .I(N__31752));
    InMux I__7748 (
            .O(N__31752),
            .I(N__31749));
    LocalMux I__7747 (
            .O(N__31749),
            .I(M_this_oam_ram_read_data_i_9));
    CascadeMux I__7746 (
            .O(N__31746),
            .I(N__31743));
    InMux I__7745 (
            .O(N__31743),
            .I(N__31740));
    LocalMux I__7744 (
            .O(N__31740),
            .I(N__31737));
    Odrv12 I__7743 (
            .O(N__31737),
            .I(M_this_data_tmp_qZ0Z_1));
    InMux I__7742 (
            .O(N__31734),
            .I(N__31731));
    LocalMux I__7741 (
            .O(N__31731),
            .I(N__31728));
    Span4Mux_v I__7740 (
            .O(N__31728),
            .I(N__31725));
    Odrv4 I__7739 (
            .O(N__31725),
            .I(N_747_0));
    CascadeMux I__7738 (
            .O(N__31722),
            .I(N__31719));
    InMux I__7737 (
            .O(N__31719),
            .I(N__31716));
    LocalMux I__7736 (
            .O(N__31716),
            .I(M_this_data_tmp_qZ0Z_10));
    InMux I__7735 (
            .O(N__31713),
            .I(N__31710));
    LocalMux I__7734 (
            .O(N__31710),
            .I(N__31707));
    Odrv4 I__7733 (
            .O(N__31707),
            .I(M_this_oam_ram_write_data_10));
    InMux I__7732 (
            .O(N__31704),
            .I(N__31701));
    LocalMux I__7731 (
            .O(N__31701),
            .I(N__31698));
    Span4Mux_h I__7730 (
            .O(N__31698),
            .I(N__31695));
    Span4Mux_h I__7729 (
            .O(N__31695),
            .I(N__31692));
    Span4Mux_h I__7728 (
            .O(N__31692),
            .I(N__31689));
    Span4Mux_h I__7727 (
            .O(N__31689),
            .I(N__31686));
    Odrv4 I__7726 (
            .O(N__31686),
            .I(M_this_map_ram_read_data_3));
    CascadeMux I__7725 (
            .O(N__31683),
            .I(N__31679));
    CascadeMux I__7724 (
            .O(N__31682),
            .I(N__31674));
    InMux I__7723 (
            .O(N__31679),
            .I(N__31668));
    CascadeMux I__7722 (
            .O(N__31678),
            .I(N__31664));
    CascadeMux I__7721 (
            .O(N__31677),
            .I(N__31660));
    InMux I__7720 (
            .O(N__31674),
            .I(N__31657));
    CascadeMux I__7719 (
            .O(N__31673),
            .I(N__31654));
    InMux I__7718 (
            .O(N__31672),
            .I(N__31649));
    InMux I__7717 (
            .O(N__31671),
            .I(N__31646));
    LocalMux I__7716 (
            .O(N__31668),
            .I(N__31643));
    CascadeMux I__7715 (
            .O(N__31667),
            .I(N__31639));
    InMux I__7714 (
            .O(N__31664),
            .I(N__31636));
    CascadeMux I__7713 (
            .O(N__31663),
            .I(N__31633));
    InMux I__7712 (
            .O(N__31660),
            .I(N__31630));
    LocalMux I__7711 (
            .O(N__31657),
            .I(N__31627));
    InMux I__7710 (
            .O(N__31654),
            .I(N__31624));
    CascadeMux I__7709 (
            .O(N__31653),
            .I(N__31621));
    CascadeMux I__7708 (
            .O(N__31652),
            .I(N__31618));
    LocalMux I__7707 (
            .O(N__31649),
            .I(N__31615));
    LocalMux I__7706 (
            .O(N__31646),
            .I(N__31612));
    Span4Mux_h I__7705 (
            .O(N__31643),
            .I(N__31609));
    InMux I__7704 (
            .O(N__31642),
            .I(N__31604));
    InMux I__7703 (
            .O(N__31639),
            .I(N__31604));
    LocalMux I__7702 (
            .O(N__31636),
            .I(N__31601));
    InMux I__7701 (
            .O(N__31633),
            .I(N__31598));
    LocalMux I__7700 (
            .O(N__31630),
            .I(N__31595));
    Span4Mux_h I__7699 (
            .O(N__31627),
            .I(N__31592));
    LocalMux I__7698 (
            .O(N__31624),
            .I(N__31589));
    InMux I__7697 (
            .O(N__31621),
            .I(N__31586));
    InMux I__7696 (
            .O(N__31618),
            .I(N__31583));
    Span4Mux_v I__7695 (
            .O(N__31615),
            .I(N__31579));
    Span4Mux_v I__7694 (
            .O(N__31612),
            .I(N__31571));
    Span4Mux_h I__7693 (
            .O(N__31609),
            .I(N__31571));
    LocalMux I__7692 (
            .O(N__31604),
            .I(N__31571));
    Span4Mux_h I__7691 (
            .O(N__31601),
            .I(N__31566));
    LocalMux I__7690 (
            .O(N__31598),
            .I(N__31566));
    Span4Mux_h I__7689 (
            .O(N__31595),
            .I(N__31563));
    Span4Mux_v I__7688 (
            .O(N__31592),
            .I(N__31556));
    Span4Mux_h I__7687 (
            .O(N__31589),
            .I(N__31556));
    LocalMux I__7686 (
            .O(N__31586),
            .I(N__31556));
    LocalMux I__7685 (
            .O(N__31583),
            .I(N__31553));
    InMux I__7684 (
            .O(N__31582),
            .I(N__31549));
    Span4Mux_v I__7683 (
            .O(N__31579),
            .I(N__31546));
    InMux I__7682 (
            .O(N__31578),
            .I(N__31543));
    Span4Mux_v I__7681 (
            .O(N__31571),
            .I(N__31536));
    Span4Mux_h I__7680 (
            .O(N__31566),
            .I(N__31536));
    Span4Mux_h I__7679 (
            .O(N__31563),
            .I(N__31536));
    Span4Mux_v I__7678 (
            .O(N__31556),
            .I(N__31531));
    Span4Mux_h I__7677 (
            .O(N__31553),
            .I(N__31531));
    InMux I__7676 (
            .O(N__31552),
            .I(N__31528));
    LocalMux I__7675 (
            .O(N__31549),
            .I(N__31525));
    Span4Mux_v I__7674 (
            .O(N__31546),
            .I(N__31520));
    LocalMux I__7673 (
            .O(N__31543),
            .I(N__31520));
    Span4Mux_v I__7672 (
            .O(N__31536),
            .I(N__31517));
    Span4Mux_h I__7671 (
            .O(N__31531),
            .I(N__31512));
    LocalMux I__7670 (
            .O(N__31528),
            .I(N__31512));
    Odrv4 I__7669 (
            .O(N__31525),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    Odrv4 I__7668 (
            .O(N__31520),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    Odrv4 I__7667 (
            .O(N__31517),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    Odrv4 I__7666 (
            .O(N__31512),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    CascadeMux I__7665 (
            .O(N__31503),
            .I(N__31496));
    InMux I__7664 (
            .O(N__31502),
            .I(N__31493));
    InMux I__7663 (
            .O(N__31501),
            .I(N__31489));
    InMux I__7662 (
            .O(N__31500),
            .I(N__31486));
    InMux I__7661 (
            .O(N__31499),
            .I(N__31483));
    InMux I__7660 (
            .O(N__31496),
            .I(N__31474));
    LocalMux I__7659 (
            .O(N__31493),
            .I(N__31471));
    InMux I__7658 (
            .O(N__31492),
            .I(N__31468));
    LocalMux I__7657 (
            .O(N__31489),
            .I(N__31465));
    LocalMux I__7656 (
            .O(N__31486),
            .I(N__31461));
    LocalMux I__7655 (
            .O(N__31483),
            .I(N__31458));
    InMux I__7654 (
            .O(N__31482),
            .I(N__31454));
    InMux I__7653 (
            .O(N__31481),
            .I(N__31449));
    InMux I__7652 (
            .O(N__31480),
            .I(N__31446));
    InMux I__7651 (
            .O(N__31479),
            .I(N__31441));
    InMux I__7650 (
            .O(N__31478),
            .I(N__31441));
    InMux I__7649 (
            .O(N__31477),
            .I(N__31438));
    LocalMux I__7648 (
            .O(N__31474),
            .I(N__31434));
    Span4Mux_h I__7647 (
            .O(N__31471),
            .I(N__31429));
    LocalMux I__7646 (
            .O(N__31468),
            .I(N__31429));
    Span4Mux_v I__7645 (
            .O(N__31465),
            .I(N__31426));
    InMux I__7644 (
            .O(N__31464),
            .I(N__31423));
    Span4Mux_h I__7643 (
            .O(N__31461),
            .I(N__31418));
    Span4Mux_h I__7642 (
            .O(N__31458),
            .I(N__31418));
    InMux I__7641 (
            .O(N__31457),
            .I(N__31415));
    LocalMux I__7640 (
            .O(N__31454),
            .I(N__31412));
    InMux I__7639 (
            .O(N__31453),
            .I(N__31407));
    InMux I__7638 (
            .O(N__31452),
            .I(N__31407));
    LocalMux I__7637 (
            .O(N__31449),
            .I(N__31404));
    LocalMux I__7636 (
            .O(N__31446),
            .I(N__31399));
    LocalMux I__7635 (
            .O(N__31441),
            .I(N__31399));
    LocalMux I__7634 (
            .O(N__31438),
            .I(N__31396));
    InMux I__7633 (
            .O(N__31437),
            .I(N__31393));
    Span4Mux_h I__7632 (
            .O(N__31434),
            .I(N__31388));
    Span4Mux_h I__7631 (
            .O(N__31429),
            .I(N__31388));
    Sp12to4 I__7630 (
            .O(N__31426),
            .I(N__31383));
    LocalMux I__7629 (
            .O(N__31423),
            .I(N__31383));
    Sp12to4 I__7628 (
            .O(N__31418),
            .I(N__31378));
    LocalMux I__7627 (
            .O(N__31415),
            .I(N__31378));
    Span4Mux_h I__7626 (
            .O(N__31412),
            .I(N__31375));
    LocalMux I__7625 (
            .O(N__31407),
            .I(N__31372));
    Span4Mux_v I__7624 (
            .O(N__31404),
            .I(N__31367));
    Span4Mux_v I__7623 (
            .O(N__31399),
            .I(N__31367));
    Span4Mux_h I__7622 (
            .O(N__31396),
            .I(N__31364));
    LocalMux I__7621 (
            .O(N__31393),
            .I(N__31361));
    Sp12to4 I__7620 (
            .O(N__31388),
            .I(N__31356));
    Span12Mux_h I__7619 (
            .O(N__31383),
            .I(N__31356));
    Span12Mux_v I__7618 (
            .O(N__31378),
            .I(N__31353));
    Span4Mux_h I__7617 (
            .O(N__31375),
            .I(N__31346));
    Span4Mux_h I__7616 (
            .O(N__31372),
            .I(N__31346));
    Span4Mux_v I__7615 (
            .O(N__31367),
            .I(N__31346));
    Odrv4 I__7614 (
            .O(N__31364),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv12 I__7613 (
            .O(N__31361),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv12 I__7612 (
            .O(N__31356),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv12 I__7611 (
            .O(N__31353),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__7610 (
            .O(N__31346),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    CascadeMux I__7609 (
            .O(N__31335),
            .I(N__31331));
    CascadeMux I__7608 (
            .O(N__31334),
            .I(N__31326));
    InMux I__7607 (
            .O(N__31331),
            .I(N__31322));
    CascadeMux I__7606 (
            .O(N__31330),
            .I(N__31319));
    CascadeMux I__7605 (
            .O(N__31329),
            .I(N__31316));
    InMux I__7604 (
            .O(N__31326),
            .I(N__31311));
    CascadeMux I__7603 (
            .O(N__31325),
            .I(N__31308));
    LocalMux I__7602 (
            .O(N__31322),
            .I(N__31304));
    InMux I__7601 (
            .O(N__31319),
            .I(N__31301));
    InMux I__7600 (
            .O(N__31316),
            .I(N__31298));
    CascadeMux I__7599 (
            .O(N__31315),
            .I(N__31295));
    CascadeMux I__7598 (
            .O(N__31314),
            .I(N__31292));
    LocalMux I__7597 (
            .O(N__31311),
            .I(N__31288));
    InMux I__7596 (
            .O(N__31308),
            .I(N__31285));
    CascadeMux I__7595 (
            .O(N__31307),
            .I(N__31282));
    Span4Mux_h I__7594 (
            .O(N__31304),
            .I(N__31278));
    LocalMux I__7593 (
            .O(N__31301),
            .I(N__31275));
    LocalMux I__7592 (
            .O(N__31298),
            .I(N__31272));
    InMux I__7591 (
            .O(N__31295),
            .I(N__31269));
    InMux I__7590 (
            .O(N__31292),
            .I(N__31266));
    CascadeMux I__7589 (
            .O(N__31291),
            .I(N__31263));
    Span4Mux_h I__7588 (
            .O(N__31288),
            .I(N__31258));
    LocalMux I__7587 (
            .O(N__31285),
            .I(N__31255));
    InMux I__7586 (
            .O(N__31282),
            .I(N__31252));
    CascadeMux I__7585 (
            .O(N__31281),
            .I(N__31249));
    Span4Mux_v I__7584 (
            .O(N__31278),
            .I(N__31243));
    Span4Mux_h I__7583 (
            .O(N__31275),
            .I(N__31243));
    Span4Mux_v I__7582 (
            .O(N__31272),
            .I(N__31240));
    LocalMux I__7581 (
            .O(N__31269),
            .I(N__31237));
    LocalMux I__7580 (
            .O(N__31266),
            .I(N__31234));
    InMux I__7579 (
            .O(N__31263),
            .I(N__31231));
    CascadeMux I__7578 (
            .O(N__31262),
            .I(N__31228));
    CascadeMux I__7577 (
            .O(N__31261),
            .I(N__31224));
    Span4Mux_v I__7576 (
            .O(N__31258),
            .I(N__31219));
    Span4Mux_h I__7575 (
            .O(N__31255),
            .I(N__31219));
    LocalMux I__7574 (
            .O(N__31252),
            .I(N__31216));
    InMux I__7573 (
            .O(N__31249),
            .I(N__31213));
    CascadeMux I__7572 (
            .O(N__31248),
            .I(N__31210));
    Span4Mux_v I__7571 (
            .O(N__31243),
            .I(N__31203));
    Span4Mux_h I__7570 (
            .O(N__31240),
            .I(N__31203));
    Span4Mux_h I__7569 (
            .O(N__31237),
            .I(N__31203));
    Span4Mux_h I__7568 (
            .O(N__31234),
            .I(N__31200));
    LocalMux I__7567 (
            .O(N__31231),
            .I(N__31197));
    InMux I__7566 (
            .O(N__31228),
            .I(N__31194));
    CascadeMux I__7565 (
            .O(N__31227),
            .I(N__31191));
    InMux I__7564 (
            .O(N__31224),
            .I(N__31187));
    Span4Mux_v I__7563 (
            .O(N__31219),
            .I(N__31182));
    Span4Mux_h I__7562 (
            .O(N__31216),
            .I(N__31182));
    LocalMux I__7561 (
            .O(N__31213),
            .I(N__31179));
    InMux I__7560 (
            .O(N__31210),
            .I(N__31176));
    Span4Mux_h I__7559 (
            .O(N__31203),
            .I(N__31173));
    Span4Mux_v I__7558 (
            .O(N__31200),
            .I(N__31168));
    Span4Mux_h I__7557 (
            .O(N__31197),
            .I(N__31168));
    LocalMux I__7556 (
            .O(N__31194),
            .I(N__31165));
    InMux I__7555 (
            .O(N__31191),
            .I(N__31162));
    CascadeMux I__7554 (
            .O(N__31190),
            .I(N__31159));
    LocalMux I__7553 (
            .O(N__31187),
            .I(N__31156));
    Span4Mux_v I__7552 (
            .O(N__31182),
            .I(N__31151));
    Span4Mux_h I__7551 (
            .O(N__31179),
            .I(N__31151));
    LocalMux I__7550 (
            .O(N__31176),
            .I(N__31148));
    Span4Mux_h I__7549 (
            .O(N__31173),
            .I(N__31145));
    Span4Mux_v I__7548 (
            .O(N__31168),
            .I(N__31140));
    Span4Mux_h I__7547 (
            .O(N__31165),
            .I(N__31140));
    LocalMux I__7546 (
            .O(N__31162),
            .I(N__31137));
    InMux I__7545 (
            .O(N__31159),
            .I(N__31134));
    Span12Mux_h I__7544 (
            .O(N__31156),
            .I(N__31130));
    Span4Mux_v I__7543 (
            .O(N__31151),
            .I(N__31125));
    Span4Mux_h I__7542 (
            .O(N__31148),
            .I(N__31125));
    Span4Mux_h I__7541 (
            .O(N__31145),
            .I(N__31118));
    Span4Mux_v I__7540 (
            .O(N__31140),
            .I(N__31118));
    Span4Mux_h I__7539 (
            .O(N__31137),
            .I(N__31118));
    LocalMux I__7538 (
            .O(N__31134),
            .I(N__31115));
    CascadeMux I__7537 (
            .O(N__31133),
            .I(N__31112));
    Span12Mux_v I__7536 (
            .O(N__31130),
            .I(N__31109));
    Span4Mux_v I__7535 (
            .O(N__31125),
            .I(N__31106));
    Span4Mux_v I__7534 (
            .O(N__31118),
            .I(N__31101));
    Span4Mux_h I__7533 (
            .O(N__31115),
            .I(N__31101));
    InMux I__7532 (
            .O(N__31112),
            .I(N__31098));
    Odrv12 I__7531 (
            .O(N__31109),
            .I(M_this_ppu_sprites_addr_9));
    Odrv4 I__7530 (
            .O(N__31106),
            .I(M_this_ppu_sprites_addr_9));
    Odrv4 I__7529 (
            .O(N__31101),
            .I(M_this_ppu_sprites_addr_9));
    LocalMux I__7528 (
            .O(N__31098),
            .I(M_this_ppu_sprites_addr_9));
    CascadeMux I__7527 (
            .O(N__31089),
            .I(N__31086));
    InMux I__7526 (
            .O(N__31086),
            .I(N__31083));
    LocalMux I__7525 (
            .O(N__31083),
            .I(N__31080));
    Span4Mux_v I__7524 (
            .O(N__31080),
            .I(N__31077));
    Odrv4 I__7523 (
            .O(N__31077),
            .I(M_this_data_tmp_qZ0Z_12));
    InMux I__7522 (
            .O(N__31074),
            .I(N__31071));
    LocalMux I__7521 (
            .O(N__31071),
            .I(N_740_0));
    InMux I__7520 (
            .O(N__31068),
            .I(N__31064));
    InMux I__7519 (
            .O(N__31067),
            .I(N__31060));
    LocalMux I__7518 (
            .O(N__31064),
            .I(N__31057));
    InMux I__7517 (
            .O(N__31063),
            .I(N__31054));
    LocalMux I__7516 (
            .O(N__31060),
            .I(N__31051));
    Span4Mux_h I__7515 (
            .O(N__31057),
            .I(N__31047));
    LocalMux I__7514 (
            .O(N__31054),
            .I(N__31042));
    Span4Mux_h I__7513 (
            .O(N__31051),
            .I(N__31042));
    InMux I__7512 (
            .O(N__31050),
            .I(N__31039));
    Span4Mux_h I__7511 (
            .O(N__31047),
            .I(N__31036));
    Span4Mux_h I__7510 (
            .O(N__31042),
            .I(N__31033));
    LocalMux I__7509 (
            .O(N__31039),
            .I(M_this_oam_ram_read_data_13));
    Odrv4 I__7508 (
            .O(N__31036),
            .I(M_this_oam_ram_read_data_13));
    Odrv4 I__7507 (
            .O(N__31033),
            .I(M_this_oam_ram_read_data_13));
    CascadeMux I__7506 (
            .O(N__31026),
            .I(N__31022));
    InMux I__7505 (
            .O(N__31025),
            .I(N__31018));
    InMux I__7504 (
            .O(N__31022),
            .I(N__31013));
    InMux I__7503 (
            .O(N__31021),
            .I(N__31013));
    LocalMux I__7502 (
            .O(N__31018),
            .I(N__31009));
    LocalMux I__7501 (
            .O(N__31013),
            .I(N__31006));
    InMux I__7500 (
            .O(N__31012),
            .I(N__31003));
    Span4Mux_h I__7499 (
            .O(N__31009),
            .I(N__30999));
    Span4Mux_h I__7498 (
            .O(N__31006),
            .I(N__30994));
    LocalMux I__7497 (
            .O(N__31003),
            .I(N__30994));
    InMux I__7496 (
            .O(N__31002),
            .I(N__30991));
    Span4Mux_h I__7495 (
            .O(N__30999),
            .I(N__30988));
    Span4Mux_h I__7494 (
            .O(N__30994),
            .I(N__30985));
    LocalMux I__7493 (
            .O(N__30991),
            .I(M_this_oam_ram_read_data_12));
    Odrv4 I__7492 (
            .O(N__30988),
            .I(M_this_oam_ram_read_data_12));
    Odrv4 I__7491 (
            .O(N__30985),
            .I(M_this_oam_ram_read_data_12));
    CascadeMux I__7490 (
            .O(N__30978),
            .I(N__30975));
    InMux I__7489 (
            .O(N__30975),
            .I(N__30971));
    InMux I__7488 (
            .O(N__30974),
            .I(N__30967));
    LocalMux I__7487 (
            .O(N__30971),
            .I(N__30964));
    CascadeMux I__7486 (
            .O(N__30970),
            .I(N__30961));
    LocalMux I__7485 (
            .O(N__30967),
            .I(N__30956));
    Span4Mux_h I__7484 (
            .O(N__30964),
            .I(N__30956));
    InMux I__7483 (
            .O(N__30961),
            .I(N__30953));
    Span4Mux_h I__7482 (
            .O(N__30956),
            .I(N__30950));
    LocalMux I__7481 (
            .O(N__30953),
            .I(M_this_oam_ram_read_data_14));
    Odrv4 I__7480 (
            .O(N__30950),
            .I(M_this_oam_ram_read_data_14));
    InMux I__7479 (
            .O(N__30945),
            .I(N__30937));
    InMux I__7478 (
            .O(N__30944),
            .I(N__30937));
    InMux I__7477 (
            .O(N__30943),
            .I(N__30934));
    InMux I__7476 (
            .O(N__30942),
            .I(N__30931));
    LocalMux I__7475 (
            .O(N__30937),
            .I(N__30927));
    LocalMux I__7474 (
            .O(N__30934),
            .I(N__30922));
    LocalMux I__7473 (
            .O(N__30931),
            .I(N__30922));
    InMux I__7472 (
            .O(N__30930),
            .I(N__30919));
    Span4Mux_v I__7471 (
            .O(N__30927),
            .I(N__30915));
    Span4Mux_h I__7470 (
            .O(N__30922),
            .I(N__30910));
    LocalMux I__7469 (
            .O(N__30919),
            .I(N__30910));
    InMux I__7468 (
            .O(N__30918),
            .I(N__30907));
    Span4Mux_h I__7467 (
            .O(N__30915),
            .I(N__30902));
    Span4Mux_v I__7466 (
            .O(N__30910),
            .I(N__30902));
    LocalMux I__7465 (
            .O(N__30907),
            .I(M_this_oam_ram_read_data_11));
    Odrv4 I__7464 (
            .O(N__30902),
            .I(M_this_oam_ram_read_data_11));
    CascadeMux I__7463 (
            .O(N__30897),
            .I(N__30894));
    InMux I__7462 (
            .O(N__30894),
            .I(N__30891));
    LocalMux I__7461 (
            .O(N__30891),
            .I(N__30888));
    Span12Mux_v I__7460 (
            .O(N__30888),
            .I(N__30885));
    Odrv12 I__7459 (
            .O(N__30885),
            .I(\this_ppu.un1_M_haddress_q_2_6 ));
    CascadeMux I__7458 (
            .O(N__30882),
            .I(N__30879));
    InMux I__7457 (
            .O(N__30879),
            .I(N__30876));
    LocalMux I__7456 (
            .O(N__30876),
            .I(N__30873));
    Span4Mux_v I__7455 (
            .O(N__30873),
            .I(N__30870));
    Odrv4 I__7454 (
            .O(N__30870),
            .I(M_this_data_tmp_qZ0Z_19));
    InMux I__7453 (
            .O(N__30867),
            .I(N__30864));
    LocalMux I__7452 (
            .O(N__30864),
            .I(N__30861));
    Span4Mux_v I__7451 (
            .O(N__30861),
            .I(N__30858));
    Odrv4 I__7450 (
            .O(N__30858),
            .I(M_this_oam_ram_write_data_19));
    CascadeMux I__7449 (
            .O(N__30855),
            .I(N__30852));
    InMux I__7448 (
            .O(N__30852),
            .I(N__30849));
    LocalMux I__7447 (
            .O(N__30849),
            .I(N__30846));
    Span4Mux_h I__7446 (
            .O(N__30846),
            .I(N__30843));
    Span4Mux_h I__7445 (
            .O(N__30843),
            .I(N__30837));
    InMux I__7444 (
            .O(N__30842),
            .I(N__30834));
    InMux I__7443 (
            .O(N__30841),
            .I(N__30831));
    InMux I__7442 (
            .O(N__30840),
            .I(N__30828));
    Span4Mux_h I__7441 (
            .O(N__30837),
            .I(N__30825));
    LocalMux I__7440 (
            .O(N__30834),
            .I(N__30818));
    LocalMux I__7439 (
            .O(N__30831),
            .I(N__30813));
    LocalMux I__7438 (
            .O(N__30828),
            .I(N__30813));
    Sp12to4 I__7437 (
            .O(N__30825),
            .I(N__30809));
    InMux I__7436 (
            .O(N__30824),
            .I(N__30802));
    InMux I__7435 (
            .O(N__30823),
            .I(N__30802));
    InMux I__7434 (
            .O(N__30822),
            .I(N__30802));
    InMux I__7433 (
            .O(N__30821),
            .I(N__30799));
    Span4Mux_v I__7432 (
            .O(N__30818),
            .I(N__30794));
    Span4Mux_h I__7431 (
            .O(N__30813),
            .I(N__30794));
    InMux I__7430 (
            .O(N__30812),
            .I(N__30791));
    Odrv12 I__7429 (
            .O(N__30809),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__7428 (
            .O(N__30802),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__7427 (
            .O(N__30799),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__7426 (
            .O(N__30794),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__7425 (
            .O(N__30791),
            .I(M_this_ppu_vram_addr_7));
    CascadeMux I__7424 (
            .O(N__30780),
            .I(N__30775));
    CascadeMux I__7423 (
            .O(N__30779),
            .I(N__30772));
    InMux I__7422 (
            .O(N__30778),
            .I(N__30769));
    InMux I__7421 (
            .O(N__30775),
            .I(N__30766));
    InMux I__7420 (
            .O(N__30772),
            .I(N__30762));
    LocalMux I__7419 (
            .O(N__30769),
            .I(N__30759));
    LocalMux I__7418 (
            .O(N__30766),
            .I(N__30756));
    InMux I__7417 (
            .O(N__30765),
            .I(N__30753));
    LocalMux I__7416 (
            .O(N__30762),
            .I(N__30750));
    Span4Mux_h I__7415 (
            .O(N__30759),
            .I(N__30747));
    Span4Mux_h I__7414 (
            .O(N__30756),
            .I(N__30744));
    LocalMux I__7413 (
            .O(N__30753),
            .I(N__30741));
    Span4Mux_h I__7412 (
            .O(N__30750),
            .I(N__30738));
    Span4Mux_v I__7411 (
            .O(N__30747),
            .I(N__30735));
    Sp12to4 I__7410 (
            .O(N__30744),
            .I(N__30732));
    Span4Mux_v I__7409 (
            .O(N__30741),
            .I(N__30729));
    Span4Mux_v I__7408 (
            .O(N__30738),
            .I(N__30726));
    Span4Mux_v I__7407 (
            .O(N__30735),
            .I(N__30723));
    Span12Mux_v I__7406 (
            .O(N__30732),
            .I(N__30720));
    Span4Mux_v I__7405 (
            .O(N__30729),
            .I(N__30715));
    Span4Mux_h I__7404 (
            .O(N__30726),
            .I(N__30715));
    Odrv4 I__7403 (
            .O(N__30723),
            .I(M_this_oam_ram_read_data_16));
    Odrv12 I__7402 (
            .O(N__30720),
            .I(M_this_oam_ram_read_data_16));
    Odrv4 I__7401 (
            .O(N__30715),
            .I(M_this_oam_ram_read_data_16));
    CascadeMux I__7400 (
            .O(N__30708),
            .I(N__30705));
    InMux I__7399 (
            .O(N__30705),
            .I(N__30702));
    LocalMux I__7398 (
            .O(N__30702),
            .I(\this_ppu.M_this_oam_ram_read_data_i_16 ));
    InMux I__7397 (
            .O(N__30699),
            .I(N__30696));
    LocalMux I__7396 (
            .O(N__30696),
            .I(N__30691));
    CascadeMux I__7395 (
            .O(N__30695),
            .I(N__30687));
    CascadeMux I__7394 (
            .O(N__30694),
            .I(N__30684));
    Span4Mux_v I__7393 (
            .O(N__30691),
            .I(N__30680));
    InMux I__7392 (
            .O(N__30690),
            .I(N__30677));
    InMux I__7391 (
            .O(N__30687),
            .I(N__30671));
    InMux I__7390 (
            .O(N__30684),
            .I(N__30671));
    InMux I__7389 (
            .O(N__30683),
            .I(N__30668));
    Sp12to4 I__7388 (
            .O(N__30680),
            .I(N__30663));
    LocalMux I__7387 (
            .O(N__30677),
            .I(N__30663));
    InMux I__7386 (
            .O(N__30676),
            .I(N__30660));
    LocalMux I__7385 (
            .O(N__30671),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    LocalMux I__7384 (
            .O(N__30668),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv12 I__7383 (
            .O(N__30663),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    LocalMux I__7382 (
            .O(N__30660),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    InMux I__7381 (
            .O(N__30651),
            .I(N__30648));
    LocalMux I__7380 (
            .O(N__30648),
            .I(\this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0 ));
    InMux I__7379 (
            .O(N__30645),
            .I(\this_ppu.un2_vscroll_cry_0 ));
    InMux I__7378 (
            .O(N__30642),
            .I(N__30639));
    LocalMux I__7377 (
            .O(N__30639),
            .I(N__30636));
    Span4Mux_v I__7376 (
            .O(N__30636),
            .I(N__30628));
    InMux I__7375 (
            .O(N__30635),
            .I(N__30625));
    InMux I__7374 (
            .O(N__30634),
            .I(N__30617));
    InMux I__7373 (
            .O(N__30633),
            .I(N__30617));
    InMux I__7372 (
            .O(N__30632),
            .I(N__30617));
    InMux I__7371 (
            .O(N__30631),
            .I(N__30614));
    Sp12to4 I__7370 (
            .O(N__30628),
            .I(N__30609));
    LocalMux I__7369 (
            .O(N__30625),
            .I(N__30609));
    InMux I__7368 (
            .O(N__30624),
            .I(N__30606));
    LocalMux I__7367 (
            .O(N__30617),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    LocalMux I__7366 (
            .O(N__30614),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    Odrv12 I__7365 (
            .O(N__30609),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    LocalMux I__7364 (
            .O(N__30606),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    CascadeMux I__7363 (
            .O(N__30597),
            .I(N__30594));
    InMux I__7362 (
            .O(N__30594),
            .I(N__30591));
    LocalMux I__7361 (
            .O(N__30591),
            .I(N__30586));
    CascadeMux I__7360 (
            .O(N__30590),
            .I(N__30583));
    InMux I__7359 (
            .O(N__30589),
            .I(N__30580));
    Span4Mux_v I__7358 (
            .O(N__30586),
            .I(N__30577));
    InMux I__7357 (
            .O(N__30583),
            .I(N__30574));
    LocalMux I__7356 (
            .O(N__30580),
            .I(N__30571));
    Sp12to4 I__7355 (
            .O(N__30577),
            .I(N__30566));
    LocalMux I__7354 (
            .O(N__30574),
            .I(N__30566));
    Span12Mux_v I__7353 (
            .O(N__30571),
            .I(N__30563));
    Span12Mux_h I__7352 (
            .O(N__30566),
            .I(N__30560));
    Odrv12 I__7351 (
            .O(N__30563),
            .I(M_this_oam_ram_read_data_18));
    Odrv12 I__7350 (
            .O(N__30560),
            .I(M_this_oam_ram_read_data_18));
    InMux I__7349 (
            .O(N__30555),
            .I(\this_ppu.un2_vscroll_cry_1 ));
    InMux I__7348 (
            .O(N__30552),
            .I(N__30549));
    LocalMux I__7347 (
            .O(N__30549),
            .I(N__30546));
    Odrv4 I__7346 (
            .O(N__30546),
            .I(\this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0 ));
    InMux I__7345 (
            .O(N__30543),
            .I(N__30540));
    LocalMux I__7344 (
            .O(N__30540),
            .I(N__30537));
    Span4Mux_v I__7343 (
            .O(N__30537),
            .I(N__30534));
    Span4Mux_v I__7342 (
            .O(N__30534),
            .I(N__30531));
    Span4Mux_h I__7341 (
            .O(N__30531),
            .I(N__30528));
    Sp12to4 I__7340 (
            .O(N__30528),
            .I(N__30525));
    Span12Mux_h I__7339 (
            .O(N__30525),
            .I(N__30522));
    Odrv12 I__7338 (
            .O(N__30522),
            .I(M_this_map_ram_read_data_4));
    CascadeMux I__7337 (
            .O(N__30519),
            .I(N__30516));
    InMux I__7336 (
            .O(N__30516),
            .I(N__30511));
    CascadeMux I__7335 (
            .O(N__30515),
            .I(N__30508));
    CascadeMux I__7334 (
            .O(N__30514),
            .I(N__30504));
    LocalMux I__7333 (
            .O(N__30511),
            .I(N__30501));
    InMux I__7332 (
            .O(N__30508),
            .I(N__30498));
    CascadeMux I__7331 (
            .O(N__30507),
            .I(N__30495));
    InMux I__7330 (
            .O(N__30504),
            .I(N__30490));
    Span4Mux_h I__7329 (
            .O(N__30501),
            .I(N__30485));
    LocalMux I__7328 (
            .O(N__30498),
            .I(N__30485));
    InMux I__7327 (
            .O(N__30495),
            .I(N__30482));
    CascadeMux I__7326 (
            .O(N__30494),
            .I(N__30479));
    CascadeMux I__7325 (
            .O(N__30493),
            .I(N__30476));
    LocalMux I__7324 (
            .O(N__30490),
            .I(N__30471));
    Span4Mux_v I__7323 (
            .O(N__30485),
            .I(N__30466));
    LocalMux I__7322 (
            .O(N__30482),
            .I(N__30466));
    InMux I__7321 (
            .O(N__30479),
            .I(N__30463));
    InMux I__7320 (
            .O(N__30476),
            .I(N__30460));
    CascadeMux I__7319 (
            .O(N__30475),
            .I(N__30457));
    CascadeMux I__7318 (
            .O(N__30474),
            .I(N__30454));
    Span4Mux_h I__7317 (
            .O(N__30471),
            .I(N__30449));
    Span4Mux_v I__7316 (
            .O(N__30466),
            .I(N__30444));
    LocalMux I__7315 (
            .O(N__30463),
            .I(N__30444));
    LocalMux I__7314 (
            .O(N__30460),
            .I(N__30441));
    InMux I__7313 (
            .O(N__30457),
            .I(N__30438));
    InMux I__7312 (
            .O(N__30454),
            .I(N__30435));
    CascadeMux I__7311 (
            .O(N__30453),
            .I(N__30432));
    CascadeMux I__7310 (
            .O(N__30452),
            .I(N__30429));
    Span4Mux_v I__7309 (
            .O(N__30449),
            .I(N__30420));
    Span4Mux_h I__7308 (
            .O(N__30444),
            .I(N__30420));
    Span4Mux_s1_v I__7307 (
            .O(N__30441),
            .I(N__30413));
    LocalMux I__7306 (
            .O(N__30438),
            .I(N__30413));
    LocalMux I__7305 (
            .O(N__30435),
            .I(N__30413));
    InMux I__7304 (
            .O(N__30432),
            .I(N__30410));
    InMux I__7303 (
            .O(N__30429),
            .I(N__30407));
    CascadeMux I__7302 (
            .O(N__30428),
            .I(N__30404));
    CascadeMux I__7301 (
            .O(N__30427),
            .I(N__30401));
    CascadeMux I__7300 (
            .O(N__30426),
            .I(N__30398));
    CascadeMux I__7299 (
            .O(N__30425),
            .I(N__30395));
    Span4Mux_h I__7298 (
            .O(N__30420),
            .I(N__30391));
    Span4Mux_v I__7297 (
            .O(N__30413),
            .I(N__30386));
    LocalMux I__7296 (
            .O(N__30410),
            .I(N__30386));
    LocalMux I__7295 (
            .O(N__30407),
            .I(N__30383));
    InMux I__7294 (
            .O(N__30404),
            .I(N__30380));
    InMux I__7293 (
            .O(N__30401),
            .I(N__30377));
    InMux I__7292 (
            .O(N__30398),
            .I(N__30374));
    InMux I__7291 (
            .O(N__30395),
            .I(N__30371));
    CascadeMux I__7290 (
            .O(N__30394),
            .I(N__30368));
    Span4Mux_h I__7289 (
            .O(N__30391),
            .I(N__30364));
    Span4Mux_v I__7288 (
            .O(N__30386),
            .I(N__30355));
    Span4Mux_v I__7287 (
            .O(N__30383),
            .I(N__30355));
    LocalMux I__7286 (
            .O(N__30380),
            .I(N__30355));
    LocalMux I__7285 (
            .O(N__30377),
            .I(N__30355));
    LocalMux I__7284 (
            .O(N__30374),
            .I(N__30350));
    LocalMux I__7283 (
            .O(N__30371),
            .I(N__30350));
    InMux I__7282 (
            .O(N__30368),
            .I(N__30347));
    CascadeMux I__7281 (
            .O(N__30367),
            .I(N__30344));
    Span4Mux_h I__7280 (
            .O(N__30364),
            .I(N__30341));
    Span4Mux_v I__7279 (
            .O(N__30355),
            .I(N__30334));
    Span4Mux_v I__7278 (
            .O(N__30350),
            .I(N__30334));
    LocalMux I__7277 (
            .O(N__30347),
            .I(N__30334));
    InMux I__7276 (
            .O(N__30344),
            .I(N__30331));
    Odrv4 I__7275 (
            .O(N__30341),
            .I(M_this_ppu_sprites_addr_10));
    Odrv4 I__7274 (
            .O(N__30334),
            .I(M_this_ppu_sprites_addr_10));
    LocalMux I__7273 (
            .O(N__30331),
            .I(M_this_ppu_sprites_addr_10));
    InMux I__7272 (
            .O(N__30324),
            .I(N__30321));
    LocalMux I__7271 (
            .O(N__30321),
            .I(N__30314));
    InMux I__7270 (
            .O(N__30320),
            .I(N__30311));
    InMux I__7269 (
            .O(N__30319),
            .I(N__30308));
    InMux I__7268 (
            .O(N__30318),
            .I(N__30303));
    InMux I__7267 (
            .O(N__30317),
            .I(N__30303));
    Span4Mux_v I__7266 (
            .O(N__30314),
            .I(N__30296));
    LocalMux I__7265 (
            .O(N__30311),
            .I(N__30296));
    LocalMux I__7264 (
            .O(N__30308),
            .I(N__30296));
    LocalMux I__7263 (
            .O(N__30303),
            .I(N__30290));
    Span4Mux_v I__7262 (
            .O(N__30296),
            .I(N__30287));
    InMux I__7261 (
            .O(N__30295),
            .I(N__30284));
    InMux I__7260 (
            .O(N__30294),
            .I(N__30281));
    InMux I__7259 (
            .O(N__30293),
            .I(N__30276));
    Span4Mux_h I__7258 (
            .O(N__30290),
            .I(N__30273));
    Sp12to4 I__7257 (
            .O(N__30287),
            .I(N__30268));
    LocalMux I__7256 (
            .O(N__30284),
            .I(N__30268));
    LocalMux I__7255 (
            .O(N__30281),
            .I(N__30265));
    InMux I__7254 (
            .O(N__30280),
            .I(N__30262));
    InMux I__7253 (
            .O(N__30279),
            .I(N__30259));
    LocalMux I__7252 (
            .O(N__30276),
            .I(N__30256));
    Odrv4 I__7251 (
            .O(N__30273),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv12 I__7250 (
            .O(N__30268),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv4 I__7249 (
            .O(N__30265),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__7248 (
            .O(N__30262),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__7247 (
            .O(N__30259),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv4 I__7246 (
            .O(N__30256),
            .I(M_this_sprites_address_qZ0Z_11));
    InMux I__7245 (
            .O(N__30243),
            .I(N__30235));
    InMux I__7244 (
            .O(N__30242),
            .I(N__30232));
    InMux I__7243 (
            .O(N__30241),
            .I(N__30229));
    InMux I__7242 (
            .O(N__30240),
            .I(N__30226));
    InMux I__7241 (
            .O(N__30239),
            .I(N__30221));
    InMux I__7240 (
            .O(N__30238),
            .I(N__30221));
    LocalMux I__7239 (
            .O(N__30235),
            .I(N__30216));
    LocalMux I__7238 (
            .O(N__30232),
            .I(N__30213));
    LocalMux I__7237 (
            .O(N__30229),
            .I(N__30208));
    LocalMux I__7236 (
            .O(N__30226),
            .I(N__30208));
    LocalMux I__7235 (
            .O(N__30221),
            .I(N__30205));
    InMux I__7234 (
            .O(N__30220),
            .I(N__30202));
    InMux I__7233 (
            .O(N__30219),
            .I(N__30199));
    Span4Mux_h I__7232 (
            .O(N__30216),
            .I(N__30194));
    Span4Mux_v I__7231 (
            .O(N__30213),
            .I(N__30189));
    Span4Mux_v I__7230 (
            .O(N__30208),
            .I(N__30189));
    Span12Mux_h I__7229 (
            .O(N__30205),
            .I(N__30184));
    LocalMux I__7228 (
            .O(N__30202),
            .I(N__30184));
    LocalMux I__7227 (
            .O(N__30199),
            .I(N__30181));
    InMux I__7226 (
            .O(N__30198),
            .I(N__30178));
    InMux I__7225 (
            .O(N__30197),
            .I(N__30175));
    Odrv4 I__7224 (
            .O(N__30194),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__7223 (
            .O(N__30189),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv12 I__7222 (
            .O(N__30184),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__7221 (
            .O(N__30181),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__7220 (
            .O(N__30178),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__7219 (
            .O(N__30175),
            .I(M_this_sprites_address_qZ0Z_12));
    CascadeMux I__7218 (
            .O(N__30162),
            .I(N__30154));
    CascadeMux I__7217 (
            .O(N__30161),
            .I(N__30151));
    CascadeMux I__7216 (
            .O(N__30160),
            .I(N__30148));
    CascadeMux I__7215 (
            .O(N__30159),
            .I(N__30145));
    CascadeMux I__7214 (
            .O(N__30158),
            .I(N__30141));
    CascadeMux I__7213 (
            .O(N__30157),
            .I(N__30138));
    InMux I__7212 (
            .O(N__30154),
            .I(N__30133));
    InMux I__7211 (
            .O(N__30151),
            .I(N__30133));
    InMux I__7210 (
            .O(N__30148),
            .I(N__30130));
    InMux I__7209 (
            .O(N__30145),
            .I(N__30127));
    CascadeMux I__7208 (
            .O(N__30144),
            .I(N__30124));
    InMux I__7207 (
            .O(N__30141),
            .I(N__30120));
    InMux I__7206 (
            .O(N__30138),
            .I(N__30117));
    LocalMux I__7205 (
            .O(N__30133),
            .I(N__30114));
    LocalMux I__7204 (
            .O(N__30130),
            .I(N__30109));
    LocalMux I__7203 (
            .O(N__30127),
            .I(N__30109));
    InMux I__7202 (
            .O(N__30124),
            .I(N__30106));
    CascadeMux I__7201 (
            .O(N__30123),
            .I(N__30103));
    LocalMux I__7200 (
            .O(N__30120),
            .I(N__30099));
    LocalMux I__7199 (
            .O(N__30117),
            .I(N__30096));
    Span4Mux_v I__7198 (
            .O(N__30114),
            .I(N__30093));
    Span4Mux_v I__7197 (
            .O(N__30109),
            .I(N__30088));
    LocalMux I__7196 (
            .O(N__30106),
            .I(N__30088));
    InMux I__7195 (
            .O(N__30103),
            .I(N__30085));
    InMux I__7194 (
            .O(N__30102),
            .I(N__30081));
    Span4Mux_h I__7193 (
            .O(N__30099),
            .I(N__30076));
    Span4Mux_h I__7192 (
            .O(N__30096),
            .I(N__30076));
    Span4Mux_h I__7191 (
            .O(N__30093),
            .I(N__30071));
    Span4Mux_h I__7190 (
            .O(N__30088),
            .I(N__30071));
    LocalMux I__7189 (
            .O(N__30085),
            .I(N__30068));
    InMux I__7188 (
            .O(N__30084),
            .I(N__30065));
    LocalMux I__7187 (
            .O(N__30081),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__7186 (
            .O(N__30076),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__7185 (
            .O(N__30071),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__7184 (
            .O(N__30068),
            .I(M_this_sprites_address_qZ0Z_13));
    LocalMux I__7183 (
            .O(N__30065),
            .I(M_this_sprites_address_qZ0Z_13));
    InMux I__7182 (
            .O(N__30054),
            .I(N__30044));
    InMux I__7181 (
            .O(N__30053),
            .I(N__30041));
    InMux I__7180 (
            .O(N__30052),
            .I(N__30038));
    InMux I__7179 (
            .O(N__30051),
            .I(N__30035));
    InMux I__7178 (
            .O(N__30050),
            .I(N__30032));
    InMux I__7177 (
            .O(N__30049),
            .I(N__30029));
    InMux I__7176 (
            .O(N__30048),
            .I(N__30024));
    InMux I__7175 (
            .O(N__30047),
            .I(N__30024));
    LocalMux I__7174 (
            .O(N__30044),
            .I(N__30021));
    LocalMux I__7173 (
            .O(N__30041),
            .I(N__30018));
    LocalMux I__7172 (
            .O(N__30038),
            .I(N__30015));
    LocalMux I__7171 (
            .O(N__30035),
            .I(N__30010));
    LocalMux I__7170 (
            .O(N__30032),
            .I(N__30010));
    LocalMux I__7169 (
            .O(N__30029),
            .I(N__30007));
    LocalMux I__7168 (
            .O(N__30024),
            .I(N__30004));
    Span4Mux_v I__7167 (
            .O(N__30021),
            .I(N__29999));
    Span4Mux_v I__7166 (
            .O(N__30018),
            .I(N__29999));
    Span4Mux_v I__7165 (
            .O(N__30015),
            .I(N__29990));
    Span4Mux_v I__7164 (
            .O(N__30010),
            .I(N__29990));
    Span4Mux_h I__7163 (
            .O(N__30007),
            .I(N__29990));
    Span4Mux_h I__7162 (
            .O(N__30004),
            .I(N__29990));
    Odrv4 I__7161 (
            .O(N__29999),
            .I(N_23_0));
    Odrv4 I__7160 (
            .O(N__29990),
            .I(N_23_0));
    CEMux I__7159 (
            .O(N__29985),
            .I(N__29981));
    CEMux I__7158 (
            .O(N__29984),
            .I(N__29978));
    LocalMux I__7157 (
            .O(N__29981),
            .I(\this_sprites_ram.mem_WE_2 ));
    LocalMux I__7156 (
            .O(N__29978),
            .I(\this_sprites_ram.mem_WE_2 ));
    InMux I__7155 (
            .O(N__29973),
            .I(N__29970));
    LocalMux I__7154 (
            .O(N__29970),
            .I(N__29966));
    CascadeMux I__7153 (
            .O(N__29969),
            .I(N__29962));
    Span4Mux_h I__7152 (
            .O(N__29966),
            .I(N__29958));
    InMux I__7151 (
            .O(N__29965),
            .I(N__29955));
    InMux I__7150 (
            .O(N__29962),
            .I(N__29952));
    InMux I__7149 (
            .O(N__29961),
            .I(N__29944));
    Span4Mux_h I__7148 (
            .O(N__29958),
            .I(N__29939));
    LocalMux I__7147 (
            .O(N__29955),
            .I(N__29939));
    LocalMux I__7146 (
            .O(N__29952),
            .I(N__29936));
    InMux I__7145 (
            .O(N__29951),
            .I(N__29931));
    InMux I__7144 (
            .O(N__29950),
            .I(N__29931));
    InMux I__7143 (
            .O(N__29949),
            .I(N__29924));
    InMux I__7142 (
            .O(N__29948),
            .I(N__29924));
    InMux I__7141 (
            .O(N__29947),
            .I(N__29924));
    LocalMux I__7140 (
            .O(N__29944),
            .I(N__29921));
    Span4Mux_v I__7139 (
            .O(N__29939),
            .I(N__29918));
    Span12Mux_h I__7138 (
            .O(N__29936),
            .I(N__29915));
    LocalMux I__7137 (
            .O(N__29931),
            .I(N__29906));
    LocalMux I__7136 (
            .O(N__29924),
            .I(N__29906));
    Span4Mux_v I__7135 (
            .O(N__29921),
            .I(N__29906));
    Span4Mux_v I__7134 (
            .O(N__29918),
            .I(N__29906));
    Odrv12 I__7133 (
            .O(N__29915),
            .I(M_this_ppu_vram_addr_0));
    Odrv4 I__7132 (
            .O(N__29906),
            .I(M_this_ppu_vram_addr_0));
    CascadeMux I__7131 (
            .O(N__29901),
            .I(N__29898));
    InMux I__7130 (
            .O(N__29898),
            .I(N__29892));
    CascadeMux I__7129 (
            .O(N__29897),
            .I(N__29889));
    InMux I__7128 (
            .O(N__29896),
            .I(N__29886));
    InMux I__7127 (
            .O(N__29895),
            .I(N__29883));
    LocalMux I__7126 (
            .O(N__29892),
            .I(N__29880));
    InMux I__7125 (
            .O(N__29889),
            .I(N__29877));
    LocalMux I__7124 (
            .O(N__29886),
            .I(N__29874));
    LocalMux I__7123 (
            .O(N__29883),
            .I(N__29871));
    Span4Mux_h I__7122 (
            .O(N__29880),
            .I(N__29866));
    LocalMux I__7121 (
            .O(N__29877),
            .I(N__29866));
    Span12Mux_h I__7120 (
            .O(N__29874),
            .I(N__29863));
    Span4Mux_h I__7119 (
            .O(N__29871),
            .I(N__29858));
    Span4Mux_h I__7118 (
            .O(N__29866),
            .I(N__29858));
    Span12Mux_v I__7117 (
            .O(N__29863),
            .I(N__29855));
    Span4Mux_v I__7116 (
            .O(N__29858),
            .I(N__29852));
    Odrv12 I__7115 (
            .O(N__29855),
            .I(M_this_oam_ram_read_data_8));
    Odrv4 I__7114 (
            .O(N__29852),
            .I(M_this_oam_ram_read_data_8));
    CascadeMux I__7113 (
            .O(N__29847),
            .I(N__29844));
    InMux I__7112 (
            .O(N__29844),
            .I(N__29841));
    LocalMux I__7111 (
            .O(N__29841),
            .I(\this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ));
    InMux I__7110 (
            .O(N__29838),
            .I(N__29833));
    InMux I__7109 (
            .O(N__29837),
            .I(N__29830));
    CascadeMux I__7108 (
            .O(N__29836),
            .I(N__29827));
    LocalMux I__7107 (
            .O(N__29833),
            .I(N__29821));
    LocalMux I__7106 (
            .O(N__29830),
            .I(N__29821));
    InMux I__7105 (
            .O(N__29827),
            .I(N__29817));
    InMux I__7104 (
            .O(N__29826),
            .I(N__29814));
    Span4Mux_h I__7103 (
            .O(N__29821),
            .I(N__29811));
    InMux I__7102 (
            .O(N__29820),
            .I(N__29808));
    LocalMux I__7101 (
            .O(N__29817),
            .I(N__29805));
    LocalMux I__7100 (
            .O(N__29814),
            .I(N__29801));
    Span4Mux_h I__7099 (
            .O(N__29811),
            .I(N__29796));
    LocalMux I__7098 (
            .O(N__29808),
            .I(N__29796));
    Sp12to4 I__7097 (
            .O(N__29805),
            .I(N__29793));
    InMux I__7096 (
            .O(N__29804),
            .I(N__29789));
    Span4Mux_v I__7095 (
            .O(N__29801),
            .I(N__29784));
    Span4Mux_v I__7094 (
            .O(N__29796),
            .I(N__29784));
    Span12Mux_s10_v I__7093 (
            .O(N__29793),
            .I(N__29781));
    InMux I__7092 (
            .O(N__29792),
            .I(N__29778));
    LocalMux I__7091 (
            .O(N__29789),
            .I(N__29773));
    Span4Mux_v I__7090 (
            .O(N__29784),
            .I(N__29773));
    Odrv12 I__7089 (
            .O(N__29781),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__7088 (
            .O(N__29778),
            .I(M_this_ppu_vram_addr_1));
    Odrv4 I__7087 (
            .O(N__29773),
            .I(M_this_ppu_vram_addr_1));
    InMux I__7086 (
            .O(N__29766),
            .I(N__29763));
    LocalMux I__7085 (
            .O(N__29763),
            .I(\this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0 ));
    InMux I__7084 (
            .O(N__29760),
            .I(\this_ppu.un2_hscroll_cry_0 ));
    CascadeMux I__7083 (
            .O(N__29757),
            .I(N__29754));
    InMux I__7082 (
            .O(N__29754),
            .I(N__29750));
    InMux I__7081 (
            .O(N__29753),
            .I(N__29747));
    LocalMux I__7080 (
            .O(N__29750),
            .I(N__29744));
    LocalMux I__7079 (
            .O(N__29747),
            .I(N__29738));
    Span4Mux_v I__7078 (
            .O(N__29744),
            .I(N__29735));
    CascadeMux I__7077 (
            .O(N__29743),
            .I(N__29731));
    CascadeMux I__7076 (
            .O(N__29742),
            .I(N__29728));
    InMux I__7075 (
            .O(N__29741),
            .I(N__29723));
    Sp12to4 I__7074 (
            .O(N__29738),
            .I(N__29720));
    Sp12to4 I__7073 (
            .O(N__29735),
            .I(N__29717));
    InMux I__7072 (
            .O(N__29734),
            .I(N__29714));
    InMux I__7071 (
            .O(N__29731),
            .I(N__29707));
    InMux I__7070 (
            .O(N__29728),
            .I(N__29707));
    InMux I__7069 (
            .O(N__29727),
            .I(N__29707));
    InMux I__7068 (
            .O(N__29726),
            .I(N__29704));
    LocalMux I__7067 (
            .O(N__29723),
            .I(N__29699));
    Span12Mux_v I__7066 (
            .O(N__29720),
            .I(N__29699));
    Span12Mux_h I__7065 (
            .O(N__29717),
            .I(N__29694));
    LocalMux I__7064 (
            .O(N__29714),
            .I(N__29694));
    LocalMux I__7063 (
            .O(N__29707),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__7062 (
            .O(N__29704),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__7061 (
            .O(N__29699),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__7060 (
            .O(N__29694),
            .I(M_this_ppu_vram_addr_2));
    InMux I__7059 (
            .O(N__29685),
            .I(N__29682));
    LocalMux I__7058 (
            .O(N__29682),
            .I(N__29679));
    Odrv4 I__7057 (
            .O(N__29679),
            .I(M_this_oam_ram_write_data_30));
    InMux I__7056 (
            .O(N__29676),
            .I(N__29673));
    LocalMux I__7055 (
            .O(N__29673),
            .I(\this_sprites_ram.mem_out_bus5_1 ));
    InMux I__7054 (
            .O(N__29670),
            .I(N__29667));
    LocalMux I__7053 (
            .O(N__29667),
            .I(N__29664));
    Span4Mux_v I__7052 (
            .O(N__29664),
            .I(N__29661));
    Odrv4 I__7051 (
            .O(N__29661),
            .I(\this_sprites_ram.mem_out_bus1_1 ));
    InMux I__7050 (
            .O(N__29658),
            .I(N__29653));
    InMux I__7049 (
            .O(N__29657),
            .I(N__29643));
    InMux I__7048 (
            .O(N__29656),
            .I(N__29643));
    LocalMux I__7047 (
            .O(N__29653),
            .I(N__29640));
    InMux I__7046 (
            .O(N__29652),
            .I(N__29637));
    InMux I__7045 (
            .O(N__29651),
            .I(N__29634));
    CascadeMux I__7044 (
            .O(N__29650),
            .I(N__29624));
    InMux I__7043 (
            .O(N__29649),
            .I(N__29618));
    InMux I__7042 (
            .O(N__29648),
            .I(N__29618));
    LocalMux I__7041 (
            .O(N__29643),
            .I(N__29611));
    Span4Mux_v I__7040 (
            .O(N__29640),
            .I(N__29611));
    LocalMux I__7039 (
            .O(N__29637),
            .I(N__29611));
    LocalMux I__7038 (
            .O(N__29634),
            .I(N__29608));
    InMux I__7037 (
            .O(N__29633),
            .I(N__29605));
    InMux I__7036 (
            .O(N__29632),
            .I(N__29600));
    InMux I__7035 (
            .O(N__29631),
            .I(N__29600));
    InMux I__7034 (
            .O(N__29630),
            .I(N__29597));
    InMux I__7033 (
            .O(N__29629),
            .I(N__29594));
    InMux I__7032 (
            .O(N__29628),
            .I(N__29591));
    InMux I__7031 (
            .O(N__29627),
            .I(N__29584));
    InMux I__7030 (
            .O(N__29624),
            .I(N__29584));
    InMux I__7029 (
            .O(N__29623),
            .I(N__29584));
    LocalMux I__7028 (
            .O(N__29618),
            .I(N__29581));
    Span4Mux_h I__7027 (
            .O(N__29611),
            .I(N__29574));
    Span4Mux_v I__7026 (
            .O(N__29608),
            .I(N__29574));
    LocalMux I__7025 (
            .O(N__29605),
            .I(N__29574));
    LocalMux I__7024 (
            .O(N__29600),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    LocalMux I__7023 (
            .O(N__29597),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    LocalMux I__7022 (
            .O(N__29594),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    LocalMux I__7021 (
            .O(N__29591),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    LocalMux I__7020 (
            .O(N__29584),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__7019 (
            .O(N__29581),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__7018 (
            .O(N__29574),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    InMux I__7017 (
            .O(N__29559),
            .I(N__29556));
    LocalMux I__7016 (
            .O(N__29556),
            .I(N__29553));
    Span4Mux_h I__7015 (
            .O(N__29553),
            .I(N__29550));
    Odrv4 I__7014 (
            .O(N__29550),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ));
    CascadeMux I__7013 (
            .O(N__29547),
            .I(N__29544));
    InMux I__7012 (
            .O(N__29544),
            .I(N__29539));
    CascadeMux I__7011 (
            .O(N__29543),
            .I(N__29536));
    CascadeMux I__7010 (
            .O(N__29542),
            .I(N__29532));
    LocalMux I__7009 (
            .O(N__29539),
            .I(N__29529));
    InMux I__7008 (
            .O(N__29536),
            .I(N__29526));
    CascadeMux I__7007 (
            .O(N__29535),
            .I(N__29523));
    InMux I__7006 (
            .O(N__29532),
            .I(N__29516));
    Span4Mux_h I__7005 (
            .O(N__29529),
            .I(N__29511));
    LocalMux I__7004 (
            .O(N__29526),
            .I(N__29511));
    InMux I__7003 (
            .O(N__29523),
            .I(N__29508));
    CascadeMux I__7002 (
            .O(N__29522),
            .I(N__29504));
    CascadeMux I__7001 (
            .O(N__29521),
            .I(N__29500));
    CascadeMux I__7000 (
            .O(N__29520),
            .I(N__29496));
    CascadeMux I__6999 (
            .O(N__29519),
            .I(N__29493));
    LocalMux I__6998 (
            .O(N__29516),
            .I(N__29484));
    Span4Mux_v I__6997 (
            .O(N__29511),
            .I(N__29484));
    LocalMux I__6996 (
            .O(N__29508),
            .I(N__29484));
    CascadeMux I__6995 (
            .O(N__29507),
            .I(N__29481));
    InMux I__6994 (
            .O(N__29504),
            .I(N__29478));
    CascadeMux I__6993 (
            .O(N__29503),
            .I(N__29475));
    InMux I__6992 (
            .O(N__29500),
            .I(N__29471));
    CascadeMux I__6991 (
            .O(N__29499),
            .I(N__29468));
    InMux I__6990 (
            .O(N__29496),
            .I(N__29465));
    InMux I__6989 (
            .O(N__29493),
            .I(N__29462));
    CascadeMux I__6988 (
            .O(N__29492),
            .I(N__29459));
    CascadeMux I__6987 (
            .O(N__29491),
            .I(N__29456));
    Span4Mux_v I__6986 (
            .O(N__29484),
            .I(N__29452));
    InMux I__6985 (
            .O(N__29481),
            .I(N__29449));
    LocalMux I__6984 (
            .O(N__29478),
            .I(N__29446));
    InMux I__6983 (
            .O(N__29475),
            .I(N__29443));
    CascadeMux I__6982 (
            .O(N__29474),
            .I(N__29440));
    LocalMux I__6981 (
            .O(N__29471),
            .I(N__29437));
    InMux I__6980 (
            .O(N__29468),
            .I(N__29434));
    LocalMux I__6979 (
            .O(N__29465),
            .I(N__29429));
    LocalMux I__6978 (
            .O(N__29462),
            .I(N__29429));
    InMux I__6977 (
            .O(N__29459),
            .I(N__29426));
    InMux I__6976 (
            .O(N__29456),
            .I(N__29423));
    CascadeMux I__6975 (
            .O(N__29455),
            .I(N__29420));
    Sp12to4 I__6974 (
            .O(N__29452),
            .I(N__29414));
    LocalMux I__6973 (
            .O(N__29449),
            .I(N__29414));
    Span4Mux_s3_v I__6972 (
            .O(N__29446),
            .I(N__29409));
    LocalMux I__6971 (
            .O(N__29443),
            .I(N__29409));
    InMux I__6970 (
            .O(N__29440),
            .I(N__29406));
    Span4Mux_v I__6969 (
            .O(N__29437),
            .I(N__29401));
    LocalMux I__6968 (
            .O(N__29434),
            .I(N__29401));
    Span4Mux_v I__6967 (
            .O(N__29429),
            .I(N__29394));
    LocalMux I__6966 (
            .O(N__29426),
            .I(N__29394));
    LocalMux I__6965 (
            .O(N__29423),
            .I(N__29394));
    InMux I__6964 (
            .O(N__29420),
            .I(N__29391));
    CascadeMux I__6963 (
            .O(N__29419),
            .I(N__29388));
    Span12Mux_h I__6962 (
            .O(N__29414),
            .I(N__29385));
    Span4Mux_v I__6961 (
            .O(N__29409),
            .I(N__29380));
    LocalMux I__6960 (
            .O(N__29406),
            .I(N__29380));
    Span4Mux_v I__6959 (
            .O(N__29401),
            .I(N__29373));
    Span4Mux_v I__6958 (
            .O(N__29394),
            .I(N__29373));
    LocalMux I__6957 (
            .O(N__29391),
            .I(N__29373));
    InMux I__6956 (
            .O(N__29388),
            .I(N__29370));
    Odrv12 I__6955 (
            .O(N__29385),
            .I(M_this_ppu_sprites_addr_2));
    Odrv4 I__6954 (
            .O(N__29380),
            .I(M_this_ppu_sprites_addr_2));
    Odrv4 I__6953 (
            .O(N__29373),
            .I(M_this_ppu_sprites_addr_2));
    LocalMux I__6952 (
            .O(N__29370),
            .I(M_this_ppu_sprites_addr_2));
    CEMux I__6951 (
            .O(N__29361),
            .I(N__29358));
    LocalMux I__6950 (
            .O(N__29358),
            .I(N__29355));
    Span4Mux_v I__6949 (
            .O(N__29355),
            .I(N__29351));
    CEMux I__6948 (
            .O(N__29354),
            .I(N__29348));
    Odrv4 I__6947 (
            .O(N__29351),
            .I(\this_sprites_ram.mem_WE_4 ));
    LocalMux I__6946 (
            .O(N__29348),
            .I(\this_sprites_ram.mem_WE_4 ));
    CEMux I__6945 (
            .O(N__29343),
            .I(N__29339));
    CEMux I__6944 (
            .O(N__29342),
            .I(N__29336));
    LocalMux I__6943 (
            .O(N__29339),
            .I(N__29331));
    LocalMux I__6942 (
            .O(N__29336),
            .I(N__29331));
    Span4Mux_v I__6941 (
            .O(N__29331),
            .I(N__29328));
    Odrv4 I__6940 (
            .O(N__29328),
            .I(\this_sprites_ram.mem_WE_12 ));
    CascadeMux I__6939 (
            .O(N__29325),
            .I(N__29320));
    CascadeMux I__6938 (
            .O(N__29324),
            .I(N__29317));
    CascadeMux I__6937 (
            .O(N__29323),
            .I(N__29312));
    InMux I__6936 (
            .O(N__29320),
            .I(N__29309));
    InMux I__6935 (
            .O(N__29317),
            .I(N__29306));
    CascadeMux I__6934 (
            .O(N__29316),
            .I(N__29303));
    CascadeMux I__6933 (
            .O(N__29315),
            .I(N__29300));
    InMux I__6932 (
            .O(N__29312),
            .I(N__29294));
    LocalMux I__6931 (
            .O(N__29309),
            .I(N__29291));
    LocalMux I__6930 (
            .O(N__29306),
            .I(N__29288));
    InMux I__6929 (
            .O(N__29303),
            .I(N__29285));
    InMux I__6928 (
            .O(N__29300),
            .I(N__29281));
    CascadeMux I__6927 (
            .O(N__29299),
            .I(N__29278));
    CascadeMux I__6926 (
            .O(N__29298),
            .I(N__29274));
    CascadeMux I__6925 (
            .O(N__29297),
            .I(N__29269));
    LocalMux I__6924 (
            .O(N__29294),
            .I(N__29265));
    Span4Mux_v I__6923 (
            .O(N__29291),
            .I(N__29258));
    Span4Mux_h I__6922 (
            .O(N__29288),
            .I(N__29258));
    LocalMux I__6921 (
            .O(N__29285),
            .I(N__29258));
    CascadeMux I__6920 (
            .O(N__29284),
            .I(N__29255));
    LocalMux I__6919 (
            .O(N__29281),
            .I(N__29252));
    InMux I__6918 (
            .O(N__29278),
            .I(N__29249));
    CascadeMux I__6917 (
            .O(N__29277),
            .I(N__29246));
    InMux I__6916 (
            .O(N__29274),
            .I(N__29243));
    CascadeMux I__6915 (
            .O(N__29273),
            .I(N__29240));
    CascadeMux I__6914 (
            .O(N__29272),
            .I(N__29237));
    InMux I__6913 (
            .O(N__29269),
            .I(N__29233));
    CascadeMux I__6912 (
            .O(N__29268),
            .I(N__29230));
    Span4Mux_v I__6911 (
            .O(N__29265),
            .I(N__29224));
    Span4Mux_v I__6910 (
            .O(N__29258),
            .I(N__29224));
    InMux I__6909 (
            .O(N__29255),
            .I(N__29221));
    Span4Mux_s3_v I__6908 (
            .O(N__29252),
            .I(N__29216));
    LocalMux I__6907 (
            .O(N__29249),
            .I(N__29216));
    InMux I__6906 (
            .O(N__29246),
            .I(N__29213));
    LocalMux I__6905 (
            .O(N__29243),
            .I(N__29210));
    InMux I__6904 (
            .O(N__29240),
            .I(N__29207));
    InMux I__6903 (
            .O(N__29237),
            .I(N__29204));
    CascadeMux I__6902 (
            .O(N__29236),
            .I(N__29201));
    LocalMux I__6901 (
            .O(N__29233),
            .I(N__29198));
    InMux I__6900 (
            .O(N__29230),
            .I(N__29195));
    CascadeMux I__6899 (
            .O(N__29229),
            .I(N__29192));
    Sp12to4 I__6898 (
            .O(N__29224),
            .I(N__29188));
    LocalMux I__6897 (
            .O(N__29221),
            .I(N__29185));
    Span4Mux_v I__6896 (
            .O(N__29216),
            .I(N__29180));
    LocalMux I__6895 (
            .O(N__29213),
            .I(N__29180));
    Span4Mux_v I__6894 (
            .O(N__29210),
            .I(N__29173));
    LocalMux I__6893 (
            .O(N__29207),
            .I(N__29173));
    LocalMux I__6892 (
            .O(N__29204),
            .I(N__29173));
    InMux I__6891 (
            .O(N__29201),
            .I(N__29170));
    Span4Mux_v I__6890 (
            .O(N__29198),
            .I(N__29165));
    LocalMux I__6889 (
            .O(N__29195),
            .I(N__29165));
    InMux I__6888 (
            .O(N__29192),
            .I(N__29162));
    CascadeMux I__6887 (
            .O(N__29191),
            .I(N__29159));
    Span12Mux_h I__6886 (
            .O(N__29188),
            .I(N__29156));
    Span12Mux_h I__6885 (
            .O(N__29185),
            .I(N__29153));
    Span4Mux_v I__6884 (
            .O(N__29180),
            .I(N__29146));
    Span4Mux_v I__6883 (
            .O(N__29173),
            .I(N__29146));
    LocalMux I__6882 (
            .O(N__29170),
            .I(N__29146));
    Span4Mux_v I__6881 (
            .O(N__29165),
            .I(N__29141));
    LocalMux I__6880 (
            .O(N__29162),
            .I(N__29141));
    InMux I__6879 (
            .O(N__29159),
            .I(N__29138));
    Odrv12 I__6878 (
            .O(N__29156),
            .I(M_this_ppu_sprites_addr_5));
    Odrv12 I__6877 (
            .O(N__29153),
            .I(M_this_ppu_sprites_addr_5));
    Odrv4 I__6876 (
            .O(N__29146),
            .I(M_this_ppu_sprites_addr_5));
    Odrv4 I__6875 (
            .O(N__29141),
            .I(M_this_ppu_sprites_addr_5));
    LocalMux I__6874 (
            .O(N__29138),
            .I(M_this_ppu_sprites_addr_5));
    InMux I__6873 (
            .O(N__29127),
            .I(N__29122));
    InMux I__6872 (
            .O(N__29126),
            .I(N__29117));
    InMux I__6871 (
            .O(N__29125),
            .I(N__29117));
    LocalMux I__6870 (
            .O(N__29122),
            .I(N__29106));
    LocalMux I__6869 (
            .O(N__29117),
            .I(N__29106));
    InMux I__6868 (
            .O(N__29116),
            .I(N__29101));
    InMux I__6867 (
            .O(N__29115),
            .I(N__29101));
    InMux I__6866 (
            .O(N__29114),
            .I(N__29098));
    InMux I__6865 (
            .O(N__29113),
            .I(N__29095));
    InMux I__6864 (
            .O(N__29112),
            .I(N__29092));
    InMux I__6863 (
            .O(N__29111),
            .I(N__29088));
    Span4Mux_v I__6862 (
            .O(N__29106),
            .I(N__29078));
    LocalMux I__6861 (
            .O(N__29101),
            .I(N__29078));
    LocalMux I__6860 (
            .O(N__29098),
            .I(N__29078));
    LocalMux I__6859 (
            .O(N__29095),
            .I(N__29078));
    LocalMux I__6858 (
            .O(N__29092),
            .I(N__29075));
    InMux I__6857 (
            .O(N__29091),
            .I(N__29072));
    LocalMux I__6856 (
            .O(N__29088),
            .I(N__29068));
    InMux I__6855 (
            .O(N__29087),
            .I(N__29065));
    Span4Mux_h I__6854 (
            .O(N__29078),
            .I(N__29062));
    Span4Mux_h I__6853 (
            .O(N__29075),
            .I(N__29057));
    LocalMux I__6852 (
            .O(N__29072),
            .I(N__29057));
    InMux I__6851 (
            .O(N__29071),
            .I(N__29054));
    Odrv12 I__6850 (
            .O(N__29068),
            .I(N_809));
    LocalMux I__6849 (
            .O(N__29065),
            .I(N_809));
    Odrv4 I__6848 (
            .O(N__29062),
            .I(N_809));
    Odrv4 I__6847 (
            .O(N__29057),
            .I(N_809));
    LocalMux I__6846 (
            .O(N__29054),
            .I(N_809));
    InMux I__6845 (
            .O(N__29043),
            .I(N__29040));
    LocalMux I__6844 (
            .O(N__29040),
            .I(N__29037));
    Span4Mux_v I__6843 (
            .O(N__29037),
            .I(N__29034));
    Odrv4 I__6842 (
            .O(N__29034),
            .I(M_this_sprites_address_q_RNO_0Z0Z_5));
    CascadeMux I__6841 (
            .O(N__29031),
            .I(N__29028));
    InMux I__6840 (
            .O(N__29028),
            .I(N__29025));
    LocalMux I__6839 (
            .O(N__29025),
            .I(N_595));
    CascadeMux I__6838 (
            .O(N__29022),
            .I(N__29013));
    CascadeMux I__6837 (
            .O(N__29021),
            .I(N__29004));
    CascadeMux I__6836 (
            .O(N__29020),
            .I(N__29000));
    CascadeMux I__6835 (
            .O(N__29019),
            .I(N__28996));
    InMux I__6834 (
            .O(N__29018),
            .I(N__28986));
    InMux I__6833 (
            .O(N__29017),
            .I(N__28986));
    InMux I__6832 (
            .O(N__29016),
            .I(N__28986));
    InMux I__6831 (
            .O(N__29013),
            .I(N__28983));
    InMux I__6830 (
            .O(N__29012),
            .I(N__28980));
    InMux I__6829 (
            .O(N__29011),
            .I(N__28973));
    InMux I__6828 (
            .O(N__29010),
            .I(N__28973));
    InMux I__6827 (
            .O(N__29009),
            .I(N__28973));
    InMux I__6826 (
            .O(N__29008),
            .I(N__28968));
    InMux I__6825 (
            .O(N__29007),
            .I(N__28968));
    InMux I__6824 (
            .O(N__29004),
            .I(N__28963));
    InMux I__6823 (
            .O(N__29003),
            .I(N__28963));
    InMux I__6822 (
            .O(N__29000),
            .I(N__28956));
    InMux I__6821 (
            .O(N__28999),
            .I(N__28956));
    InMux I__6820 (
            .O(N__28996),
            .I(N__28956));
    InMux I__6819 (
            .O(N__28995),
            .I(N__28951));
    InMux I__6818 (
            .O(N__28994),
            .I(N__28951));
    InMux I__6817 (
            .O(N__28993),
            .I(N__28948));
    LocalMux I__6816 (
            .O(N__28986),
            .I(N__28943));
    LocalMux I__6815 (
            .O(N__28983),
            .I(N__28938));
    LocalMux I__6814 (
            .O(N__28980),
            .I(N__28933));
    LocalMux I__6813 (
            .O(N__28973),
            .I(N__28933));
    LocalMux I__6812 (
            .O(N__28968),
            .I(N__28928));
    LocalMux I__6811 (
            .O(N__28963),
            .I(N__28928));
    LocalMux I__6810 (
            .O(N__28956),
            .I(N__28921));
    LocalMux I__6809 (
            .O(N__28951),
            .I(N__28921));
    LocalMux I__6808 (
            .O(N__28948),
            .I(N__28921));
    InMux I__6807 (
            .O(N__28947),
            .I(N__28918));
    CascadeMux I__6806 (
            .O(N__28946),
            .I(N__28915));
    Span4Mux_v I__6805 (
            .O(N__28943),
            .I(N__28911));
    InMux I__6804 (
            .O(N__28942),
            .I(N__28908));
    InMux I__6803 (
            .O(N__28941),
            .I(N__28905));
    Span4Mux_h I__6802 (
            .O(N__28938),
            .I(N__28894));
    Span4Mux_h I__6801 (
            .O(N__28933),
            .I(N__28894));
    Span4Mux_v I__6800 (
            .O(N__28928),
            .I(N__28894));
    Span4Mux_v I__6799 (
            .O(N__28921),
            .I(N__28894));
    LocalMux I__6798 (
            .O(N__28918),
            .I(N__28894));
    InMux I__6797 (
            .O(N__28915),
            .I(N__28891));
    InMux I__6796 (
            .O(N__28914),
            .I(N__28888));
    Sp12to4 I__6795 (
            .O(N__28911),
            .I(N__28881));
    LocalMux I__6794 (
            .O(N__28908),
            .I(N__28881));
    LocalMux I__6793 (
            .O(N__28905),
            .I(N__28881));
    Span4Mux_h I__6792 (
            .O(N__28894),
            .I(N__28878));
    LocalMux I__6791 (
            .O(N__28891),
            .I(N_383_0));
    LocalMux I__6790 (
            .O(N__28888),
            .I(N_383_0));
    Odrv12 I__6789 (
            .O(N__28881),
            .I(N_383_0));
    Odrv4 I__6788 (
            .O(N__28878),
            .I(N_383_0));
    CascadeMux I__6787 (
            .O(N__28869),
            .I(N__28865));
    CascadeMux I__6786 (
            .O(N__28868),
            .I(N__28862));
    InMux I__6785 (
            .O(N__28865),
            .I(N__28855));
    InMux I__6784 (
            .O(N__28862),
            .I(N__28852));
    CascadeMux I__6783 (
            .O(N__28861),
            .I(N__28849));
    CascadeMux I__6782 (
            .O(N__28860),
            .I(N__28846));
    CascadeMux I__6781 (
            .O(N__28859),
            .I(N__28842));
    CascadeMux I__6780 (
            .O(N__28858),
            .I(N__28839));
    LocalMux I__6779 (
            .O(N__28855),
            .I(N__28834));
    LocalMux I__6778 (
            .O(N__28852),
            .I(N__28831));
    InMux I__6777 (
            .O(N__28849),
            .I(N__28828));
    InMux I__6776 (
            .O(N__28846),
            .I(N__28825));
    CascadeMux I__6775 (
            .O(N__28845),
            .I(N__28821));
    InMux I__6774 (
            .O(N__28842),
            .I(N__28816));
    InMux I__6773 (
            .O(N__28839),
            .I(N__28813));
    CascadeMux I__6772 (
            .O(N__28838),
            .I(N__28810));
    CascadeMux I__6771 (
            .O(N__28837),
            .I(N__28807));
    Span4Mux_v I__6770 (
            .O(N__28834),
            .I(N__28798));
    Span4Mux_h I__6769 (
            .O(N__28831),
            .I(N__28798));
    LocalMux I__6768 (
            .O(N__28828),
            .I(N__28798));
    LocalMux I__6767 (
            .O(N__28825),
            .I(N__28795));
    CascadeMux I__6766 (
            .O(N__28824),
            .I(N__28792));
    InMux I__6765 (
            .O(N__28821),
            .I(N__28789));
    CascadeMux I__6764 (
            .O(N__28820),
            .I(N__28786));
    CascadeMux I__6763 (
            .O(N__28819),
            .I(N__28783));
    LocalMux I__6762 (
            .O(N__28816),
            .I(N__28778));
    LocalMux I__6761 (
            .O(N__28813),
            .I(N__28778));
    InMux I__6760 (
            .O(N__28810),
            .I(N__28775));
    InMux I__6759 (
            .O(N__28807),
            .I(N__28772));
    CascadeMux I__6758 (
            .O(N__28806),
            .I(N__28769));
    CascadeMux I__6757 (
            .O(N__28805),
            .I(N__28766));
    Span4Mux_v I__6756 (
            .O(N__28798),
            .I(N__28759));
    Span4Mux_v I__6755 (
            .O(N__28795),
            .I(N__28759));
    InMux I__6754 (
            .O(N__28792),
            .I(N__28756));
    LocalMux I__6753 (
            .O(N__28789),
            .I(N__28753));
    InMux I__6752 (
            .O(N__28786),
            .I(N__28750));
    InMux I__6751 (
            .O(N__28783),
            .I(N__28747));
    Span4Mux_v I__6750 (
            .O(N__28778),
            .I(N__28740));
    LocalMux I__6749 (
            .O(N__28775),
            .I(N__28740));
    LocalMux I__6748 (
            .O(N__28772),
            .I(N__28740));
    InMux I__6747 (
            .O(N__28769),
            .I(N__28737));
    InMux I__6746 (
            .O(N__28766),
            .I(N__28734));
    CascadeMux I__6745 (
            .O(N__28765),
            .I(N__28731));
    InMux I__6744 (
            .O(N__28764),
            .I(N__28727));
    Sp12to4 I__6743 (
            .O(N__28759),
            .I(N__28722));
    LocalMux I__6742 (
            .O(N__28756),
            .I(N__28722));
    Span4Mux_v I__6741 (
            .O(N__28753),
            .I(N__28715));
    LocalMux I__6740 (
            .O(N__28750),
            .I(N__28715));
    LocalMux I__6739 (
            .O(N__28747),
            .I(N__28715));
    Span4Mux_v I__6738 (
            .O(N__28740),
            .I(N__28708));
    LocalMux I__6737 (
            .O(N__28737),
            .I(N__28708));
    LocalMux I__6736 (
            .O(N__28734),
            .I(N__28708));
    InMux I__6735 (
            .O(N__28731),
            .I(N__28705));
    CascadeMux I__6734 (
            .O(N__28730),
            .I(N__28702));
    LocalMux I__6733 (
            .O(N__28727),
            .I(N__28698));
    Span12Mux_h I__6732 (
            .O(N__28722),
            .I(N__28695));
    Span4Mux_v I__6731 (
            .O(N__28715),
            .I(N__28688));
    Span4Mux_v I__6730 (
            .O(N__28708),
            .I(N__28688));
    LocalMux I__6729 (
            .O(N__28705),
            .I(N__28688));
    InMux I__6728 (
            .O(N__28702),
            .I(N__28685));
    InMux I__6727 (
            .O(N__28701),
            .I(N__28682));
    Span4Mux_h I__6726 (
            .O(N__28698),
            .I(N__28679));
    Odrv12 I__6725 (
            .O(N__28695),
            .I(M_this_sprites_address_qZ0Z_5));
    Odrv4 I__6724 (
            .O(N__28688),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__6723 (
            .O(N__28685),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__6722 (
            .O(N__28682),
            .I(M_this_sprites_address_qZ0Z_5));
    Odrv4 I__6721 (
            .O(N__28679),
            .I(M_this_sprites_address_qZ0Z_5));
    SRMux I__6720 (
            .O(N__28668),
            .I(N__28632));
    SRMux I__6719 (
            .O(N__28667),
            .I(N__28632));
    SRMux I__6718 (
            .O(N__28666),
            .I(N__28632));
    SRMux I__6717 (
            .O(N__28665),
            .I(N__28632));
    SRMux I__6716 (
            .O(N__28664),
            .I(N__28632));
    SRMux I__6715 (
            .O(N__28663),
            .I(N__28632));
    SRMux I__6714 (
            .O(N__28662),
            .I(N__28632));
    SRMux I__6713 (
            .O(N__28661),
            .I(N__28632));
    SRMux I__6712 (
            .O(N__28660),
            .I(N__28632));
    SRMux I__6711 (
            .O(N__28659),
            .I(N__28632));
    SRMux I__6710 (
            .O(N__28658),
            .I(N__28632));
    SRMux I__6709 (
            .O(N__28657),
            .I(N__28632));
    GlobalMux I__6708 (
            .O(N__28632),
            .I(N__28629));
    gio2CtrlBuf I__6707 (
            .O(N__28629),
            .I(N_515_g));
    CEMux I__6706 (
            .O(N__28626),
            .I(N__28622));
    CEMux I__6705 (
            .O(N__28625),
            .I(N__28619));
    LocalMux I__6704 (
            .O(N__28622),
            .I(N__28614));
    LocalMux I__6703 (
            .O(N__28619),
            .I(N__28614));
    Span4Mux_v I__6702 (
            .O(N__28614),
            .I(N__28611));
    Odrv4 I__6701 (
            .O(N__28611),
            .I(\this_sprites_ram.mem_WE_0 ));
    CascadeMux I__6700 (
            .O(N__28608),
            .I(N__28605));
    InMux I__6699 (
            .O(N__28605),
            .I(N__28600));
    CascadeMux I__6698 (
            .O(N__28604),
            .I(N__28597));
    CascadeMux I__6697 (
            .O(N__28603),
            .I(N__28594));
    LocalMux I__6696 (
            .O(N__28600),
            .I(N__28588));
    InMux I__6695 (
            .O(N__28597),
            .I(N__28585));
    InMux I__6694 (
            .O(N__28594),
            .I(N__28582));
    CascadeMux I__6693 (
            .O(N__28593),
            .I(N__28579));
    CascadeMux I__6692 (
            .O(N__28592),
            .I(N__28575));
    CascadeMux I__6691 (
            .O(N__28591),
            .I(N__28571));
    Span4Mux_h I__6690 (
            .O(N__28588),
            .I(N__28565));
    LocalMux I__6689 (
            .O(N__28585),
            .I(N__28565));
    LocalMux I__6688 (
            .O(N__28582),
            .I(N__28562));
    InMux I__6687 (
            .O(N__28579),
            .I(N__28559));
    CascadeMux I__6686 (
            .O(N__28578),
            .I(N__28556));
    InMux I__6685 (
            .O(N__28575),
            .I(N__28551));
    CascadeMux I__6684 (
            .O(N__28574),
            .I(N__28548));
    InMux I__6683 (
            .O(N__28571),
            .I(N__28544));
    CascadeMux I__6682 (
            .O(N__28570),
            .I(N__28541));
    Span4Mux_v I__6681 (
            .O(N__28565),
            .I(N__28533));
    Span4Mux_h I__6680 (
            .O(N__28562),
            .I(N__28533));
    LocalMux I__6679 (
            .O(N__28559),
            .I(N__28533));
    InMux I__6678 (
            .O(N__28556),
            .I(N__28530));
    CascadeMux I__6677 (
            .O(N__28555),
            .I(N__28527));
    CascadeMux I__6676 (
            .O(N__28554),
            .I(N__28524));
    LocalMux I__6675 (
            .O(N__28551),
            .I(N__28521));
    InMux I__6674 (
            .O(N__28548),
            .I(N__28518));
    CascadeMux I__6673 (
            .O(N__28547),
            .I(N__28515));
    LocalMux I__6672 (
            .O(N__28544),
            .I(N__28511));
    InMux I__6671 (
            .O(N__28541),
            .I(N__28508));
    CascadeMux I__6670 (
            .O(N__28540),
            .I(N__28505));
    Span4Mux_v I__6669 (
            .O(N__28533),
            .I(N__28501));
    LocalMux I__6668 (
            .O(N__28530),
            .I(N__28498));
    InMux I__6667 (
            .O(N__28527),
            .I(N__28495));
    InMux I__6666 (
            .O(N__28524),
            .I(N__28492));
    Span4Mux_v I__6665 (
            .O(N__28521),
            .I(N__28487));
    LocalMux I__6664 (
            .O(N__28518),
            .I(N__28487));
    InMux I__6663 (
            .O(N__28515),
            .I(N__28484));
    CascadeMux I__6662 (
            .O(N__28514),
            .I(N__28481));
    Span4Mux_s3_v I__6661 (
            .O(N__28511),
            .I(N__28476));
    LocalMux I__6660 (
            .O(N__28508),
            .I(N__28476));
    InMux I__6659 (
            .O(N__28505),
            .I(N__28473));
    CascadeMux I__6658 (
            .O(N__28504),
            .I(N__28470));
    Sp12to4 I__6657 (
            .O(N__28501),
            .I(N__28466));
    Sp12to4 I__6656 (
            .O(N__28498),
            .I(N__28463));
    LocalMux I__6655 (
            .O(N__28495),
            .I(N__28458));
    LocalMux I__6654 (
            .O(N__28492),
            .I(N__28458));
    Span4Mux_v I__6653 (
            .O(N__28487),
            .I(N__28453));
    LocalMux I__6652 (
            .O(N__28484),
            .I(N__28453));
    InMux I__6651 (
            .O(N__28481),
            .I(N__28450));
    Span4Mux_v I__6650 (
            .O(N__28476),
            .I(N__28445));
    LocalMux I__6649 (
            .O(N__28473),
            .I(N__28445));
    InMux I__6648 (
            .O(N__28470),
            .I(N__28442));
    CascadeMux I__6647 (
            .O(N__28469),
            .I(N__28439));
    Span12Mux_h I__6646 (
            .O(N__28466),
            .I(N__28436));
    Span12Mux_h I__6645 (
            .O(N__28463),
            .I(N__28433));
    Span4Mux_v I__6644 (
            .O(N__28458),
            .I(N__28426));
    Span4Mux_v I__6643 (
            .O(N__28453),
            .I(N__28426));
    LocalMux I__6642 (
            .O(N__28450),
            .I(N__28426));
    Span4Mux_v I__6641 (
            .O(N__28445),
            .I(N__28421));
    LocalMux I__6640 (
            .O(N__28442),
            .I(N__28421));
    InMux I__6639 (
            .O(N__28439),
            .I(N__28418));
    Odrv12 I__6638 (
            .O(N__28436),
            .I(M_this_ppu_sprites_addr_4));
    Odrv12 I__6637 (
            .O(N__28433),
            .I(M_this_ppu_sprites_addr_4));
    Odrv4 I__6636 (
            .O(N__28426),
            .I(M_this_ppu_sprites_addr_4));
    Odrv4 I__6635 (
            .O(N__28421),
            .I(M_this_ppu_sprites_addr_4));
    LocalMux I__6634 (
            .O(N__28418),
            .I(M_this_ppu_sprites_addr_4));
    InMux I__6633 (
            .O(N__28407),
            .I(N__28404));
    LocalMux I__6632 (
            .O(N__28404),
            .I(N__28401));
    Span4Mux_v I__6631 (
            .O(N__28401),
            .I(N__28398));
    Odrv4 I__6630 (
            .O(N__28398),
            .I(N_32_0));
    CascadeMux I__6629 (
            .O(N__28395),
            .I(N__28392));
    InMux I__6628 (
            .O(N__28392),
            .I(N__28389));
    LocalMux I__6627 (
            .O(N__28389),
            .I(N__28386));
    Odrv4 I__6626 (
            .O(N__28386),
            .I(M_this_data_tmp_qZ0Z_11));
    InMux I__6625 (
            .O(N__28383),
            .I(N__28380));
    LocalMux I__6624 (
            .O(N__28380),
            .I(N__28377));
    Odrv4 I__6623 (
            .O(N__28377),
            .I(M_this_oam_ram_write_data_11));
    CascadeMux I__6622 (
            .O(N__28374),
            .I(N__28371));
    InMux I__6621 (
            .O(N__28371),
            .I(N__28368));
    LocalMux I__6620 (
            .O(N__28368),
            .I(N__28365));
    Odrv4 I__6619 (
            .O(N__28365),
            .I(M_this_data_tmp_qZ0Z_0));
    InMux I__6618 (
            .O(N__28362),
            .I(N__28359));
    LocalMux I__6617 (
            .O(N__28359),
            .I(N__28356));
    Span4Mux_h I__6616 (
            .O(N__28356),
            .I(N__28353));
    Odrv4 I__6615 (
            .O(N__28353),
            .I(N_748_0));
    InMux I__6614 (
            .O(N__28350),
            .I(N__28347));
    LocalMux I__6613 (
            .O(N__28347),
            .I(N__28344));
    Span4Mux_v I__6612 (
            .O(N__28344),
            .I(N__28341));
    Odrv4 I__6611 (
            .O(N__28341),
            .I(N_44_0));
    CascadeMux I__6610 (
            .O(N__28338),
            .I(N__28335));
    InMux I__6609 (
            .O(N__28335),
            .I(N__28332));
    LocalMux I__6608 (
            .O(N__28332),
            .I(M_this_data_tmp_qZ0Z_17));
    CEMux I__6607 (
            .O(N__28329),
            .I(N__28322));
    CEMux I__6606 (
            .O(N__28328),
            .I(N__28319));
    CEMux I__6605 (
            .O(N__28327),
            .I(N__28316));
    CEMux I__6604 (
            .O(N__28326),
            .I(N__28313));
    CEMux I__6603 (
            .O(N__28325),
            .I(N__28310));
    LocalMux I__6602 (
            .O(N__28322),
            .I(N__28307));
    LocalMux I__6601 (
            .O(N__28319),
            .I(N__28304));
    LocalMux I__6600 (
            .O(N__28316),
            .I(N__28301));
    LocalMux I__6599 (
            .O(N__28313),
            .I(N__28298));
    LocalMux I__6598 (
            .O(N__28310),
            .I(N__28295));
    Span4Mux_v I__6597 (
            .O(N__28307),
            .I(N__28292));
    Span4Mux_v I__6596 (
            .O(N__28304),
            .I(N__28289));
    Span4Mux_v I__6595 (
            .O(N__28301),
            .I(N__28286));
    Span4Mux_h I__6594 (
            .O(N__28298),
            .I(N__28283));
    Span4Mux_v I__6593 (
            .O(N__28295),
            .I(N__28280));
    Odrv4 I__6592 (
            .O(N__28292),
            .I(N_1174_0));
    Odrv4 I__6591 (
            .O(N__28289),
            .I(N_1174_0));
    Odrv4 I__6590 (
            .O(N__28286),
            .I(N_1174_0));
    Odrv4 I__6589 (
            .O(N__28283),
            .I(N_1174_0));
    Odrv4 I__6588 (
            .O(N__28280),
            .I(N_1174_0));
    InMux I__6587 (
            .O(N__28269),
            .I(N__28266));
    LocalMux I__6586 (
            .O(N__28266),
            .I(N__28263));
    Odrv4 I__6585 (
            .O(N__28263),
            .I(M_this_data_tmp_qZ0Z_23));
    InMux I__6584 (
            .O(N__28260),
            .I(N__28257));
    LocalMux I__6583 (
            .O(N__28257),
            .I(N__28254));
    Span4Mux_h I__6582 (
            .O(N__28254),
            .I(N__28251));
    Odrv4 I__6581 (
            .O(N__28251),
            .I(M_this_oam_ram_write_data_23));
    CascadeMux I__6580 (
            .O(N__28248),
            .I(N__28245));
    InMux I__6579 (
            .O(N__28245),
            .I(N__28242));
    LocalMux I__6578 (
            .O(N__28242),
            .I(M_this_data_tmp_qZ0Z_20));
    InMux I__6577 (
            .O(N__28239),
            .I(N__28236));
    LocalMux I__6576 (
            .O(N__28236),
            .I(N__28233));
    Span4Mux_h I__6575 (
            .O(N__28233),
            .I(N__28230));
    Odrv4 I__6574 (
            .O(N__28230),
            .I(N_42_0));
    CascadeMux I__6573 (
            .O(N__28227),
            .I(N__28224));
    InMux I__6572 (
            .O(N__28224),
            .I(N__28221));
    LocalMux I__6571 (
            .O(N__28221),
            .I(M_this_data_tmp_qZ0Z_8));
    CEMux I__6570 (
            .O(N__28218),
            .I(N__28214));
    CEMux I__6569 (
            .O(N__28217),
            .I(N__28210));
    LocalMux I__6568 (
            .O(N__28214),
            .I(N__28207));
    CEMux I__6567 (
            .O(N__28213),
            .I(N__28204));
    LocalMux I__6566 (
            .O(N__28210),
            .I(N__28201));
    Span4Mux_v I__6565 (
            .O(N__28207),
            .I(N__28198));
    LocalMux I__6564 (
            .O(N__28204),
            .I(N__28195));
    Span4Mux_h I__6563 (
            .O(N__28201),
            .I(N__28192));
    Span4Mux_h I__6562 (
            .O(N__28198),
            .I(N__28187));
    Span4Mux_h I__6561 (
            .O(N__28195),
            .I(N__28187));
    Odrv4 I__6560 (
            .O(N__28192),
            .I(N_1182_0));
    Odrv4 I__6559 (
            .O(N__28187),
            .I(N_1182_0));
    CascadeMux I__6558 (
            .O(N__28182),
            .I(N__28179));
    InMux I__6557 (
            .O(N__28179),
            .I(N__28176));
    LocalMux I__6556 (
            .O(N__28176),
            .I(M_this_data_tmp_qZ0Z_3));
    InMux I__6555 (
            .O(N__28173),
            .I(N__28170));
    LocalMux I__6554 (
            .O(N__28170),
            .I(N__28167));
    Span4Mux_h I__6553 (
            .O(N__28167),
            .I(N__28164));
    Odrv4 I__6552 (
            .O(N__28164),
            .I(N_745_0));
    CascadeMux I__6551 (
            .O(N__28161),
            .I(N__28158));
    InMux I__6550 (
            .O(N__28158),
            .I(N__28155));
    LocalMux I__6549 (
            .O(N__28155),
            .I(N__28152));
    Odrv4 I__6548 (
            .O(N__28152),
            .I(M_this_data_tmp_qZ0Z_14));
    InMux I__6547 (
            .O(N__28149),
            .I(N__28146));
    LocalMux I__6546 (
            .O(N__28146),
            .I(N__28143));
    Span4Mux_h I__6545 (
            .O(N__28143),
            .I(N__28140));
    Odrv4 I__6544 (
            .O(N__28140),
            .I(N_739_0));
    CascadeMux I__6543 (
            .O(N__28137),
            .I(N__28134));
    InMux I__6542 (
            .O(N__28134),
            .I(N__28131));
    LocalMux I__6541 (
            .O(N__28131),
            .I(N__28128));
    Odrv4 I__6540 (
            .O(N__28128),
            .I(M_this_data_tmp_qZ0Z_5));
    InMux I__6539 (
            .O(N__28125),
            .I(N__28122));
    LocalMux I__6538 (
            .O(N__28122),
            .I(N__28119));
    Span4Mux_h I__6537 (
            .O(N__28119),
            .I(N__28116));
    Odrv4 I__6536 (
            .O(N__28116),
            .I(N_743_0));
    CascadeMux I__6535 (
            .O(N__28113),
            .I(N_101_cascade_));
    InMux I__6534 (
            .O(N__28110),
            .I(N__28107));
    LocalMux I__6533 (
            .O(N__28107),
            .I(N__28104));
    Odrv4 I__6532 (
            .O(N__28104),
            .I(M_this_sprites_address_q_RNO_0Z0Z_6));
    CascadeMux I__6531 (
            .O(N__28101),
            .I(N__28095));
    CascadeMux I__6530 (
            .O(N__28100),
            .I(N__28092));
    CascadeMux I__6529 (
            .O(N__28099),
            .I(N__28087));
    CascadeMux I__6528 (
            .O(N__28098),
            .I(N__28080));
    InMux I__6527 (
            .O(N__28095),
            .I(N__28075));
    InMux I__6526 (
            .O(N__28092),
            .I(N__28072));
    CascadeMux I__6525 (
            .O(N__28091),
            .I(N__28069));
    CascadeMux I__6524 (
            .O(N__28090),
            .I(N__28066));
    InMux I__6523 (
            .O(N__28087),
            .I(N__28061));
    CascadeMux I__6522 (
            .O(N__28086),
            .I(N__28058));
    CascadeMux I__6521 (
            .O(N__28085),
            .I(N__28055));
    CascadeMux I__6520 (
            .O(N__28084),
            .I(N__28052));
    CascadeMux I__6519 (
            .O(N__28083),
            .I(N__28049));
    InMux I__6518 (
            .O(N__28080),
            .I(N__28046));
    CascadeMux I__6517 (
            .O(N__28079),
            .I(N__28043));
    CascadeMux I__6516 (
            .O(N__28078),
            .I(N__28040));
    LocalMux I__6515 (
            .O(N__28075),
            .I(N__28036));
    LocalMux I__6514 (
            .O(N__28072),
            .I(N__28033));
    InMux I__6513 (
            .O(N__28069),
            .I(N__28030));
    InMux I__6512 (
            .O(N__28066),
            .I(N__28027));
    CascadeMux I__6511 (
            .O(N__28065),
            .I(N__28024));
    CascadeMux I__6510 (
            .O(N__28064),
            .I(N__28021));
    LocalMux I__6509 (
            .O(N__28061),
            .I(N__28017));
    InMux I__6508 (
            .O(N__28058),
            .I(N__28014));
    InMux I__6507 (
            .O(N__28055),
            .I(N__28011));
    InMux I__6506 (
            .O(N__28052),
            .I(N__28008));
    InMux I__6505 (
            .O(N__28049),
            .I(N__28005));
    LocalMux I__6504 (
            .O(N__28046),
            .I(N__28002));
    InMux I__6503 (
            .O(N__28043),
            .I(N__27999));
    InMux I__6502 (
            .O(N__28040),
            .I(N__27996));
    CascadeMux I__6501 (
            .O(N__28039),
            .I(N__27993));
    Span4Mux_v I__6500 (
            .O(N__28036),
            .I(N__27984));
    Span4Mux_v I__6499 (
            .O(N__28033),
            .I(N__27984));
    LocalMux I__6498 (
            .O(N__28030),
            .I(N__27984));
    LocalMux I__6497 (
            .O(N__28027),
            .I(N__27984));
    InMux I__6496 (
            .O(N__28024),
            .I(N__27981));
    InMux I__6495 (
            .O(N__28021),
            .I(N__27978));
    CascadeMux I__6494 (
            .O(N__28020),
            .I(N__27975));
    Span4Mux_v I__6493 (
            .O(N__28017),
            .I(N__27968));
    LocalMux I__6492 (
            .O(N__28014),
            .I(N__27968));
    LocalMux I__6491 (
            .O(N__28011),
            .I(N__27968));
    LocalMux I__6490 (
            .O(N__28008),
            .I(N__27963));
    LocalMux I__6489 (
            .O(N__28005),
            .I(N__27963));
    Span4Mux_v I__6488 (
            .O(N__28002),
            .I(N__27956));
    LocalMux I__6487 (
            .O(N__27999),
            .I(N__27956));
    LocalMux I__6486 (
            .O(N__27996),
            .I(N__27956));
    InMux I__6485 (
            .O(N__27993),
            .I(N__27953));
    Span4Mux_v I__6484 (
            .O(N__27984),
            .I(N__27946));
    LocalMux I__6483 (
            .O(N__27981),
            .I(N__27946));
    LocalMux I__6482 (
            .O(N__27978),
            .I(N__27946));
    InMux I__6481 (
            .O(N__27975),
            .I(N__27943));
    Span4Mux_v I__6480 (
            .O(N__27968),
            .I(N__27938));
    Span4Mux_v I__6479 (
            .O(N__27963),
            .I(N__27938));
    Span4Mux_v I__6478 (
            .O(N__27956),
            .I(N__27929));
    LocalMux I__6477 (
            .O(N__27953),
            .I(N__27929));
    Span4Mux_v I__6476 (
            .O(N__27946),
            .I(N__27929));
    LocalMux I__6475 (
            .O(N__27943),
            .I(N__27929));
    Sp12to4 I__6474 (
            .O(N__27938),
            .I(N__27925));
    Span4Mux_v I__6473 (
            .O(N__27929),
            .I(N__27922));
    InMux I__6472 (
            .O(N__27928),
            .I(N__27918));
    Span12Mux_h I__6471 (
            .O(N__27925),
            .I(N__27915));
    Sp12to4 I__6470 (
            .O(N__27922),
            .I(N__27912));
    InMux I__6469 (
            .O(N__27921),
            .I(N__27909));
    LocalMux I__6468 (
            .O(N__27918),
            .I(N__27906));
    Odrv12 I__6467 (
            .O(N__27915),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv12 I__6466 (
            .O(N__27912),
            .I(M_this_sprites_address_qZ0Z_6));
    LocalMux I__6465 (
            .O(N__27909),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv4 I__6464 (
            .O(N__27906),
            .I(M_this_sprites_address_qZ0Z_6));
    InMux I__6463 (
            .O(N__27897),
            .I(N__27894));
    LocalMux I__6462 (
            .O(N__27894),
            .I(\this_vga_signals.M_this_sprites_address_q_3_bmZ0Z_1 ));
    CascadeMux I__6461 (
            .O(N__27891),
            .I(N__27881));
    CascadeMux I__6460 (
            .O(N__27890),
            .I(N__27878));
    CascadeMux I__6459 (
            .O(N__27889),
            .I(N__27873));
    CascadeMux I__6458 (
            .O(N__27888),
            .I(N__27868));
    CascadeMux I__6457 (
            .O(N__27887),
            .I(N__27865));
    CascadeMux I__6456 (
            .O(N__27886),
            .I(N__27862));
    CascadeMux I__6455 (
            .O(N__27885),
            .I(N__27859));
    CascadeMux I__6454 (
            .O(N__27884),
            .I(N__27856));
    InMux I__6453 (
            .O(N__27881),
            .I(N__27852));
    InMux I__6452 (
            .O(N__27878),
            .I(N__27849));
    CascadeMux I__6451 (
            .O(N__27877),
            .I(N__27846));
    CascadeMux I__6450 (
            .O(N__27876),
            .I(N__27843));
    InMux I__6449 (
            .O(N__27873),
            .I(N__27839));
    CascadeMux I__6448 (
            .O(N__27872),
            .I(N__27836));
    CascadeMux I__6447 (
            .O(N__27871),
            .I(N__27833));
    InMux I__6446 (
            .O(N__27868),
            .I(N__27828));
    InMux I__6445 (
            .O(N__27865),
            .I(N__27825));
    InMux I__6444 (
            .O(N__27862),
            .I(N__27822));
    InMux I__6443 (
            .O(N__27859),
            .I(N__27819));
    InMux I__6442 (
            .O(N__27856),
            .I(N__27816));
    CascadeMux I__6441 (
            .O(N__27855),
            .I(N__27813));
    LocalMux I__6440 (
            .O(N__27852),
            .I(N__27810));
    LocalMux I__6439 (
            .O(N__27849),
            .I(N__27807));
    InMux I__6438 (
            .O(N__27846),
            .I(N__27804));
    InMux I__6437 (
            .O(N__27843),
            .I(N__27801));
    CascadeMux I__6436 (
            .O(N__27842),
            .I(N__27798));
    LocalMux I__6435 (
            .O(N__27839),
            .I(N__27795));
    InMux I__6434 (
            .O(N__27836),
            .I(N__27792));
    InMux I__6433 (
            .O(N__27833),
            .I(N__27789));
    CascadeMux I__6432 (
            .O(N__27832),
            .I(N__27786));
    CascadeMux I__6431 (
            .O(N__27831),
            .I(N__27783));
    LocalMux I__6430 (
            .O(N__27828),
            .I(N__27776));
    LocalMux I__6429 (
            .O(N__27825),
            .I(N__27776));
    LocalMux I__6428 (
            .O(N__27822),
            .I(N__27776));
    LocalMux I__6427 (
            .O(N__27819),
            .I(N__27771));
    LocalMux I__6426 (
            .O(N__27816),
            .I(N__27771));
    InMux I__6425 (
            .O(N__27813),
            .I(N__27767));
    Span4Mux_v I__6424 (
            .O(N__27810),
            .I(N__27757));
    Span4Mux_v I__6423 (
            .O(N__27807),
            .I(N__27757));
    LocalMux I__6422 (
            .O(N__27804),
            .I(N__27757));
    LocalMux I__6421 (
            .O(N__27801),
            .I(N__27757));
    InMux I__6420 (
            .O(N__27798),
            .I(N__27754));
    Span4Mux_v I__6419 (
            .O(N__27795),
            .I(N__27747));
    LocalMux I__6418 (
            .O(N__27792),
            .I(N__27747));
    LocalMux I__6417 (
            .O(N__27789),
            .I(N__27747));
    InMux I__6416 (
            .O(N__27786),
            .I(N__27744));
    InMux I__6415 (
            .O(N__27783),
            .I(N__27741));
    Span12Mux_v I__6414 (
            .O(N__27776),
            .I(N__27735));
    Span12Mux_v I__6413 (
            .O(N__27771),
            .I(N__27735));
    CascadeMux I__6412 (
            .O(N__27770),
            .I(N__27732));
    LocalMux I__6411 (
            .O(N__27767),
            .I(N__27729));
    InMux I__6410 (
            .O(N__27766),
            .I(N__27726));
    Span4Mux_v I__6409 (
            .O(N__27757),
            .I(N__27721));
    LocalMux I__6408 (
            .O(N__27754),
            .I(N__27721));
    Span4Mux_v I__6407 (
            .O(N__27747),
            .I(N__27714));
    LocalMux I__6406 (
            .O(N__27744),
            .I(N__27714));
    LocalMux I__6405 (
            .O(N__27741),
            .I(N__27714));
    InMux I__6404 (
            .O(N__27740),
            .I(N__27711));
    Span12Mux_h I__6403 (
            .O(N__27735),
            .I(N__27708));
    InMux I__6402 (
            .O(N__27732),
            .I(N__27705));
    Span4Mux_h I__6401 (
            .O(N__27729),
            .I(N__27700));
    LocalMux I__6400 (
            .O(N__27726),
            .I(N__27700));
    Span4Mux_v I__6399 (
            .O(N__27721),
            .I(N__27693));
    Span4Mux_v I__6398 (
            .O(N__27714),
            .I(N__27693));
    LocalMux I__6397 (
            .O(N__27711),
            .I(N__27693));
    Odrv12 I__6396 (
            .O(N__27708),
            .I(M_this_sprites_address_qZ0Z_1));
    LocalMux I__6395 (
            .O(N__27705),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv4 I__6394 (
            .O(N__27700),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv4 I__6393 (
            .O(N__27693),
            .I(M_this_sprites_address_qZ0Z_1));
    InMux I__6392 (
            .O(N__27684),
            .I(N__27673));
    InMux I__6391 (
            .O(N__27683),
            .I(N__27670));
    InMux I__6390 (
            .O(N__27682),
            .I(N__27663));
    InMux I__6389 (
            .O(N__27681),
            .I(N__27658));
    InMux I__6388 (
            .O(N__27680),
            .I(N__27658));
    InMux I__6387 (
            .O(N__27679),
            .I(N__27653));
    InMux I__6386 (
            .O(N__27678),
            .I(N__27653));
    InMux I__6385 (
            .O(N__27677),
            .I(N__27648));
    InMux I__6384 (
            .O(N__27676),
            .I(N__27648));
    LocalMux I__6383 (
            .O(N__27673),
            .I(N__27643));
    LocalMux I__6382 (
            .O(N__27670),
            .I(N__27643));
    InMux I__6381 (
            .O(N__27669),
            .I(N__27640));
    InMux I__6380 (
            .O(N__27668),
            .I(N__27637));
    CascadeMux I__6379 (
            .O(N__27667),
            .I(N__27633));
    CascadeMux I__6378 (
            .O(N__27666),
            .I(N__27629));
    LocalMux I__6377 (
            .O(N__27663),
            .I(N__27626));
    LocalMux I__6376 (
            .O(N__27658),
            .I(N__27622));
    LocalMux I__6375 (
            .O(N__27653),
            .I(N__27611));
    LocalMux I__6374 (
            .O(N__27648),
            .I(N__27611));
    Span4Mux_v I__6373 (
            .O(N__27643),
            .I(N__27611));
    LocalMux I__6372 (
            .O(N__27640),
            .I(N__27611));
    LocalMux I__6371 (
            .O(N__27637),
            .I(N__27611));
    InMux I__6370 (
            .O(N__27636),
            .I(N__27608));
    InMux I__6369 (
            .O(N__27633),
            .I(N__27604));
    InMux I__6368 (
            .O(N__27632),
            .I(N__27601));
    InMux I__6367 (
            .O(N__27629),
            .I(N__27598));
    Span4Mux_v I__6366 (
            .O(N__27626),
            .I(N__27595));
    InMux I__6365 (
            .O(N__27625),
            .I(N__27592));
    Span4Mux_v I__6364 (
            .O(N__27622),
            .I(N__27585));
    Span4Mux_h I__6363 (
            .O(N__27611),
            .I(N__27585));
    LocalMux I__6362 (
            .O(N__27608),
            .I(N__27585));
    InMux I__6361 (
            .O(N__27607),
            .I(N__27581));
    LocalMux I__6360 (
            .O(N__27604),
            .I(N__27570));
    LocalMux I__6359 (
            .O(N__27601),
            .I(N__27570));
    LocalMux I__6358 (
            .O(N__27598),
            .I(N__27570));
    Sp12to4 I__6357 (
            .O(N__27595),
            .I(N__27570));
    LocalMux I__6356 (
            .O(N__27592),
            .I(N__27570));
    Span4Mux_h I__6355 (
            .O(N__27585),
            .I(N__27567));
    InMux I__6354 (
            .O(N__27584),
            .I(N__27564));
    LocalMux I__6353 (
            .O(N__27581),
            .I(M_this_state_qZ0Z_2));
    Odrv12 I__6352 (
            .O(N__27570),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__6351 (
            .O(N__27567),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__6350 (
            .O(N__27564),
            .I(M_this_state_qZ0Z_2));
    InMux I__6349 (
            .O(N__27555),
            .I(N__27539));
    InMux I__6348 (
            .O(N__27554),
            .I(N__27533));
    InMux I__6347 (
            .O(N__27553),
            .I(N__27528));
    InMux I__6346 (
            .O(N__27552),
            .I(N__27528));
    InMux I__6345 (
            .O(N__27551),
            .I(N__27522));
    InMux I__6344 (
            .O(N__27550),
            .I(N__27522));
    InMux I__6343 (
            .O(N__27549),
            .I(N__27515));
    InMux I__6342 (
            .O(N__27548),
            .I(N__27511));
    InMux I__6341 (
            .O(N__27547),
            .I(N__27506));
    InMux I__6340 (
            .O(N__27546),
            .I(N__27506));
    InMux I__6339 (
            .O(N__27545),
            .I(N__27498));
    InMux I__6338 (
            .O(N__27544),
            .I(N__27498));
    InMux I__6337 (
            .O(N__27543),
            .I(N__27493));
    InMux I__6336 (
            .O(N__27542),
            .I(N__27493));
    LocalMux I__6335 (
            .O(N__27539),
            .I(N__27490));
    InMux I__6334 (
            .O(N__27538),
            .I(N__27487));
    InMux I__6333 (
            .O(N__27537),
            .I(N__27484));
    InMux I__6332 (
            .O(N__27536),
            .I(N__27481));
    LocalMux I__6331 (
            .O(N__27533),
            .I(N__27478));
    LocalMux I__6330 (
            .O(N__27528),
            .I(N__27475));
    InMux I__6329 (
            .O(N__27527),
            .I(N__27472));
    LocalMux I__6328 (
            .O(N__27522),
            .I(N__27469));
    InMux I__6327 (
            .O(N__27521),
            .I(N__27466));
    InMux I__6326 (
            .O(N__27520),
            .I(N__27461));
    InMux I__6325 (
            .O(N__27519),
            .I(N__27461));
    InMux I__6324 (
            .O(N__27518),
            .I(N__27454));
    LocalMux I__6323 (
            .O(N__27515),
            .I(N__27451));
    InMux I__6322 (
            .O(N__27514),
            .I(N__27448));
    LocalMux I__6321 (
            .O(N__27511),
            .I(N__27443));
    LocalMux I__6320 (
            .O(N__27506),
            .I(N__27443));
    InMux I__6319 (
            .O(N__27505),
            .I(N__27440));
    InMux I__6318 (
            .O(N__27504),
            .I(N__27435));
    InMux I__6317 (
            .O(N__27503),
            .I(N__27435));
    LocalMux I__6316 (
            .O(N__27498),
            .I(N__27426));
    LocalMux I__6315 (
            .O(N__27493),
            .I(N__27426));
    Span4Mux_v I__6314 (
            .O(N__27490),
            .I(N__27426));
    LocalMux I__6313 (
            .O(N__27487),
            .I(N__27426));
    LocalMux I__6312 (
            .O(N__27484),
            .I(N__27423));
    LocalMux I__6311 (
            .O(N__27481),
            .I(N__27420));
    Span4Mux_h I__6310 (
            .O(N__27478),
            .I(N__27409));
    Span4Mux_v I__6309 (
            .O(N__27475),
            .I(N__27409));
    LocalMux I__6308 (
            .O(N__27472),
            .I(N__27409));
    Span4Mux_v I__6307 (
            .O(N__27469),
            .I(N__27406));
    LocalMux I__6306 (
            .O(N__27466),
            .I(N__27401));
    LocalMux I__6305 (
            .O(N__27461),
            .I(N__27401));
    InMux I__6304 (
            .O(N__27460),
            .I(N__27394));
    InMux I__6303 (
            .O(N__27459),
            .I(N__27394));
    InMux I__6302 (
            .O(N__27458),
            .I(N__27394));
    InMux I__6301 (
            .O(N__27457),
            .I(N__27391));
    LocalMux I__6300 (
            .O(N__27454),
            .I(N__27378));
    Span4Mux_h I__6299 (
            .O(N__27451),
            .I(N__27378));
    LocalMux I__6298 (
            .O(N__27448),
            .I(N__27378));
    Span4Mux_h I__6297 (
            .O(N__27443),
            .I(N__27378));
    LocalMux I__6296 (
            .O(N__27440),
            .I(N__27378));
    LocalMux I__6295 (
            .O(N__27435),
            .I(N__27378));
    Span4Mux_h I__6294 (
            .O(N__27426),
            .I(N__27371));
    Span4Mux_h I__6293 (
            .O(N__27423),
            .I(N__27371));
    Span4Mux_h I__6292 (
            .O(N__27420),
            .I(N__27371));
    InMux I__6291 (
            .O(N__27419),
            .I(N__27362));
    InMux I__6290 (
            .O(N__27418),
            .I(N__27362));
    InMux I__6289 (
            .O(N__27417),
            .I(N__27362));
    InMux I__6288 (
            .O(N__27416),
            .I(N__27362));
    Odrv4 I__6287 (
            .O(N__27409),
            .I(N_87_0));
    Odrv4 I__6286 (
            .O(N__27406),
            .I(N_87_0));
    Odrv12 I__6285 (
            .O(N__27401),
            .I(N_87_0));
    LocalMux I__6284 (
            .O(N__27394),
            .I(N_87_0));
    LocalMux I__6283 (
            .O(N__27391),
            .I(N_87_0));
    Odrv4 I__6282 (
            .O(N__27378),
            .I(N_87_0));
    Odrv4 I__6281 (
            .O(N__27371),
            .I(N_87_0));
    LocalMux I__6280 (
            .O(N__27362),
            .I(N_87_0));
    InMux I__6279 (
            .O(N__27345),
            .I(N__27342));
    LocalMux I__6278 (
            .O(N__27342),
            .I(N__27339));
    Odrv4 I__6277 (
            .O(N__27339),
            .I(\this_vga_signals.M_this_sprites_address_q_3_amZ0Z_1 ));
    InMux I__6276 (
            .O(N__27336),
            .I(N__27333));
    LocalMux I__6275 (
            .O(N__27333),
            .I(N__27330));
    Span4Mux_h I__6274 (
            .O(N__27330),
            .I(N__27324));
    InMux I__6273 (
            .O(N__27329),
            .I(N__27319));
    InMux I__6272 (
            .O(N__27328),
            .I(N__27319));
    InMux I__6271 (
            .O(N__27327),
            .I(N__27316));
    Odrv4 I__6270 (
            .O(N__27324),
            .I(\this_vga_signals.un1_M_this_state_q_3_0_i_0_0 ));
    LocalMux I__6269 (
            .O(N__27319),
            .I(\this_vga_signals.un1_M_this_state_q_3_0_i_0_0 ));
    LocalMux I__6268 (
            .O(N__27316),
            .I(\this_vga_signals.un1_M_this_state_q_3_0_i_0_0 ));
    InMux I__6267 (
            .O(N__27309),
            .I(N__27306));
    LocalMux I__6266 (
            .O(N__27306),
            .I(N__27302));
    InMux I__6265 (
            .O(N__27305),
            .I(N__27299));
    Span4Mux_h I__6264 (
            .O(N__27302),
            .I(N__27293));
    LocalMux I__6263 (
            .O(N__27299),
            .I(N__27290));
    InMux I__6262 (
            .O(N__27298),
            .I(N__27283));
    InMux I__6261 (
            .O(N__27297),
            .I(N__27283));
    InMux I__6260 (
            .O(N__27296),
            .I(N__27283));
    Odrv4 I__6259 (
            .O(N__27293),
            .I(\this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2 ));
    Odrv4 I__6258 (
            .O(N__27290),
            .I(\this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2 ));
    LocalMux I__6257 (
            .O(N__27283),
            .I(\this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2 ));
    InMux I__6256 (
            .O(N__27276),
            .I(N__27270));
    InMux I__6255 (
            .O(N__27275),
            .I(N__27266));
    InMux I__6254 (
            .O(N__27274),
            .I(N__27263));
    InMux I__6253 (
            .O(N__27273),
            .I(N__27259));
    LocalMux I__6252 (
            .O(N__27270),
            .I(N__27256));
    InMux I__6251 (
            .O(N__27269),
            .I(N__27253));
    LocalMux I__6250 (
            .O(N__27266),
            .I(N__27246));
    LocalMux I__6249 (
            .O(N__27263),
            .I(N__27246));
    InMux I__6248 (
            .O(N__27262),
            .I(N__27243));
    LocalMux I__6247 (
            .O(N__27259),
            .I(N__27240));
    Span4Mux_h I__6246 (
            .O(N__27256),
            .I(N__27237));
    LocalMux I__6245 (
            .O(N__27253),
            .I(N__27234));
    InMux I__6244 (
            .O(N__27252),
            .I(N__27231));
    InMux I__6243 (
            .O(N__27251),
            .I(N__27228));
    Span12Mux_v I__6242 (
            .O(N__27246),
            .I(N__27223));
    LocalMux I__6241 (
            .O(N__27243),
            .I(N__27223));
    Span12Mux_h I__6240 (
            .O(N__27240),
            .I(N__27220));
    Span4Mux_v I__6239 (
            .O(N__27237),
            .I(N__27217));
    Span4Mux_h I__6238 (
            .O(N__27234),
            .I(N__27214));
    LocalMux I__6237 (
            .O(N__27231),
            .I(N__27211));
    LocalMux I__6236 (
            .O(N__27228),
            .I(N__27208));
    Span12Mux_h I__6235 (
            .O(N__27223),
            .I(N__27203));
    Span12Mux_v I__6234 (
            .O(N__27220),
            .I(N__27203));
    Span4Mux_v I__6233 (
            .O(N__27217),
            .I(N__27200));
    Span4Mux_v I__6232 (
            .O(N__27214),
            .I(N__27193));
    Span4Mux_h I__6231 (
            .O(N__27211),
            .I(N__27193));
    Span4Mux_h I__6230 (
            .O(N__27208),
            .I(N__27193));
    Odrv12 I__6229 (
            .O(N__27203),
            .I(M_this_sprites_ram_write_data_iv_i_i_3));
    Odrv4 I__6228 (
            .O(N__27200),
            .I(M_this_sprites_ram_write_data_iv_i_i_3));
    Odrv4 I__6227 (
            .O(N__27193),
            .I(M_this_sprites_ram_write_data_iv_i_i_3));
    InMux I__6226 (
            .O(N__27186),
            .I(N__27183));
    LocalMux I__6225 (
            .O(N__27183),
            .I(\this_ppu.un2_vscroll_axb_0 ));
    CascadeMux I__6224 (
            .O(N__27180),
            .I(N__27176));
    CascadeMux I__6223 (
            .O(N__27179),
            .I(N__27173));
    InMux I__6222 (
            .O(N__27176),
            .I(N__27168));
    InMux I__6221 (
            .O(N__27173),
            .I(N__27165));
    CascadeMux I__6220 (
            .O(N__27172),
            .I(N__27162));
    CascadeMux I__6219 (
            .O(N__27171),
            .I(N__27156));
    LocalMux I__6218 (
            .O(N__27168),
            .I(N__27151));
    LocalMux I__6217 (
            .O(N__27165),
            .I(N__27151));
    InMux I__6216 (
            .O(N__27162),
            .I(N__27148));
    CascadeMux I__6215 (
            .O(N__27161),
            .I(N__27145));
    CascadeMux I__6214 (
            .O(N__27160),
            .I(N__27141));
    CascadeMux I__6213 (
            .O(N__27159),
            .I(N__27138));
    InMux I__6212 (
            .O(N__27156),
            .I(N__27134));
    Span4Mux_s2_v I__6211 (
            .O(N__27151),
            .I(N__27129));
    LocalMux I__6210 (
            .O(N__27148),
            .I(N__27129));
    InMux I__6209 (
            .O(N__27145),
            .I(N__27126));
    CascadeMux I__6208 (
            .O(N__27144),
            .I(N__27123));
    InMux I__6207 (
            .O(N__27141),
            .I(N__27119));
    InMux I__6206 (
            .O(N__27138),
            .I(N__27116));
    CascadeMux I__6205 (
            .O(N__27137),
            .I(N__27113));
    LocalMux I__6204 (
            .O(N__27134),
            .I(N__27110));
    Span4Mux_v I__6203 (
            .O(N__27129),
            .I(N__27105));
    LocalMux I__6202 (
            .O(N__27126),
            .I(N__27105));
    InMux I__6201 (
            .O(N__27123),
            .I(N__27102));
    CascadeMux I__6200 (
            .O(N__27122),
            .I(N__27099));
    LocalMux I__6199 (
            .O(N__27119),
            .I(N__27094));
    LocalMux I__6198 (
            .O(N__27116),
            .I(N__27091));
    InMux I__6197 (
            .O(N__27113),
            .I(N__27088));
    Span4Mux_h I__6196 (
            .O(N__27110),
            .I(N__27085));
    Span4Mux_h I__6195 (
            .O(N__27105),
            .I(N__27080));
    LocalMux I__6194 (
            .O(N__27102),
            .I(N__27080));
    InMux I__6193 (
            .O(N__27099),
            .I(N__27077));
    CascadeMux I__6192 (
            .O(N__27098),
            .I(N__27074));
    CascadeMux I__6191 (
            .O(N__27097),
            .I(N__27070));
    Span4Mux_h I__6190 (
            .O(N__27094),
            .I(N__27067));
    Span4Mux_v I__6189 (
            .O(N__27091),
            .I(N__27062));
    LocalMux I__6188 (
            .O(N__27088),
            .I(N__27062));
    Span4Mux_h I__6187 (
            .O(N__27085),
            .I(N__27058));
    Span4Mux_v I__6186 (
            .O(N__27080),
            .I(N__27053));
    LocalMux I__6185 (
            .O(N__27077),
            .I(N__27053));
    InMux I__6184 (
            .O(N__27074),
            .I(N__27050));
    CascadeMux I__6183 (
            .O(N__27073),
            .I(N__27047));
    InMux I__6182 (
            .O(N__27070),
            .I(N__27043));
    Span4Mux_v I__6181 (
            .O(N__27067),
            .I(N__27038));
    Span4Mux_h I__6180 (
            .O(N__27062),
            .I(N__27038));
    CascadeMux I__6179 (
            .O(N__27061),
            .I(N__27035));
    Span4Mux_h I__6178 (
            .O(N__27058),
            .I(N__27032));
    Span4Mux_h I__6177 (
            .O(N__27053),
            .I(N__27027));
    LocalMux I__6176 (
            .O(N__27050),
            .I(N__27027));
    InMux I__6175 (
            .O(N__27047),
            .I(N__27024));
    CascadeMux I__6174 (
            .O(N__27046),
            .I(N__27021));
    LocalMux I__6173 (
            .O(N__27043),
            .I(N__27017));
    Span4Mux_v I__6172 (
            .O(N__27038),
            .I(N__27014));
    InMux I__6171 (
            .O(N__27035),
            .I(N__27011));
    Span4Mux_h I__6170 (
            .O(N__27032),
            .I(N__27004));
    Span4Mux_v I__6169 (
            .O(N__27027),
            .I(N__27004));
    LocalMux I__6168 (
            .O(N__27024),
            .I(N__27004));
    InMux I__6167 (
            .O(N__27021),
            .I(N__27001));
    CascadeMux I__6166 (
            .O(N__27020),
            .I(N__26998));
    Span12Mux_h I__6165 (
            .O(N__27017),
            .I(N__26995));
    Sp12to4 I__6164 (
            .O(N__27014),
            .I(N__26992));
    LocalMux I__6163 (
            .O(N__27011),
            .I(N__26989));
    Span4Mux_h I__6162 (
            .O(N__27004),
            .I(N__26984));
    LocalMux I__6161 (
            .O(N__27001),
            .I(N__26984));
    InMux I__6160 (
            .O(N__26998),
            .I(N__26981));
    Span12Mux_v I__6159 (
            .O(N__26995),
            .I(N__26978));
    Span12Mux_h I__6158 (
            .O(N__26992),
            .I(N__26975));
    Span4Mux_v I__6157 (
            .O(N__26989),
            .I(N__26968));
    Span4Mux_v I__6156 (
            .O(N__26984),
            .I(N__26968));
    LocalMux I__6155 (
            .O(N__26981),
            .I(N__26968));
    Odrv12 I__6154 (
            .O(N__26978),
            .I(M_this_ppu_sprites_addr_1));
    Odrv12 I__6153 (
            .O(N__26975),
            .I(M_this_ppu_sprites_addr_1));
    Odrv4 I__6152 (
            .O(N__26968),
            .I(M_this_ppu_sprites_addr_1));
    CascadeMux I__6151 (
            .O(N__26961),
            .I(N__26958));
    InMux I__6150 (
            .O(N__26958),
            .I(N__26955));
    LocalMux I__6149 (
            .O(N__26955),
            .I(M_this_data_tmp_qZ0Z_4));
    InMux I__6148 (
            .O(N__26952),
            .I(N__26949));
    LocalMux I__6147 (
            .O(N__26949),
            .I(N__26946));
    Span4Mux_v I__6146 (
            .O(N__26946),
            .I(N__26943));
    Odrv4 I__6145 (
            .O(N__26943),
            .I(N_744_0));
    InMux I__6144 (
            .O(N__26940),
            .I(N__26937));
    LocalMux I__6143 (
            .O(N__26937),
            .I(N__26934));
    Odrv4 I__6142 (
            .O(N__26934),
            .I(M_this_data_tmp_qZ0Z_7));
    InMux I__6141 (
            .O(N__26931),
            .I(N__26928));
    LocalMux I__6140 (
            .O(N__26928),
            .I(N__26925));
    Span4Mux_h I__6139 (
            .O(N__26925),
            .I(N__26922));
    Odrv4 I__6138 (
            .O(N__26922),
            .I(N_56_0));
    CascadeMux I__6137 (
            .O(N__26919),
            .I(N__26916));
    InMux I__6136 (
            .O(N__26916),
            .I(N__26913));
    LocalMux I__6135 (
            .O(N__26913),
            .I(M_this_data_tmp_qZ0Z_16));
    InMux I__6134 (
            .O(N__26910),
            .I(N__26907));
    LocalMux I__6133 (
            .O(N__26907),
            .I(N__26904));
    Span4Mux_h I__6132 (
            .O(N__26904),
            .I(N__26901));
    Odrv4 I__6131 (
            .O(N__26901),
            .I(N_738_0));
    CascadeMux I__6130 (
            .O(N__26898),
            .I(N__26895));
    InMux I__6129 (
            .O(N__26895),
            .I(N__26892));
    LocalMux I__6128 (
            .O(N__26892),
            .I(M_this_data_tmp_qZ0Z_22));
    InMux I__6127 (
            .O(N__26889),
            .I(N__26886));
    LocalMux I__6126 (
            .O(N__26886),
            .I(N__26883));
    Span4Mux_h I__6125 (
            .O(N__26883),
            .I(N__26880));
    Odrv4 I__6124 (
            .O(N__26880),
            .I(N_40_0));
    InMux I__6123 (
            .O(N__26877),
            .I(N__26874));
    LocalMux I__6122 (
            .O(N__26874),
            .I(N__26871));
    Span4Mux_h I__6121 (
            .O(N__26871),
            .I(N__26868));
    Span4Mux_v I__6120 (
            .O(N__26868),
            .I(N__26865));
    Odrv4 I__6119 (
            .O(N__26865),
            .I(\this_sprites_ram.mem_out_bus6_0 ));
    InMux I__6118 (
            .O(N__26862),
            .I(N__26859));
    LocalMux I__6117 (
            .O(N__26859),
            .I(N__26856));
    Span4Mux_v I__6116 (
            .O(N__26856),
            .I(N__26853));
    Odrv4 I__6115 (
            .O(N__26853),
            .I(\this_sprites_ram.mem_out_bus2_0 ));
    InMux I__6114 (
            .O(N__26850),
            .I(N__26847));
    LocalMux I__6113 (
            .O(N__26847),
            .I(N__26844));
    Odrv12 I__6112 (
            .O(N__26844),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ));
    CascadeMux I__6111 (
            .O(N__26841),
            .I(N__26838));
    InMux I__6110 (
            .O(N__26838),
            .I(N__26835));
    LocalMux I__6109 (
            .O(N__26835),
            .I(N_102));
    InMux I__6108 (
            .O(N__26832),
            .I(N__26829));
    LocalMux I__6107 (
            .O(N__26829),
            .I(N__26826));
    Odrv4 I__6106 (
            .O(N__26826),
            .I(M_this_sprites_address_q_RNO_0Z0Z_4));
    CascadeMux I__6105 (
            .O(N__26823),
            .I(N__26817));
    CascadeMux I__6104 (
            .O(N__26822),
            .I(N__26812));
    CascadeMux I__6103 (
            .O(N__26821),
            .I(N__26805));
    CascadeMux I__6102 (
            .O(N__26820),
            .I(N__26802));
    InMux I__6101 (
            .O(N__26817),
            .I(N__26797));
    CascadeMux I__6100 (
            .O(N__26816),
            .I(N__26794));
    CascadeMux I__6099 (
            .O(N__26815),
            .I(N__26791));
    InMux I__6098 (
            .O(N__26812),
            .I(N__26787));
    CascadeMux I__6097 (
            .O(N__26811),
            .I(N__26784));
    CascadeMux I__6096 (
            .O(N__26810),
            .I(N__26781));
    CascadeMux I__6095 (
            .O(N__26809),
            .I(N__26778));
    CascadeMux I__6094 (
            .O(N__26808),
            .I(N__26775));
    InMux I__6093 (
            .O(N__26805),
            .I(N__26772));
    InMux I__6092 (
            .O(N__26802),
            .I(N__26769));
    CascadeMux I__6091 (
            .O(N__26801),
            .I(N__26766));
    CascadeMux I__6090 (
            .O(N__26800),
            .I(N__26763));
    LocalMux I__6089 (
            .O(N__26797),
            .I(N__26760));
    InMux I__6088 (
            .O(N__26794),
            .I(N__26757));
    InMux I__6087 (
            .O(N__26791),
            .I(N__26754));
    CascadeMux I__6086 (
            .O(N__26790),
            .I(N__26751));
    LocalMux I__6085 (
            .O(N__26787),
            .I(N__26745));
    InMux I__6084 (
            .O(N__26784),
            .I(N__26742));
    InMux I__6083 (
            .O(N__26781),
            .I(N__26739));
    InMux I__6082 (
            .O(N__26778),
            .I(N__26736));
    InMux I__6081 (
            .O(N__26775),
            .I(N__26733));
    LocalMux I__6080 (
            .O(N__26772),
            .I(N__26728));
    LocalMux I__6079 (
            .O(N__26769),
            .I(N__26728));
    InMux I__6078 (
            .O(N__26766),
            .I(N__26725));
    InMux I__6077 (
            .O(N__26763),
            .I(N__26722));
    Span4Mux_v I__6076 (
            .O(N__26760),
            .I(N__26715));
    LocalMux I__6075 (
            .O(N__26757),
            .I(N__26715));
    LocalMux I__6074 (
            .O(N__26754),
            .I(N__26715));
    InMux I__6073 (
            .O(N__26751),
            .I(N__26712));
    CascadeMux I__6072 (
            .O(N__26750),
            .I(N__26709));
    CascadeMux I__6071 (
            .O(N__26749),
            .I(N__26706));
    CascadeMux I__6070 (
            .O(N__26748),
            .I(N__26703));
    Span4Mux_v I__6069 (
            .O(N__26745),
            .I(N__26698));
    LocalMux I__6068 (
            .O(N__26742),
            .I(N__26698));
    LocalMux I__6067 (
            .O(N__26739),
            .I(N__26695));
    LocalMux I__6066 (
            .O(N__26736),
            .I(N__26690));
    LocalMux I__6065 (
            .O(N__26733),
            .I(N__26690));
    Span4Mux_v I__6064 (
            .O(N__26728),
            .I(N__26683));
    LocalMux I__6063 (
            .O(N__26725),
            .I(N__26683));
    LocalMux I__6062 (
            .O(N__26722),
            .I(N__26683));
    Span4Mux_v I__6061 (
            .O(N__26715),
            .I(N__26678));
    LocalMux I__6060 (
            .O(N__26712),
            .I(N__26678));
    InMux I__6059 (
            .O(N__26709),
            .I(N__26675));
    InMux I__6058 (
            .O(N__26706),
            .I(N__26672));
    InMux I__6057 (
            .O(N__26703),
            .I(N__26669));
    Span4Mux_v I__6056 (
            .O(N__26698),
            .I(N__26662));
    Span4Mux_v I__6055 (
            .O(N__26695),
            .I(N__26662));
    Span4Mux_v I__6054 (
            .O(N__26690),
            .I(N__26662));
    Span4Mux_v I__6053 (
            .O(N__26683),
            .I(N__26655));
    Span4Mux_v I__6052 (
            .O(N__26678),
            .I(N__26655));
    LocalMux I__6051 (
            .O(N__26675),
            .I(N__26655));
    LocalMux I__6050 (
            .O(N__26672),
            .I(N__26651));
    LocalMux I__6049 (
            .O(N__26669),
            .I(N__26648));
    Sp12to4 I__6048 (
            .O(N__26662),
            .I(N__26644));
    Span4Mux_v I__6047 (
            .O(N__26655),
            .I(N__26641));
    InMux I__6046 (
            .O(N__26654),
            .I(N__26638));
    Span4Mux_h I__6045 (
            .O(N__26651),
            .I(N__26633));
    Span4Mux_h I__6044 (
            .O(N__26648),
            .I(N__26633));
    InMux I__6043 (
            .O(N__26647),
            .I(N__26630));
    Span12Mux_h I__6042 (
            .O(N__26644),
            .I(N__26623));
    Sp12to4 I__6041 (
            .O(N__26641),
            .I(N__26623));
    LocalMux I__6040 (
            .O(N__26638),
            .I(N__26623));
    Odrv4 I__6039 (
            .O(N__26633),
            .I(M_this_sprites_address_qZ0Z_4));
    LocalMux I__6038 (
            .O(N__26630),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv12 I__6037 (
            .O(N__26623),
            .I(M_this_sprites_address_qZ0Z_4));
    InMux I__6036 (
            .O(N__26616),
            .I(N__26613));
    LocalMux I__6035 (
            .O(N__26613),
            .I(N__26610));
    Span4Mux_h I__6034 (
            .O(N__26610),
            .I(N__26607));
    Sp12to4 I__6033 (
            .O(N__26607),
            .I(N__26604));
    Span12Mux_v I__6032 (
            .O(N__26604),
            .I(N__26601));
    Odrv12 I__6031 (
            .O(N__26601),
            .I(port_address_in_3));
    InMux I__6030 (
            .O(N__26598),
            .I(N__26595));
    LocalMux I__6029 (
            .O(N__26595),
            .I(N__26592));
    Span12Mux_v I__6028 (
            .O(N__26592),
            .I(N__26589));
    Odrv12 I__6027 (
            .O(N__26589),
            .I(port_address_in_2));
    CascadeMux I__6026 (
            .O(N__26586),
            .I(N__26583));
    InMux I__6025 (
            .O(N__26583),
            .I(N__26580));
    LocalMux I__6024 (
            .O(N__26580),
            .I(N__26577));
    Span4Mux_v I__6023 (
            .O(N__26577),
            .I(N__26574));
    Span4Mux_h I__6022 (
            .O(N__26574),
            .I(N__26571));
    Sp12to4 I__6021 (
            .O(N__26571),
            .I(N__26568));
    Span12Mux_h I__6020 (
            .O(N__26568),
            .I(N__26564));
    InMux I__6019 (
            .O(N__26567),
            .I(N__26561));
    Odrv12 I__6018 (
            .O(N__26564),
            .I(port_rw_in));
    LocalMux I__6017 (
            .O(N__26561),
            .I(port_rw_in));
    InMux I__6016 (
            .O(N__26556),
            .I(N__26553));
    LocalMux I__6015 (
            .O(N__26553),
            .I(N__26550));
    Span4Mux_v I__6014 (
            .O(N__26550),
            .I(N__26547));
    Sp12to4 I__6013 (
            .O(N__26547),
            .I(N__26544));
    Odrv12 I__6012 (
            .O(N__26544),
            .I(port_address_in_6));
    CascadeMux I__6011 (
            .O(N__26541),
            .I(N__26537));
    CascadeMux I__6010 (
            .O(N__26540),
            .I(N__26534));
    InMux I__6009 (
            .O(N__26537),
            .I(N__26529));
    InMux I__6008 (
            .O(N__26534),
            .I(N__26529));
    LocalMux I__6007 (
            .O(N__26529),
            .I(N__26526));
    Span4Mux_v I__6006 (
            .O(N__26526),
            .I(N__26523));
    Span4Mux_h I__6005 (
            .O(N__26523),
            .I(N__26520));
    Odrv4 I__6004 (
            .O(N__26520),
            .I(\this_vga_signals.M_this_state_q_srsts_0_0_a2_1_4_0 ));
    InMux I__6003 (
            .O(N__26517),
            .I(N__26514));
    LocalMux I__6002 (
            .O(N__26514),
            .I(N__26511));
    Span4Mux_h I__6001 (
            .O(N__26511),
            .I(N__26508));
    Odrv4 I__6000 (
            .O(N__26508),
            .I(N_54_0));
    InMux I__5999 (
            .O(N__26505),
            .I(N__26502));
    LocalMux I__5998 (
            .O(N__26502),
            .I(\this_ppu.un1_oam_data_1_c2 ));
    CascadeMux I__5997 (
            .O(N__26499),
            .I(N__26493));
    InMux I__5996 (
            .O(N__26498),
            .I(N__26484));
    InMux I__5995 (
            .O(N__26497),
            .I(N__26484));
    InMux I__5994 (
            .O(N__26496),
            .I(N__26484));
    InMux I__5993 (
            .O(N__26493),
            .I(N__26480));
    InMux I__5992 (
            .O(N__26492),
            .I(N__26475));
    InMux I__5991 (
            .O(N__26491),
            .I(N__26475));
    LocalMux I__5990 (
            .O(N__26484),
            .I(N__26472));
    InMux I__5989 (
            .O(N__26483),
            .I(N__26469));
    LocalMux I__5988 (
            .O(N__26480),
            .I(N__26466));
    LocalMux I__5987 (
            .O(N__26475),
            .I(N__26463));
    Span4Mux_h I__5986 (
            .O(N__26472),
            .I(N__26458));
    LocalMux I__5985 (
            .O(N__26469),
            .I(N__26458));
    Span4Mux_v I__5984 (
            .O(N__26466),
            .I(N__26455));
    Span4Mux_v I__5983 (
            .O(N__26463),
            .I(N__26450));
    Span4Mux_v I__5982 (
            .O(N__26458),
            .I(N__26450));
    Odrv4 I__5981 (
            .O(N__26455),
            .I(N_163));
    Odrv4 I__5980 (
            .O(N__26450),
            .I(N_163));
    InMux I__5979 (
            .O(N__26445),
            .I(N__26442));
    LocalMux I__5978 (
            .O(N__26442),
            .I(N__26438));
    InMux I__5977 (
            .O(N__26441),
            .I(N__26434));
    Span4Mux_v I__5976 (
            .O(N__26438),
            .I(N__26431));
    InMux I__5975 (
            .O(N__26437),
            .I(N__26428));
    LocalMux I__5974 (
            .O(N__26434),
            .I(un1_M_this_oam_address_q_c2));
    Odrv4 I__5973 (
            .O(N__26431),
            .I(un1_M_this_oam_address_q_c2));
    LocalMux I__5972 (
            .O(N__26428),
            .I(un1_M_this_oam_address_q_c2));
    CascadeMux I__5971 (
            .O(N__26421),
            .I(N__26418));
    CascadeBuf I__5970 (
            .O(N__26418),
            .I(N__26415));
    CascadeMux I__5969 (
            .O(N__26415),
            .I(N__26412));
    InMux I__5968 (
            .O(N__26412),
            .I(N__26408));
    InMux I__5967 (
            .O(N__26411),
            .I(N__26403));
    LocalMux I__5966 (
            .O(N__26408),
            .I(N__26400));
    InMux I__5965 (
            .O(N__26407),
            .I(N__26397));
    InMux I__5964 (
            .O(N__26406),
            .I(N__26394));
    LocalMux I__5963 (
            .O(N__26403),
            .I(N__26389));
    Span12Mux_s11_v I__5962 (
            .O(N__26400),
            .I(N__26389));
    LocalMux I__5961 (
            .O(N__26397),
            .I(M_this_oam_address_qZ0Z_2));
    LocalMux I__5960 (
            .O(N__26394),
            .I(M_this_oam_address_qZ0Z_2));
    Odrv12 I__5959 (
            .O(N__26389),
            .I(M_this_oam_address_qZ0Z_2));
    CEMux I__5958 (
            .O(N__26382),
            .I(N__26378));
    CEMux I__5957 (
            .O(N__26381),
            .I(N__26375));
    LocalMux I__5956 (
            .O(N__26378),
            .I(N__26371));
    LocalMux I__5955 (
            .O(N__26375),
            .I(N__26368));
    CEMux I__5954 (
            .O(N__26374),
            .I(N__26365));
    Span4Mux_v I__5953 (
            .O(N__26371),
            .I(N__26358));
    Span4Mux_v I__5952 (
            .O(N__26368),
            .I(N__26358));
    LocalMux I__5951 (
            .O(N__26365),
            .I(N__26358));
    Span4Mux_v I__5950 (
            .O(N__26358),
            .I(N__26355));
    Odrv4 I__5949 (
            .O(N__26355),
            .I(N_1190_0));
    CascadeMux I__5948 (
            .O(N__26352),
            .I(N__26349));
    InMux I__5947 (
            .O(N__26349),
            .I(N__26346));
    LocalMux I__5946 (
            .O(N__26346),
            .I(M_this_data_tmp_qZ0Z_6));
    InMux I__5945 (
            .O(N__26343),
            .I(N__26340));
    LocalMux I__5944 (
            .O(N__26340),
            .I(N__26337));
    Span4Mux_h I__5943 (
            .O(N__26337),
            .I(N__26334));
    Odrv4 I__5942 (
            .O(N__26334),
            .I(N_742_0));
    InMux I__5941 (
            .O(N__26331),
            .I(N__26328));
    LocalMux I__5940 (
            .O(N__26328),
            .I(N__26325));
    Span4Mux_v I__5939 (
            .O(N__26325),
            .I(N__26322));
    Span4Mux_h I__5938 (
            .O(N__26322),
            .I(N__26319));
    Odrv4 I__5937 (
            .O(N__26319),
            .I(N_34_0));
    InMux I__5936 (
            .O(N__26316),
            .I(N__26313));
    LocalMux I__5935 (
            .O(N__26313),
            .I(M_this_sprites_address_q_RNO_0Z0Z_2));
    InMux I__5934 (
            .O(N__26310),
            .I(N__26305));
    InMux I__5933 (
            .O(N__26309),
            .I(N__26302));
    InMux I__5932 (
            .O(N__26308),
            .I(N__26299));
    LocalMux I__5931 (
            .O(N__26305),
            .I(N__26293));
    LocalMux I__5930 (
            .O(N__26302),
            .I(N__26293));
    LocalMux I__5929 (
            .O(N__26299),
            .I(N__26290));
    InMux I__5928 (
            .O(N__26298),
            .I(N__26287));
    Span4Mux_h I__5927 (
            .O(N__26293),
            .I(N__26282));
    Span4Mux_v I__5926 (
            .O(N__26290),
            .I(N__26279));
    LocalMux I__5925 (
            .O(N__26287),
            .I(N__26276));
    InMux I__5924 (
            .O(N__26286),
            .I(N__26273));
    InMux I__5923 (
            .O(N__26285),
            .I(N__26270));
    Odrv4 I__5922 (
            .O(N__26282),
            .I(N_813));
    Odrv4 I__5921 (
            .O(N__26279),
            .I(N_813));
    Odrv12 I__5920 (
            .O(N__26276),
            .I(N_813));
    LocalMux I__5919 (
            .O(N__26273),
            .I(N_813));
    LocalMux I__5918 (
            .O(N__26270),
            .I(N_813));
    InMux I__5917 (
            .O(N__26259),
            .I(N__26256));
    LocalMux I__5916 (
            .O(N__26256),
            .I(N__26253));
    Span4Mux_v I__5915 (
            .O(N__26253),
            .I(N__26250));
    Odrv4 I__5914 (
            .O(N__26250),
            .I(N_799));
    CascadeMux I__5913 (
            .O(N__26247),
            .I(M_this_sprites_address_qc_11_0_cascade_));
    InMux I__5912 (
            .O(N__26244),
            .I(N__26241));
    LocalMux I__5911 (
            .O(N__26241),
            .I(M_this_sprites_address_q_RNO_1Z0Z_9));
    CascadeMux I__5910 (
            .O(N__26238),
            .I(N__26234));
    CascadeMux I__5909 (
            .O(N__26237),
            .I(N__26231));
    InMux I__5908 (
            .O(N__26234),
            .I(N__26224));
    InMux I__5907 (
            .O(N__26231),
            .I(N__26221));
    CascadeMux I__5906 (
            .O(N__26230),
            .I(N__26218));
    CascadeMux I__5905 (
            .O(N__26229),
            .I(N__26215));
    CascadeMux I__5904 (
            .O(N__26228),
            .I(N__26212));
    CascadeMux I__5903 (
            .O(N__26227),
            .I(N__26209));
    LocalMux I__5902 (
            .O(N__26224),
            .I(N__26204));
    LocalMux I__5901 (
            .O(N__26221),
            .I(N__26201));
    InMux I__5900 (
            .O(N__26218),
            .I(N__26198));
    InMux I__5899 (
            .O(N__26215),
            .I(N__26195));
    InMux I__5898 (
            .O(N__26212),
            .I(N__26192));
    InMux I__5897 (
            .O(N__26209),
            .I(N__26189));
    CascadeMux I__5896 (
            .O(N__26208),
            .I(N__26186));
    CascadeMux I__5895 (
            .O(N__26207),
            .I(N__26183));
    Span4Mux_v I__5894 (
            .O(N__26204),
            .I(N__26172));
    Span4Mux_h I__5893 (
            .O(N__26201),
            .I(N__26172));
    LocalMux I__5892 (
            .O(N__26198),
            .I(N__26172));
    LocalMux I__5891 (
            .O(N__26195),
            .I(N__26169));
    LocalMux I__5890 (
            .O(N__26192),
            .I(N__26166));
    LocalMux I__5889 (
            .O(N__26189),
            .I(N__26163));
    InMux I__5888 (
            .O(N__26186),
            .I(N__26160));
    InMux I__5887 (
            .O(N__26183),
            .I(N__26157));
    CascadeMux I__5886 (
            .O(N__26182),
            .I(N__26154));
    CascadeMux I__5885 (
            .O(N__26181),
            .I(N__26151));
    CascadeMux I__5884 (
            .O(N__26180),
            .I(N__26147));
    CascadeMux I__5883 (
            .O(N__26179),
            .I(N__26144));
    Span4Mux_v I__5882 (
            .O(N__26172),
            .I(N__26134));
    Span4Mux_v I__5881 (
            .O(N__26169),
            .I(N__26134));
    Span4Mux_h I__5880 (
            .O(N__26166),
            .I(N__26134));
    Span4Mux_s1_v I__5879 (
            .O(N__26163),
            .I(N__26129));
    LocalMux I__5878 (
            .O(N__26160),
            .I(N__26129));
    LocalMux I__5877 (
            .O(N__26157),
            .I(N__26126));
    InMux I__5876 (
            .O(N__26154),
            .I(N__26123));
    InMux I__5875 (
            .O(N__26151),
            .I(N__26120));
    CascadeMux I__5874 (
            .O(N__26150),
            .I(N__26117));
    InMux I__5873 (
            .O(N__26147),
            .I(N__26114));
    InMux I__5872 (
            .O(N__26144),
            .I(N__26111));
    CascadeMux I__5871 (
            .O(N__26143),
            .I(N__26108));
    CascadeMux I__5870 (
            .O(N__26142),
            .I(N__26105));
    CascadeMux I__5869 (
            .O(N__26141),
            .I(N__26102));
    Span4Mux_h I__5868 (
            .O(N__26134),
            .I(N__26099));
    Span4Mux_v I__5867 (
            .O(N__26129),
            .I(N__26092));
    Span4Mux_h I__5866 (
            .O(N__26126),
            .I(N__26092));
    LocalMux I__5865 (
            .O(N__26123),
            .I(N__26092));
    LocalMux I__5864 (
            .O(N__26120),
            .I(N__26089));
    InMux I__5863 (
            .O(N__26117),
            .I(N__26086));
    LocalMux I__5862 (
            .O(N__26114),
            .I(N__26081));
    LocalMux I__5861 (
            .O(N__26111),
            .I(N__26081));
    InMux I__5860 (
            .O(N__26108),
            .I(N__26078));
    InMux I__5859 (
            .O(N__26105),
            .I(N__26075));
    InMux I__5858 (
            .O(N__26102),
            .I(N__26072));
    Span4Mux_h I__5857 (
            .O(N__26099),
            .I(N__26069));
    Span4Mux_v I__5856 (
            .O(N__26092),
            .I(N__26062));
    Span4Mux_h I__5855 (
            .O(N__26089),
            .I(N__26062));
    LocalMux I__5854 (
            .O(N__26086),
            .I(N__26062));
    Span4Mux_v I__5853 (
            .O(N__26081),
            .I(N__26055));
    LocalMux I__5852 (
            .O(N__26078),
            .I(N__26055));
    LocalMux I__5851 (
            .O(N__26075),
            .I(N__26055));
    LocalMux I__5850 (
            .O(N__26072),
            .I(N__26052));
    Span4Mux_h I__5849 (
            .O(N__26069),
            .I(N__26041));
    Span4Mux_v I__5848 (
            .O(N__26062),
            .I(N__26041));
    Span4Mux_v I__5847 (
            .O(N__26055),
            .I(N__26041));
    Span4Mux_h I__5846 (
            .O(N__26052),
            .I(N__26041));
    InMux I__5845 (
            .O(N__26051),
            .I(N__26038));
    InMux I__5844 (
            .O(N__26050),
            .I(N__26035));
    Odrv4 I__5843 (
            .O(N__26041),
            .I(M_this_sprites_address_qZ0Z_9));
    LocalMux I__5842 (
            .O(N__26038),
            .I(M_this_sprites_address_qZ0Z_9));
    LocalMux I__5841 (
            .O(N__26035),
            .I(M_this_sprites_address_qZ0Z_9));
    InMux I__5840 (
            .O(N__26028),
            .I(N__26025));
    LocalMux I__5839 (
            .O(N__26025),
            .I(M_this_sprites_address_q_RNO_0Z0Z_3));
    CascadeMux I__5838 (
            .O(N__26022),
            .I(N__26015));
    CascadeMux I__5837 (
            .O(N__26021),
            .I(N__26012));
    CascadeMux I__5836 (
            .O(N__26020),
            .I(N__26009));
    CascadeMux I__5835 (
            .O(N__26019),
            .I(N__26001));
    CascadeMux I__5834 (
            .O(N__26018),
            .I(N__25997));
    InMux I__5833 (
            .O(N__26015),
            .I(N__25994));
    InMux I__5832 (
            .O(N__26012),
            .I(N__25991));
    InMux I__5831 (
            .O(N__26009),
            .I(N__25988));
    CascadeMux I__5830 (
            .O(N__26008),
            .I(N__25985));
    CascadeMux I__5829 (
            .O(N__26007),
            .I(N__25978));
    CascadeMux I__5828 (
            .O(N__26006),
            .I(N__25974));
    CascadeMux I__5827 (
            .O(N__26005),
            .I(N__25971));
    CascadeMux I__5826 (
            .O(N__26004),
            .I(N__25968));
    InMux I__5825 (
            .O(N__26001),
            .I(N__25965));
    CascadeMux I__5824 (
            .O(N__26000),
            .I(N__25962));
    InMux I__5823 (
            .O(N__25997),
            .I(N__25959));
    LocalMux I__5822 (
            .O(N__25994),
            .I(N__25956));
    LocalMux I__5821 (
            .O(N__25991),
            .I(N__25953));
    LocalMux I__5820 (
            .O(N__25988),
            .I(N__25950));
    InMux I__5819 (
            .O(N__25985),
            .I(N__25947));
    CascadeMux I__5818 (
            .O(N__25984),
            .I(N__25944));
    CascadeMux I__5817 (
            .O(N__25983),
            .I(N__25941));
    CascadeMux I__5816 (
            .O(N__25982),
            .I(N__25938));
    CascadeMux I__5815 (
            .O(N__25981),
            .I(N__25935));
    InMux I__5814 (
            .O(N__25978),
            .I(N__25932));
    CascadeMux I__5813 (
            .O(N__25977),
            .I(N__25929));
    InMux I__5812 (
            .O(N__25974),
            .I(N__25926));
    InMux I__5811 (
            .O(N__25971),
            .I(N__25923));
    InMux I__5810 (
            .O(N__25968),
            .I(N__25920));
    LocalMux I__5809 (
            .O(N__25965),
            .I(N__25917));
    InMux I__5808 (
            .O(N__25962),
            .I(N__25914));
    LocalMux I__5807 (
            .O(N__25959),
            .I(N__25911));
    Span4Mux_v I__5806 (
            .O(N__25956),
            .I(N__25902));
    Span4Mux_v I__5805 (
            .O(N__25953),
            .I(N__25902));
    Span4Mux_h I__5804 (
            .O(N__25950),
            .I(N__25902));
    LocalMux I__5803 (
            .O(N__25947),
            .I(N__25902));
    InMux I__5802 (
            .O(N__25944),
            .I(N__25899));
    InMux I__5801 (
            .O(N__25941),
            .I(N__25896));
    InMux I__5800 (
            .O(N__25938),
            .I(N__25893));
    InMux I__5799 (
            .O(N__25935),
            .I(N__25890));
    LocalMux I__5798 (
            .O(N__25932),
            .I(N__25887));
    InMux I__5797 (
            .O(N__25929),
            .I(N__25884));
    LocalMux I__5796 (
            .O(N__25926),
            .I(N__25881));
    LocalMux I__5795 (
            .O(N__25923),
            .I(N__25878));
    LocalMux I__5794 (
            .O(N__25920),
            .I(N__25875));
    Span4Mux_h I__5793 (
            .O(N__25917),
            .I(N__25871));
    LocalMux I__5792 (
            .O(N__25914),
            .I(N__25868));
    Span4Mux_h I__5791 (
            .O(N__25911),
            .I(N__25863));
    Span4Mux_v I__5790 (
            .O(N__25902),
            .I(N__25863));
    LocalMux I__5789 (
            .O(N__25899),
            .I(N__25858));
    LocalMux I__5788 (
            .O(N__25896),
            .I(N__25858));
    LocalMux I__5787 (
            .O(N__25893),
            .I(N__25851));
    LocalMux I__5786 (
            .O(N__25890),
            .I(N__25851));
    Span4Mux_v I__5785 (
            .O(N__25887),
            .I(N__25851));
    LocalMux I__5784 (
            .O(N__25884),
            .I(N__25848));
    Sp12to4 I__5783 (
            .O(N__25881),
            .I(N__25845));
    Span4Mux_h I__5782 (
            .O(N__25878),
            .I(N__25840));
    Span4Mux_h I__5781 (
            .O(N__25875),
            .I(N__25840));
    InMux I__5780 (
            .O(N__25874),
            .I(N__25837));
    Sp12to4 I__5779 (
            .O(N__25871),
            .I(N__25832));
    Span12Mux_s8_h I__5778 (
            .O(N__25868),
            .I(N__25832));
    Span4Mux_h I__5777 (
            .O(N__25863),
            .I(N__25829));
    Span4Mux_v I__5776 (
            .O(N__25858),
            .I(N__25823));
    Span4Mux_v I__5775 (
            .O(N__25851),
            .I(N__25823));
    Span12Mux_s10_h I__5774 (
            .O(N__25848),
            .I(N__25816));
    Span12Mux_s10_h I__5773 (
            .O(N__25845),
            .I(N__25816));
    Sp12to4 I__5772 (
            .O(N__25840),
            .I(N__25816));
    LocalMux I__5771 (
            .O(N__25837),
            .I(N__25813));
    Span12Mux_v I__5770 (
            .O(N__25832),
            .I(N__25808));
    Sp12to4 I__5769 (
            .O(N__25829),
            .I(N__25808));
    InMux I__5768 (
            .O(N__25828),
            .I(N__25805));
    Odrv4 I__5767 (
            .O(N__25823),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv12 I__5766 (
            .O(N__25816),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv4 I__5765 (
            .O(N__25813),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv12 I__5764 (
            .O(N__25808),
            .I(M_this_sprites_address_qZ0Z_3));
    LocalMux I__5763 (
            .O(N__25805),
            .I(M_this_sprites_address_qZ0Z_3));
    CascadeMux I__5762 (
            .O(N__25794),
            .I(N__25791));
    InMux I__5761 (
            .O(N__25791),
            .I(N__25788));
    LocalMux I__5760 (
            .O(N__25788),
            .I(N_50));
    CascadeMux I__5759 (
            .O(N__25785),
            .I(N__25780));
    CascadeMux I__5758 (
            .O(N__25784),
            .I(N__25777));
    CascadeMux I__5757 (
            .O(N__25783),
            .I(N__25773));
    InMux I__5756 (
            .O(N__25780),
            .I(N__25768));
    InMux I__5755 (
            .O(N__25777),
            .I(N__25765));
    CascadeMux I__5754 (
            .O(N__25776),
            .I(N__25762));
    InMux I__5753 (
            .O(N__25773),
            .I(N__25758));
    CascadeMux I__5752 (
            .O(N__25772),
            .I(N__25755));
    CascadeMux I__5751 (
            .O(N__25771),
            .I(N__25752));
    LocalMux I__5750 (
            .O(N__25768),
            .I(N__25746));
    LocalMux I__5749 (
            .O(N__25765),
            .I(N__25746));
    InMux I__5748 (
            .O(N__25762),
            .I(N__25743));
    CascadeMux I__5747 (
            .O(N__25761),
            .I(N__25740));
    LocalMux I__5746 (
            .O(N__25758),
            .I(N__25736));
    InMux I__5745 (
            .O(N__25755),
            .I(N__25733));
    InMux I__5744 (
            .O(N__25752),
            .I(N__25730));
    CascadeMux I__5743 (
            .O(N__25751),
            .I(N__25727));
    Span4Mux_s2_v I__5742 (
            .O(N__25746),
            .I(N__25720));
    LocalMux I__5741 (
            .O(N__25743),
            .I(N__25720));
    InMux I__5740 (
            .O(N__25740),
            .I(N__25717));
    CascadeMux I__5739 (
            .O(N__25739),
            .I(N__25714));
    Span4Mux_h I__5738 (
            .O(N__25736),
            .I(N__25708));
    LocalMux I__5737 (
            .O(N__25733),
            .I(N__25708));
    LocalMux I__5736 (
            .O(N__25730),
            .I(N__25705));
    InMux I__5735 (
            .O(N__25727),
            .I(N__25702));
    CascadeMux I__5734 (
            .O(N__25726),
            .I(N__25698));
    CascadeMux I__5733 (
            .O(N__25725),
            .I(N__25695));
    Span4Mux_v I__5732 (
            .O(N__25720),
            .I(N__25689));
    LocalMux I__5731 (
            .O(N__25717),
            .I(N__25689));
    InMux I__5730 (
            .O(N__25714),
            .I(N__25686));
    CascadeMux I__5729 (
            .O(N__25713),
            .I(N__25683));
    Span4Mux_v I__5728 (
            .O(N__25708),
            .I(N__25675));
    Span4Mux_h I__5727 (
            .O(N__25705),
            .I(N__25675));
    LocalMux I__5726 (
            .O(N__25702),
            .I(N__25675));
    CascadeMux I__5725 (
            .O(N__25701),
            .I(N__25672));
    InMux I__5724 (
            .O(N__25698),
            .I(N__25669));
    InMux I__5723 (
            .O(N__25695),
            .I(N__25666));
    CascadeMux I__5722 (
            .O(N__25694),
            .I(N__25663));
    Span4Mux_h I__5721 (
            .O(N__25689),
            .I(N__25658));
    LocalMux I__5720 (
            .O(N__25686),
            .I(N__25658));
    InMux I__5719 (
            .O(N__25683),
            .I(N__25655));
    CascadeMux I__5718 (
            .O(N__25682),
            .I(N__25652));
    Span4Mux_v I__5717 (
            .O(N__25675),
            .I(N__25648));
    InMux I__5716 (
            .O(N__25672),
            .I(N__25645));
    LocalMux I__5715 (
            .O(N__25669),
            .I(N__25642));
    LocalMux I__5714 (
            .O(N__25666),
            .I(N__25639));
    InMux I__5713 (
            .O(N__25663),
            .I(N__25636));
    Span4Mux_v I__5712 (
            .O(N__25658),
            .I(N__25631));
    LocalMux I__5711 (
            .O(N__25655),
            .I(N__25631));
    InMux I__5710 (
            .O(N__25652),
            .I(N__25628));
    CascadeMux I__5709 (
            .O(N__25651),
            .I(N__25625));
    Sp12to4 I__5708 (
            .O(N__25648),
            .I(N__25620));
    LocalMux I__5707 (
            .O(N__25645),
            .I(N__25620));
    Span4Mux_v I__5706 (
            .O(N__25642),
            .I(N__25613));
    Span4Mux_h I__5705 (
            .O(N__25639),
            .I(N__25613));
    LocalMux I__5704 (
            .O(N__25636),
            .I(N__25613));
    Span4Mux_h I__5703 (
            .O(N__25631),
            .I(N__25608));
    LocalMux I__5702 (
            .O(N__25628),
            .I(N__25608));
    InMux I__5701 (
            .O(N__25625),
            .I(N__25605));
    Span12Mux_h I__5700 (
            .O(N__25620),
            .I(N__25602));
    Span4Mux_v I__5699 (
            .O(N__25613),
            .I(N__25595));
    Span4Mux_v I__5698 (
            .O(N__25608),
            .I(N__25595));
    LocalMux I__5697 (
            .O(N__25605),
            .I(N__25595));
    Odrv12 I__5696 (
            .O(N__25602),
            .I(M_this_ppu_sprites_addr_3));
    Odrv4 I__5695 (
            .O(N__25595),
            .I(M_this_ppu_sprites_addr_3));
    CascadeMux I__5694 (
            .O(N__25590),
            .I(N__25585));
    CascadeMux I__5693 (
            .O(N__25589),
            .I(N__25581));
    CascadeMux I__5692 (
            .O(N__25588),
            .I(N__25578));
    InMux I__5691 (
            .O(N__25585),
            .I(N__25573));
    CascadeMux I__5690 (
            .O(N__25584),
            .I(N__25570));
    InMux I__5689 (
            .O(N__25581),
            .I(N__25566));
    InMux I__5688 (
            .O(N__25578),
            .I(N__25563));
    CascadeMux I__5687 (
            .O(N__25577),
            .I(N__25560));
    CascadeMux I__5686 (
            .O(N__25576),
            .I(N__25557));
    LocalMux I__5685 (
            .O(N__25573),
            .I(N__25554));
    InMux I__5684 (
            .O(N__25570),
            .I(N__25551));
    CascadeMux I__5683 (
            .O(N__25569),
            .I(N__25548));
    LocalMux I__5682 (
            .O(N__25566),
            .I(N__25541));
    LocalMux I__5681 (
            .O(N__25563),
            .I(N__25538));
    InMux I__5680 (
            .O(N__25560),
            .I(N__25535));
    InMux I__5679 (
            .O(N__25557),
            .I(N__25532));
    Span4Mux_v I__5678 (
            .O(N__25554),
            .I(N__25526));
    LocalMux I__5677 (
            .O(N__25551),
            .I(N__25526));
    InMux I__5676 (
            .O(N__25548),
            .I(N__25523));
    CascadeMux I__5675 (
            .O(N__25547),
            .I(N__25520));
    CascadeMux I__5674 (
            .O(N__25546),
            .I(N__25516));
    CascadeMux I__5673 (
            .O(N__25545),
            .I(N__25513));
    CascadeMux I__5672 (
            .O(N__25544),
            .I(N__25508));
    Span4Mux_v I__5671 (
            .O(N__25541),
            .I(N__25501));
    Span4Mux_h I__5670 (
            .O(N__25538),
            .I(N__25501));
    LocalMux I__5669 (
            .O(N__25535),
            .I(N__25501));
    LocalMux I__5668 (
            .O(N__25532),
            .I(N__25498));
    CascadeMux I__5667 (
            .O(N__25531),
            .I(N__25495));
    Span4Mux_h I__5666 (
            .O(N__25526),
            .I(N__25490));
    LocalMux I__5665 (
            .O(N__25523),
            .I(N__25490));
    InMux I__5664 (
            .O(N__25520),
            .I(N__25487));
    CascadeMux I__5663 (
            .O(N__25519),
            .I(N__25484));
    InMux I__5662 (
            .O(N__25516),
            .I(N__25481));
    InMux I__5661 (
            .O(N__25513),
            .I(N__25478));
    CascadeMux I__5660 (
            .O(N__25512),
            .I(N__25475));
    CascadeMux I__5659 (
            .O(N__25511),
            .I(N__25472));
    InMux I__5658 (
            .O(N__25508),
            .I(N__25468));
    Span4Mux_v I__5657 (
            .O(N__25501),
            .I(N__25463));
    Span4Mux_v I__5656 (
            .O(N__25498),
            .I(N__25463));
    InMux I__5655 (
            .O(N__25495),
            .I(N__25460));
    Span4Mux_v I__5654 (
            .O(N__25490),
            .I(N__25455));
    LocalMux I__5653 (
            .O(N__25487),
            .I(N__25455));
    InMux I__5652 (
            .O(N__25484),
            .I(N__25452));
    LocalMux I__5651 (
            .O(N__25481),
            .I(N__25449));
    LocalMux I__5650 (
            .O(N__25478),
            .I(N__25446));
    InMux I__5649 (
            .O(N__25475),
            .I(N__25443));
    InMux I__5648 (
            .O(N__25472),
            .I(N__25440));
    CascadeMux I__5647 (
            .O(N__25471),
            .I(N__25437));
    LocalMux I__5646 (
            .O(N__25468),
            .I(N__25434));
    Sp12to4 I__5645 (
            .O(N__25463),
            .I(N__25429));
    LocalMux I__5644 (
            .O(N__25460),
            .I(N__25429));
    Span4Mux_h I__5643 (
            .O(N__25455),
            .I(N__25424));
    LocalMux I__5642 (
            .O(N__25452),
            .I(N__25424));
    Span4Mux_v I__5641 (
            .O(N__25449),
            .I(N__25415));
    Span4Mux_v I__5640 (
            .O(N__25446),
            .I(N__25415));
    LocalMux I__5639 (
            .O(N__25443),
            .I(N__25415));
    LocalMux I__5638 (
            .O(N__25440),
            .I(N__25415));
    InMux I__5637 (
            .O(N__25437),
            .I(N__25412));
    Span12Mux_s10_h I__5636 (
            .O(N__25434),
            .I(N__25407));
    Span12Mux_h I__5635 (
            .O(N__25429),
            .I(N__25404));
    Span4Mux_v I__5634 (
            .O(N__25424),
            .I(N__25397));
    Span4Mux_v I__5633 (
            .O(N__25415),
            .I(N__25397));
    LocalMux I__5632 (
            .O(N__25412),
            .I(N__25397));
    InMux I__5631 (
            .O(N__25411),
            .I(N__25394));
    InMux I__5630 (
            .O(N__25410),
            .I(N__25391));
    Odrv12 I__5629 (
            .O(N__25407),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv12 I__5628 (
            .O(N__25404),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv4 I__5627 (
            .O(N__25397),
            .I(M_this_sprites_address_qZ0Z_2));
    LocalMux I__5626 (
            .O(N__25394),
            .I(M_this_sprites_address_qZ0Z_2));
    LocalMux I__5625 (
            .O(N__25391),
            .I(M_this_sprites_address_qZ0Z_2));
    CascadeMux I__5624 (
            .O(N__25380),
            .I(N__25377));
    InMux I__5623 (
            .O(N__25377),
            .I(N__25374));
    LocalMux I__5622 (
            .O(N__25374),
            .I(N_103));
    InMux I__5621 (
            .O(N__25371),
            .I(N__25367));
    InMux I__5620 (
            .O(N__25370),
            .I(N__25363));
    LocalMux I__5619 (
            .O(N__25367),
            .I(N__25359));
    InMux I__5618 (
            .O(N__25366),
            .I(N__25356));
    LocalMux I__5617 (
            .O(N__25363),
            .I(N__25353));
    InMux I__5616 (
            .O(N__25362),
            .I(N__25350));
    Span4Mux_v I__5615 (
            .O(N__25359),
            .I(N__25343));
    LocalMux I__5614 (
            .O(N__25356),
            .I(N__25343));
    Span4Mux_s3_v I__5613 (
            .O(N__25353),
            .I(N__25337));
    LocalMux I__5612 (
            .O(N__25350),
            .I(N__25337));
    InMux I__5611 (
            .O(N__25349),
            .I(N__25334));
    InMux I__5610 (
            .O(N__25348),
            .I(N__25331));
    Span4Mux_v I__5609 (
            .O(N__25343),
            .I(N__25327));
    InMux I__5608 (
            .O(N__25342),
            .I(N__25324));
    Span4Mux_v I__5607 (
            .O(N__25337),
            .I(N__25317));
    LocalMux I__5606 (
            .O(N__25334),
            .I(N__25317));
    LocalMux I__5605 (
            .O(N__25331),
            .I(N__25317));
    InMux I__5604 (
            .O(N__25330),
            .I(N__25314));
    Sp12to4 I__5603 (
            .O(N__25327),
            .I(N__25311));
    LocalMux I__5602 (
            .O(N__25324),
            .I(N__25308));
    Span4Mux_v I__5601 (
            .O(N__25317),
            .I(N__25303));
    LocalMux I__5600 (
            .O(N__25314),
            .I(N__25303));
    Span12Mux_h I__5599 (
            .O(N__25311),
            .I(N__25300));
    Span4Mux_v I__5598 (
            .O(N__25308),
            .I(N__25295));
    Span4Mux_v I__5597 (
            .O(N__25303),
            .I(N__25295));
    Odrv12 I__5596 (
            .O(N__25300),
            .I(M_this_sprites_ram_write_data_iv_i_i_1));
    Odrv4 I__5595 (
            .O(N__25295),
            .I(M_this_sprites_ram_write_data_iv_i_i_1));
    CascadeMux I__5594 (
            .O(N__25290),
            .I(N__25287));
    InMux I__5593 (
            .O(N__25287),
            .I(N__25284));
    LocalMux I__5592 (
            .O(N__25284),
            .I(N__25281));
    Odrv4 I__5591 (
            .O(N__25281),
            .I(M_this_data_tmp_qZ0Z_2));
    InMux I__5590 (
            .O(N__25278),
            .I(N__25275));
    LocalMux I__5589 (
            .O(N__25275),
            .I(N__25272));
    Span4Mux_v I__5588 (
            .O(N__25272),
            .I(N__25269));
    Span4Mux_h I__5587 (
            .O(N__25269),
            .I(N__25266));
    Odrv4 I__5586 (
            .O(N__25266),
            .I(N_746_0));
    InMux I__5585 (
            .O(N__25263),
            .I(N__25260));
    LocalMux I__5584 (
            .O(N__25260),
            .I(N__25257));
    Span4Mux_h I__5583 (
            .O(N__25257),
            .I(N__25254));
    Odrv4 I__5582 (
            .O(N__25254),
            .I(M_this_oam_ram_write_data_28));
    InMux I__5581 (
            .O(N__25251),
            .I(N__25248));
    LocalMux I__5580 (
            .O(N__25248),
            .I(N__25241));
    InMux I__5579 (
            .O(N__25247),
            .I(N__25238));
    InMux I__5578 (
            .O(N__25246),
            .I(N__25235));
    InMux I__5577 (
            .O(N__25245),
            .I(N__25229));
    InMux I__5576 (
            .O(N__25244),
            .I(N__25226));
    Span4Mux_h I__5575 (
            .O(N__25241),
            .I(N__25222));
    LocalMux I__5574 (
            .O(N__25238),
            .I(N__25217));
    LocalMux I__5573 (
            .O(N__25235),
            .I(N__25217));
    InMux I__5572 (
            .O(N__25234),
            .I(N__25210));
    InMux I__5571 (
            .O(N__25233),
            .I(N__25210));
    InMux I__5570 (
            .O(N__25232),
            .I(N__25210));
    LocalMux I__5569 (
            .O(N__25229),
            .I(N__25205));
    LocalMux I__5568 (
            .O(N__25226),
            .I(N__25205));
    InMux I__5567 (
            .O(N__25225),
            .I(N__25202));
    Span4Mux_h I__5566 (
            .O(N__25222),
            .I(N__25199));
    Span4Mux_v I__5565 (
            .O(N__25217),
            .I(N__25194));
    LocalMux I__5564 (
            .O(N__25210),
            .I(N__25194));
    Span4Mux_h I__5563 (
            .O(N__25205),
            .I(N__25191));
    LocalMux I__5562 (
            .O(N__25202),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__5561 (
            .O(N__25199),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__5560 (
            .O(N__25194),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__5559 (
            .O(N__25191),
            .I(M_this_state_qZ0Z_4));
    InMux I__5558 (
            .O(N__25182),
            .I(N__25179));
    LocalMux I__5557 (
            .O(N__25179),
            .I(un1_M_this_sprites_address_q_cry_0_THRU_CO));
    CascadeMux I__5556 (
            .O(N__25176),
            .I(N__25173));
    InMux I__5555 (
            .O(N__25173),
            .I(N__25165));
    CascadeMux I__5554 (
            .O(N__25172),
            .I(N__25162));
    CascadeMux I__5553 (
            .O(N__25171),
            .I(N__25159));
    CascadeMux I__5552 (
            .O(N__25170),
            .I(N__25152));
    CascadeMux I__5551 (
            .O(N__25169),
            .I(N__25149));
    CascadeMux I__5550 (
            .O(N__25168),
            .I(N__25146));
    LocalMux I__5549 (
            .O(N__25165),
            .I(N__25143));
    InMux I__5548 (
            .O(N__25162),
            .I(N__25140));
    InMux I__5547 (
            .O(N__25159),
            .I(N__25137));
    CascadeMux I__5546 (
            .O(N__25158),
            .I(N__25134));
    CascadeMux I__5545 (
            .O(N__25157),
            .I(N__25131));
    CascadeMux I__5544 (
            .O(N__25156),
            .I(N__25124));
    CascadeMux I__5543 (
            .O(N__25155),
            .I(N__25121));
    InMux I__5542 (
            .O(N__25152),
            .I(N__25118));
    InMux I__5541 (
            .O(N__25149),
            .I(N__25115));
    InMux I__5540 (
            .O(N__25146),
            .I(N__25110));
    Span4Mux_h I__5539 (
            .O(N__25143),
            .I(N__25103));
    LocalMux I__5538 (
            .O(N__25140),
            .I(N__25103));
    LocalMux I__5537 (
            .O(N__25137),
            .I(N__25103));
    InMux I__5536 (
            .O(N__25134),
            .I(N__25100));
    InMux I__5535 (
            .O(N__25131),
            .I(N__25097));
    CascadeMux I__5534 (
            .O(N__25130),
            .I(N__25094));
    CascadeMux I__5533 (
            .O(N__25129),
            .I(N__25091));
    CascadeMux I__5532 (
            .O(N__25128),
            .I(N__25088));
    CascadeMux I__5531 (
            .O(N__25127),
            .I(N__25085));
    InMux I__5530 (
            .O(N__25124),
            .I(N__25082));
    InMux I__5529 (
            .O(N__25121),
            .I(N__25079));
    LocalMux I__5528 (
            .O(N__25118),
            .I(N__25076));
    LocalMux I__5527 (
            .O(N__25115),
            .I(N__25073));
    CascadeMux I__5526 (
            .O(N__25114),
            .I(N__25070));
    CascadeMux I__5525 (
            .O(N__25113),
            .I(N__25067));
    LocalMux I__5524 (
            .O(N__25110),
            .I(N__25064));
    Span4Mux_v I__5523 (
            .O(N__25103),
            .I(N__25059));
    LocalMux I__5522 (
            .O(N__25100),
            .I(N__25059));
    LocalMux I__5521 (
            .O(N__25097),
            .I(N__25056));
    InMux I__5520 (
            .O(N__25094),
            .I(N__25053));
    InMux I__5519 (
            .O(N__25091),
            .I(N__25050));
    InMux I__5518 (
            .O(N__25088),
            .I(N__25047));
    InMux I__5517 (
            .O(N__25085),
            .I(N__25044));
    LocalMux I__5516 (
            .O(N__25082),
            .I(N__25041));
    LocalMux I__5515 (
            .O(N__25079),
            .I(N__25038));
    Span4Mux_h I__5514 (
            .O(N__25076),
            .I(N__25033));
    Span4Mux_h I__5513 (
            .O(N__25073),
            .I(N__25033));
    InMux I__5512 (
            .O(N__25070),
            .I(N__25030));
    InMux I__5511 (
            .O(N__25067),
            .I(N__25027));
    Span4Mux_h I__5510 (
            .O(N__25064),
            .I(N__25022));
    Span4Mux_v I__5509 (
            .O(N__25059),
            .I(N__25022));
    Span4Mux_v I__5508 (
            .O(N__25056),
            .I(N__25019));
    LocalMux I__5507 (
            .O(N__25053),
            .I(N__25013));
    LocalMux I__5506 (
            .O(N__25050),
            .I(N__25013));
    LocalMux I__5505 (
            .O(N__25047),
            .I(N__25008));
    LocalMux I__5504 (
            .O(N__25044),
            .I(N__25008));
    Span4Mux_h I__5503 (
            .O(N__25041),
            .I(N__25005));
    Span4Mux_h I__5502 (
            .O(N__25038),
            .I(N__25002));
    Sp12to4 I__5501 (
            .O(N__25033),
            .I(N__24998));
    LocalMux I__5500 (
            .O(N__25030),
            .I(N__24995));
    LocalMux I__5499 (
            .O(N__25027),
            .I(N__24992));
    Sp12to4 I__5498 (
            .O(N__25022),
            .I(N__24989));
    Span4Mux_h I__5497 (
            .O(N__25019),
            .I(N__24986));
    InMux I__5496 (
            .O(N__25018),
            .I(N__24983));
    Span4Mux_v I__5495 (
            .O(N__25013),
            .I(N__24978));
    Span4Mux_v I__5494 (
            .O(N__25008),
            .I(N__24978));
    Span4Mux_v I__5493 (
            .O(N__25005),
            .I(N__24973));
    Span4Mux_v I__5492 (
            .O(N__25002),
            .I(N__24973));
    InMux I__5491 (
            .O(N__25001),
            .I(N__24970));
    Span12Mux_v I__5490 (
            .O(N__24998),
            .I(N__24967));
    Span12Mux_s11_h I__5489 (
            .O(N__24995),
            .I(N__24960));
    Span12Mux_s11_h I__5488 (
            .O(N__24992),
            .I(N__24960));
    Span12Mux_h I__5487 (
            .O(N__24989),
            .I(N__24960));
    Span4Mux_v I__5486 (
            .O(N__24986),
            .I(N__24955));
    LocalMux I__5485 (
            .O(N__24983),
            .I(N__24955));
    Odrv4 I__5484 (
            .O(N__24978),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv4 I__5483 (
            .O(N__24973),
            .I(M_this_sprites_address_qZ0Z_7));
    LocalMux I__5482 (
            .O(N__24970),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv12 I__5481 (
            .O(N__24967),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv12 I__5480 (
            .O(N__24960),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv4 I__5479 (
            .O(N__24955),
            .I(M_this_sprites_address_qZ0Z_7));
    InMux I__5478 (
            .O(N__24942),
            .I(N__24939));
    LocalMux I__5477 (
            .O(N__24939),
            .I(M_this_sprites_address_qc_9_0));
    CascadeMux I__5476 (
            .O(N__24936),
            .I(N__24933));
    InMux I__5475 (
            .O(N__24933),
            .I(N__24930));
    LocalMux I__5474 (
            .O(N__24930),
            .I(N__24927));
    Odrv12 I__5473 (
            .O(N__24927),
            .I(M_this_oam_ram_read_data_i_19));
    CascadeMux I__5472 (
            .O(N__24924),
            .I(N__24921));
    InMux I__5471 (
            .O(N__24921),
            .I(N__24918));
    LocalMux I__5470 (
            .O(N__24918),
            .I(N__24915));
    Odrv4 I__5469 (
            .O(N__24915),
            .I(M_this_oam_ram_read_data_i_11));
    CascadeMux I__5468 (
            .O(N__24912),
            .I(N__24909));
    InMux I__5467 (
            .O(N__24909),
            .I(N__24905));
    CascadeMux I__5466 (
            .O(N__24908),
            .I(N__24902));
    LocalMux I__5465 (
            .O(N__24905),
            .I(N__24899));
    InMux I__5464 (
            .O(N__24902),
            .I(N__24896));
    Span4Mux_h I__5463 (
            .O(N__24899),
            .I(N__24891));
    LocalMux I__5462 (
            .O(N__24896),
            .I(N__24891));
    Span4Mux_h I__5461 (
            .O(N__24891),
            .I(N__24888));
    Odrv4 I__5460 (
            .O(N__24888),
            .I(M_this_oam_ram_read_data_15));
    InMux I__5459 (
            .O(N__24885),
            .I(N__24882));
    LocalMux I__5458 (
            .O(N__24882),
            .I(N__24879));
    Odrv4 I__5457 (
            .O(N__24879),
            .I(\this_ppu.un1_M_haddress_q_2_7 ));
    CascadeMux I__5456 (
            .O(N__24876),
            .I(N__24873));
    CascadeBuf I__5455 (
            .O(N__24873),
            .I(N__24870));
    CascadeMux I__5454 (
            .O(N__24870),
            .I(N__24867));
    InMux I__5453 (
            .O(N__24867),
            .I(N__24864));
    LocalMux I__5452 (
            .O(N__24864),
            .I(N__24861));
    Span4Mux_h I__5451 (
            .O(N__24861),
            .I(N__24857));
    InMux I__5450 (
            .O(N__24860),
            .I(N__24854));
    Span4Mux_h I__5449 (
            .O(N__24857),
            .I(N__24850));
    LocalMux I__5448 (
            .O(N__24854),
            .I(N__24847));
    InMux I__5447 (
            .O(N__24853),
            .I(N__24844));
    Span4Mux_v I__5446 (
            .O(N__24850),
            .I(N__24841));
    Odrv12 I__5445 (
            .O(N__24847),
            .I(M_this_oam_address_qZ0Z_4));
    LocalMux I__5444 (
            .O(N__24844),
            .I(M_this_oam_address_qZ0Z_4));
    Odrv4 I__5443 (
            .O(N__24841),
            .I(M_this_oam_address_qZ0Z_4));
    InMux I__5442 (
            .O(N__24834),
            .I(N__24830));
    InMux I__5441 (
            .O(N__24833),
            .I(N__24827));
    LocalMux I__5440 (
            .O(N__24830),
            .I(un1_M_this_oam_address_q_c4));
    LocalMux I__5439 (
            .O(N__24827),
            .I(un1_M_this_oam_address_q_c4));
    CascadeMux I__5438 (
            .O(N__24822),
            .I(N__24819));
    CascadeBuf I__5437 (
            .O(N__24819),
            .I(N__24816));
    CascadeMux I__5436 (
            .O(N__24816),
            .I(N__24813));
    InMux I__5435 (
            .O(N__24813),
            .I(N__24810));
    LocalMux I__5434 (
            .O(N__24810),
            .I(N__24806));
    CascadeMux I__5433 (
            .O(N__24809),
            .I(N__24803));
    Span4Mux_v I__5432 (
            .O(N__24806),
            .I(N__24800));
    InMux I__5431 (
            .O(N__24803),
            .I(N__24797));
    Span4Mux_h I__5430 (
            .O(N__24800),
            .I(N__24794));
    LocalMux I__5429 (
            .O(N__24797),
            .I(M_this_oam_address_qZ0Z_5));
    Odrv4 I__5428 (
            .O(N__24794),
            .I(M_this_oam_address_qZ0Z_5));
    CascadeMux I__5427 (
            .O(N__24789),
            .I(N__24786));
    CascadeBuf I__5426 (
            .O(N__24786),
            .I(N__24783));
    CascadeMux I__5425 (
            .O(N__24783),
            .I(N__24780));
    InMux I__5424 (
            .O(N__24780),
            .I(N__24776));
    CascadeMux I__5423 (
            .O(N__24779),
            .I(N__24773));
    LocalMux I__5422 (
            .O(N__24776),
            .I(N__24769));
    InMux I__5421 (
            .O(N__24773),
            .I(N__24766));
    InMux I__5420 (
            .O(N__24772),
            .I(N__24763));
    Span12Mux_s11_v I__5419 (
            .O(N__24769),
            .I(N__24760));
    LocalMux I__5418 (
            .O(N__24766),
            .I(M_this_oam_address_qZ0Z_3));
    LocalMux I__5417 (
            .O(N__24763),
            .I(M_this_oam_address_qZ0Z_3));
    Odrv12 I__5416 (
            .O(N__24760),
            .I(M_this_oam_address_qZ0Z_3));
    InMux I__5415 (
            .O(N__24753),
            .I(N__24750));
    LocalMux I__5414 (
            .O(N__24750),
            .I(M_this_sprites_address_qc_2_1));
    InMux I__5413 (
            .O(N__24747),
            .I(un1_M_this_sprites_address_q_cry_12));
    InMux I__5412 (
            .O(N__24744),
            .I(N__24741));
    LocalMux I__5411 (
            .O(N__24741),
            .I(M_this_sprites_address_q_RNO_0Z0Z_12));
    CascadeMux I__5410 (
            .O(N__24738),
            .I(N_807_cascade_));
    InMux I__5409 (
            .O(N__24735),
            .I(N__24732));
    LocalMux I__5408 (
            .O(N__24732),
            .I(N__24729));
    Odrv4 I__5407 (
            .O(N__24729),
            .I(M_this_sprites_address_q_RNO_1Z0Z_7));
    InMux I__5406 (
            .O(N__24726),
            .I(N__24723));
    LocalMux I__5405 (
            .O(N__24723),
            .I(M_this_sprites_address_q_RNO_1Z0Z_8));
    CascadeMux I__5404 (
            .O(N__24720),
            .I(N_803_cascade_));
    InMux I__5403 (
            .O(N__24717),
            .I(N__24714));
    LocalMux I__5402 (
            .O(N__24714),
            .I(M_this_sprites_address_qc_10_0));
    CascadeMux I__5401 (
            .O(N__24711),
            .I(N__24708));
    InMux I__5400 (
            .O(N__24708),
            .I(N__24702));
    CascadeMux I__5399 (
            .O(N__24707),
            .I(N__24699));
    CascadeMux I__5398 (
            .O(N__24706),
            .I(N__24695));
    CascadeMux I__5397 (
            .O(N__24705),
            .I(N__24692));
    LocalMux I__5396 (
            .O(N__24702),
            .I(N__24686));
    InMux I__5395 (
            .O(N__24699),
            .I(N__24683));
    CascadeMux I__5394 (
            .O(N__24698),
            .I(N__24680));
    InMux I__5393 (
            .O(N__24695),
            .I(N__24674));
    InMux I__5392 (
            .O(N__24692),
            .I(N__24671));
    CascadeMux I__5391 (
            .O(N__24691),
            .I(N__24668));
    CascadeMux I__5390 (
            .O(N__24690),
            .I(N__24665));
    CascadeMux I__5389 (
            .O(N__24689),
            .I(N__24662));
    Span4Mux_s3_v I__5388 (
            .O(N__24686),
            .I(N__24657));
    LocalMux I__5387 (
            .O(N__24683),
            .I(N__24657));
    InMux I__5386 (
            .O(N__24680),
            .I(N__24654));
    CascadeMux I__5385 (
            .O(N__24679),
            .I(N__24651));
    CascadeMux I__5384 (
            .O(N__24678),
            .I(N__24647));
    CascadeMux I__5383 (
            .O(N__24677),
            .I(N__24644));
    LocalMux I__5382 (
            .O(N__24674),
            .I(N__24637));
    LocalMux I__5381 (
            .O(N__24671),
            .I(N__24637));
    InMux I__5380 (
            .O(N__24668),
            .I(N__24634));
    InMux I__5379 (
            .O(N__24665),
            .I(N__24631));
    InMux I__5378 (
            .O(N__24662),
            .I(N__24628));
    Span4Mux_h I__5377 (
            .O(N__24657),
            .I(N__24623));
    LocalMux I__5376 (
            .O(N__24654),
            .I(N__24623));
    InMux I__5375 (
            .O(N__24651),
            .I(N__24620));
    CascadeMux I__5374 (
            .O(N__24650),
            .I(N__24617));
    InMux I__5373 (
            .O(N__24647),
            .I(N__24613));
    InMux I__5372 (
            .O(N__24644),
            .I(N__24610));
    CascadeMux I__5371 (
            .O(N__24643),
            .I(N__24607));
    CascadeMux I__5370 (
            .O(N__24642),
            .I(N__24604));
    Span4Mux_v I__5369 (
            .O(N__24637),
            .I(N__24596));
    LocalMux I__5368 (
            .O(N__24634),
            .I(N__24596));
    LocalMux I__5367 (
            .O(N__24631),
            .I(N__24596));
    LocalMux I__5366 (
            .O(N__24628),
            .I(N__24593));
    Span4Mux_v I__5365 (
            .O(N__24623),
            .I(N__24588));
    LocalMux I__5364 (
            .O(N__24620),
            .I(N__24588));
    InMux I__5363 (
            .O(N__24617),
            .I(N__24585));
    CascadeMux I__5362 (
            .O(N__24616),
            .I(N__24582));
    LocalMux I__5361 (
            .O(N__24613),
            .I(N__24579));
    LocalMux I__5360 (
            .O(N__24610),
            .I(N__24576));
    InMux I__5359 (
            .O(N__24607),
            .I(N__24573));
    InMux I__5358 (
            .O(N__24604),
            .I(N__24570));
    CascadeMux I__5357 (
            .O(N__24603),
            .I(N__24567));
    Span4Mux_v I__5356 (
            .O(N__24596),
            .I(N__24562));
    Span4Mux_v I__5355 (
            .O(N__24593),
            .I(N__24562));
    Span4Mux_h I__5354 (
            .O(N__24588),
            .I(N__24557));
    LocalMux I__5353 (
            .O(N__24585),
            .I(N__24557));
    InMux I__5352 (
            .O(N__24582),
            .I(N__24554));
    Span4Mux_v I__5351 (
            .O(N__24579),
            .I(N__24547));
    Span4Mux_h I__5350 (
            .O(N__24576),
            .I(N__24547));
    LocalMux I__5349 (
            .O(N__24573),
            .I(N__24547));
    LocalMux I__5348 (
            .O(N__24570),
            .I(N__24544));
    InMux I__5347 (
            .O(N__24567),
            .I(N__24541));
    Sp12to4 I__5346 (
            .O(N__24562),
            .I(N__24538));
    Span4Mux_v I__5345 (
            .O(N__24557),
            .I(N__24533));
    LocalMux I__5344 (
            .O(N__24554),
            .I(N__24533));
    Span4Mux_v I__5343 (
            .O(N__24547),
            .I(N__24526));
    Span4Mux_v I__5342 (
            .O(N__24544),
            .I(N__24526));
    LocalMux I__5341 (
            .O(N__24541),
            .I(N__24526));
    Span12Mux_h I__5340 (
            .O(N__24538),
            .I(N__24521));
    Span4Mux_h I__5339 (
            .O(N__24533),
            .I(N__24516));
    Span4Mux_h I__5338 (
            .O(N__24526),
            .I(N__24516));
    InMux I__5337 (
            .O(N__24525),
            .I(N__24513));
    InMux I__5336 (
            .O(N__24524),
            .I(N__24510));
    Odrv12 I__5335 (
            .O(N__24521),
            .I(M_this_sprites_address_qZ0Z_8));
    Odrv4 I__5334 (
            .O(N__24516),
            .I(M_this_sprites_address_qZ0Z_8));
    LocalMux I__5333 (
            .O(N__24513),
            .I(M_this_sprites_address_qZ0Z_8));
    LocalMux I__5332 (
            .O(N__24510),
            .I(M_this_sprites_address_qZ0Z_8));
    InMux I__5331 (
            .O(N__24501),
            .I(N__24498));
    LocalMux I__5330 (
            .O(N__24498),
            .I(N_602));
    InMux I__5329 (
            .O(N__24495),
            .I(N__24491));
    InMux I__5328 (
            .O(N__24494),
            .I(N__24486));
    LocalMux I__5327 (
            .O(N__24491),
            .I(N__24480));
    InMux I__5326 (
            .O(N__24490),
            .I(N__24477));
    CascadeMux I__5325 (
            .O(N__24489),
            .I(N__24473));
    LocalMux I__5324 (
            .O(N__24486),
            .I(N__24470));
    InMux I__5323 (
            .O(N__24485),
            .I(N__24465));
    InMux I__5322 (
            .O(N__24484),
            .I(N__24465));
    InMux I__5321 (
            .O(N__24483),
            .I(N__24462));
    Span4Mux_v I__5320 (
            .O(N__24480),
            .I(N__24457));
    LocalMux I__5319 (
            .O(N__24477),
            .I(N__24457));
    InMux I__5318 (
            .O(N__24476),
            .I(N__24454));
    InMux I__5317 (
            .O(N__24473),
            .I(N__24451));
    Odrv4 I__5316 (
            .O(N__24470),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__5315 (
            .O(N__24465),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__5314 (
            .O(N__24462),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__5313 (
            .O(N__24457),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__5312 (
            .O(N__24454),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__5311 (
            .O(N__24451),
            .I(M_this_state_qZ0Z_9));
    InMux I__5310 (
            .O(N__24438),
            .I(N__24434));
    CascadeMux I__5309 (
            .O(N__24437),
            .I(N__24429));
    LocalMux I__5308 (
            .O(N__24434),
            .I(N__24426));
    InMux I__5307 (
            .O(N__24433),
            .I(N__24423));
    InMux I__5306 (
            .O(N__24432),
            .I(N__24418));
    InMux I__5305 (
            .O(N__24429),
            .I(N__24415));
    Span4Mux_h I__5304 (
            .O(N__24426),
            .I(N__24412));
    LocalMux I__5303 (
            .O(N__24423),
            .I(N__24409));
    InMux I__5302 (
            .O(N__24422),
            .I(N__24404));
    InMux I__5301 (
            .O(N__24421),
            .I(N__24404));
    LocalMux I__5300 (
            .O(N__24418),
            .I(N__24399));
    LocalMux I__5299 (
            .O(N__24415),
            .I(N__24399));
    Span4Mux_h I__5298 (
            .O(N__24412),
            .I(N__24396));
    Span4Mux_v I__5297 (
            .O(N__24409),
            .I(N__24393));
    LocalMux I__5296 (
            .O(N__24404),
            .I(M_this_state_qZ0Z_3));
    Odrv12 I__5295 (
            .O(N__24399),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__5294 (
            .O(N__24396),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__5293 (
            .O(N__24393),
            .I(M_this_state_qZ0Z_3));
    InMux I__5292 (
            .O(N__24384),
            .I(un1_M_this_sprites_address_q_cry_3));
    InMux I__5291 (
            .O(N__24381),
            .I(un1_M_this_sprites_address_q_cry_4));
    InMux I__5290 (
            .O(N__24378),
            .I(un1_M_this_sprites_address_q_cry_5));
    InMux I__5289 (
            .O(N__24375),
            .I(un1_M_this_sprites_address_q_cry_6));
    InMux I__5288 (
            .O(N__24372),
            .I(bfn_21_14_0_));
    InMux I__5287 (
            .O(N__24369),
            .I(un1_M_this_sprites_address_q_cry_8));
    CascadeMux I__5286 (
            .O(N__24366),
            .I(N__24361));
    CascadeMux I__5285 (
            .O(N__24365),
            .I(N__24358));
    CascadeMux I__5284 (
            .O(N__24364),
            .I(N__24353));
    InMux I__5283 (
            .O(N__24361),
            .I(N__24350));
    InMux I__5282 (
            .O(N__24358),
            .I(N__24347));
    CascadeMux I__5281 (
            .O(N__24357),
            .I(N__24344));
    CascadeMux I__5280 (
            .O(N__24356),
            .I(N__24340));
    InMux I__5279 (
            .O(N__24353),
            .I(N__24334));
    LocalMux I__5278 (
            .O(N__24350),
            .I(N__24329));
    LocalMux I__5277 (
            .O(N__24347),
            .I(N__24326));
    InMux I__5276 (
            .O(N__24344),
            .I(N__24323));
    CascadeMux I__5275 (
            .O(N__24343),
            .I(N__24320));
    InMux I__5274 (
            .O(N__24340),
            .I(N__24316));
    CascadeMux I__5273 (
            .O(N__24339),
            .I(N__24313));
    CascadeMux I__5272 (
            .O(N__24338),
            .I(N__24310));
    CascadeMux I__5271 (
            .O(N__24337),
            .I(N__24307));
    LocalMux I__5270 (
            .O(N__24334),
            .I(N__24304));
    CascadeMux I__5269 (
            .O(N__24333),
            .I(N__24301));
    CascadeMux I__5268 (
            .O(N__24332),
            .I(N__24298));
    Span4Mux_s3_v I__5267 (
            .O(N__24329),
            .I(N__24290));
    Span4Mux_h I__5266 (
            .O(N__24326),
            .I(N__24290));
    LocalMux I__5265 (
            .O(N__24323),
            .I(N__24290));
    InMux I__5264 (
            .O(N__24320),
            .I(N__24287));
    CascadeMux I__5263 (
            .O(N__24319),
            .I(N__24284));
    LocalMux I__5262 (
            .O(N__24316),
            .I(N__24280));
    InMux I__5261 (
            .O(N__24313),
            .I(N__24277));
    InMux I__5260 (
            .O(N__24310),
            .I(N__24274));
    InMux I__5259 (
            .O(N__24307),
            .I(N__24271));
    Span4Mux_v I__5258 (
            .O(N__24304),
            .I(N__24267));
    InMux I__5257 (
            .O(N__24301),
            .I(N__24264));
    InMux I__5256 (
            .O(N__24298),
            .I(N__24261));
    CascadeMux I__5255 (
            .O(N__24297),
            .I(N__24258));
    Span4Mux_v I__5254 (
            .O(N__24290),
            .I(N__24253));
    LocalMux I__5253 (
            .O(N__24287),
            .I(N__24253));
    InMux I__5252 (
            .O(N__24284),
            .I(N__24250));
    CascadeMux I__5251 (
            .O(N__24283),
            .I(N__24247));
    Span4Mux_h I__5250 (
            .O(N__24280),
            .I(N__24242));
    LocalMux I__5249 (
            .O(N__24277),
            .I(N__24242));
    LocalMux I__5248 (
            .O(N__24274),
            .I(N__24237));
    LocalMux I__5247 (
            .O(N__24271),
            .I(N__24237));
    CascadeMux I__5246 (
            .O(N__24270),
            .I(N__24234));
    Span4Mux_h I__5245 (
            .O(N__24267),
            .I(N__24227));
    LocalMux I__5244 (
            .O(N__24264),
            .I(N__24227));
    LocalMux I__5243 (
            .O(N__24261),
            .I(N__24227));
    InMux I__5242 (
            .O(N__24258),
            .I(N__24224));
    Span4Mux_h I__5241 (
            .O(N__24253),
            .I(N__24219));
    LocalMux I__5240 (
            .O(N__24250),
            .I(N__24219));
    InMux I__5239 (
            .O(N__24247),
            .I(N__24216));
    Span4Mux_v I__5238 (
            .O(N__24242),
            .I(N__24210));
    Span4Mux_v I__5237 (
            .O(N__24237),
            .I(N__24210));
    InMux I__5236 (
            .O(N__24234),
            .I(N__24207));
    Span4Mux_v I__5235 (
            .O(N__24227),
            .I(N__24198));
    LocalMux I__5234 (
            .O(N__24224),
            .I(N__24198));
    Span4Mux_v I__5233 (
            .O(N__24219),
            .I(N__24198));
    LocalMux I__5232 (
            .O(N__24216),
            .I(N__24198));
    CascadeMux I__5231 (
            .O(N__24215),
            .I(N__24195));
    Span4Mux_h I__5230 (
            .O(N__24210),
            .I(N__24191));
    LocalMux I__5229 (
            .O(N__24207),
            .I(N__24188));
    Span4Mux_v I__5228 (
            .O(N__24198),
            .I(N__24185));
    InMux I__5227 (
            .O(N__24195),
            .I(N__24182));
    InMux I__5226 (
            .O(N__24194),
            .I(N__24178));
    Sp12to4 I__5225 (
            .O(N__24191),
            .I(N__24173));
    Span12Mux_s11_h I__5224 (
            .O(N__24188),
            .I(N__24173));
    Sp12to4 I__5223 (
            .O(N__24185),
            .I(N__24168));
    LocalMux I__5222 (
            .O(N__24182),
            .I(N__24168));
    InMux I__5221 (
            .O(N__24181),
            .I(N__24165));
    LocalMux I__5220 (
            .O(N__24178),
            .I(N__24162));
    Odrv12 I__5219 (
            .O(N__24173),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv12 I__5218 (
            .O(N__24168),
            .I(M_this_sprites_address_qZ0Z_10));
    LocalMux I__5217 (
            .O(N__24165),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv4 I__5216 (
            .O(N__24162),
            .I(M_this_sprites_address_qZ0Z_10));
    InMux I__5215 (
            .O(N__24153),
            .I(N__24150));
    LocalMux I__5214 (
            .O(N__24150),
            .I(N__24147));
    Odrv4 I__5213 (
            .O(N__24147),
            .I(M_this_sprites_address_q_RNO_1Z0Z_10));
    InMux I__5212 (
            .O(N__24144),
            .I(un1_M_this_sprites_address_q_cry_9));
    InMux I__5211 (
            .O(N__24141),
            .I(N__24138));
    LocalMux I__5210 (
            .O(N__24138),
            .I(N__24135));
    Odrv4 I__5209 (
            .O(N__24135),
            .I(M_this_sprites_address_q_RNO_1Z0Z_11));
    InMux I__5208 (
            .O(N__24132),
            .I(un1_M_this_sprites_address_q_cry_10));
    InMux I__5207 (
            .O(N__24129),
            .I(un1_M_this_sprites_address_q_cry_11));
    InMux I__5206 (
            .O(N__24126),
            .I(N__24123));
    LocalMux I__5205 (
            .O(N__24123),
            .I(N__24120));
    Span4Mux_h I__5204 (
            .O(N__24120),
            .I(N__24117));
    Span4Mux_v I__5203 (
            .O(N__24117),
            .I(N__24114));
    Odrv4 I__5202 (
            .O(N__24114),
            .I(\this_sprites_ram.mem_out_bus6_1 ));
    InMux I__5201 (
            .O(N__24111),
            .I(N__24108));
    LocalMux I__5200 (
            .O(N__24108),
            .I(N__24105));
    Span4Mux_v I__5199 (
            .O(N__24105),
            .I(N__24102));
    Odrv4 I__5198 (
            .O(N__24102),
            .I(\this_sprites_ram.mem_out_bus2_1 ));
    InMux I__5197 (
            .O(N__24099),
            .I(N__24096));
    LocalMux I__5196 (
            .O(N__24096),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ));
    InMux I__5195 (
            .O(N__24093),
            .I(N__24090));
    LocalMux I__5194 (
            .O(N__24090),
            .I(N__24087));
    Span4Mux_v I__5193 (
            .O(N__24087),
            .I(N__24084));
    Odrv4 I__5192 (
            .O(N__24084),
            .I(\this_sprites_ram.mem_out_bus5_2 ));
    InMux I__5191 (
            .O(N__24081),
            .I(N__24078));
    LocalMux I__5190 (
            .O(N__24078),
            .I(N__24075));
    Span4Mux_h I__5189 (
            .O(N__24075),
            .I(N__24072));
    Odrv4 I__5188 (
            .O(N__24072),
            .I(\this_sprites_ram.mem_out_bus1_2 ));
    InMux I__5187 (
            .O(N__24069),
            .I(N__24066));
    LocalMux I__5186 (
            .O(N__24066),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ));
    CascadeMux I__5185 (
            .O(N__24063),
            .I(N__24060));
    InMux I__5184 (
            .O(N__24060),
            .I(N__24057));
    LocalMux I__5183 (
            .O(N__24057),
            .I(N__24054));
    Span4Mux_v I__5182 (
            .O(N__24054),
            .I(N__24051));
    Odrv4 I__5181 (
            .O(N__24051),
            .I(\this_sprites_ram.mem_out_bus5_0 ));
    InMux I__5180 (
            .O(N__24048),
            .I(N__24045));
    LocalMux I__5179 (
            .O(N__24045),
            .I(N__24042));
    Span4Mux_v I__5178 (
            .O(N__24042),
            .I(N__24039));
    Span4Mux_h I__5177 (
            .O(N__24039),
            .I(N__24036));
    Odrv4 I__5176 (
            .O(N__24036),
            .I(\this_sprites_ram.mem_out_bus1_0 ));
    InMux I__5175 (
            .O(N__24033),
            .I(N__24030));
    LocalMux I__5174 (
            .O(N__24030),
            .I(N__24027));
    Odrv4 I__5173 (
            .O(N__24027),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ));
    InMux I__5172 (
            .O(N__24024),
            .I(N__24021));
    LocalMux I__5171 (
            .O(N__24021),
            .I(M_this_sprites_address_qc_0_0));
    CEMux I__5170 (
            .O(N__24018),
            .I(N__24014));
    CEMux I__5169 (
            .O(N__24017),
            .I(N__24011));
    LocalMux I__5168 (
            .O(N__24014),
            .I(N__24008));
    LocalMux I__5167 (
            .O(N__24011),
            .I(N__24005));
    Span4Mux_s3_v I__5166 (
            .O(N__24008),
            .I(N__24002));
    Span4Mux_h I__5165 (
            .O(N__24005),
            .I(N__23999));
    Span4Mux_v I__5164 (
            .O(N__24002),
            .I(N__23994));
    Span4Mux_v I__5163 (
            .O(N__23999),
            .I(N__23994));
    Span4Mux_h I__5162 (
            .O(N__23994),
            .I(N__23991));
    Odrv4 I__5161 (
            .O(N__23991),
            .I(\this_sprites_ram.mem_WE_14 ));
    CascadeMux I__5160 (
            .O(N__23988),
            .I(N__23981));
    CascadeMux I__5159 (
            .O(N__23987),
            .I(N__23978));
    CascadeMux I__5158 (
            .O(N__23986),
            .I(N__23973));
    CascadeMux I__5157 (
            .O(N__23985),
            .I(N__23968));
    CascadeMux I__5156 (
            .O(N__23984),
            .I(N__23965));
    InMux I__5155 (
            .O(N__23981),
            .I(N__23960));
    InMux I__5154 (
            .O(N__23978),
            .I(N__23957));
    CascadeMux I__5153 (
            .O(N__23977),
            .I(N__23954));
    CascadeMux I__5152 (
            .O(N__23976),
            .I(N__23951));
    InMux I__5151 (
            .O(N__23973),
            .I(N__23945));
    CascadeMux I__5150 (
            .O(N__23972),
            .I(N__23942));
    CascadeMux I__5149 (
            .O(N__23971),
            .I(N__23939));
    InMux I__5148 (
            .O(N__23968),
            .I(N__23935));
    InMux I__5147 (
            .O(N__23965),
            .I(N__23932));
    CascadeMux I__5146 (
            .O(N__23964),
            .I(N__23929));
    CascadeMux I__5145 (
            .O(N__23963),
            .I(N__23926));
    LocalMux I__5144 (
            .O(N__23960),
            .I(N__23920));
    LocalMux I__5143 (
            .O(N__23957),
            .I(N__23920));
    InMux I__5142 (
            .O(N__23954),
            .I(N__23917));
    InMux I__5141 (
            .O(N__23951),
            .I(N__23914));
    CascadeMux I__5140 (
            .O(N__23950),
            .I(N__23911));
    CascadeMux I__5139 (
            .O(N__23949),
            .I(N__23908));
    CascadeMux I__5138 (
            .O(N__23948),
            .I(N__23905));
    LocalMux I__5137 (
            .O(N__23945),
            .I(N__23902));
    InMux I__5136 (
            .O(N__23942),
            .I(N__23899));
    InMux I__5135 (
            .O(N__23939),
            .I(N__23896));
    CascadeMux I__5134 (
            .O(N__23938),
            .I(N__23893));
    LocalMux I__5133 (
            .O(N__23935),
            .I(N__23890));
    LocalMux I__5132 (
            .O(N__23932),
            .I(N__23887));
    InMux I__5131 (
            .O(N__23929),
            .I(N__23884));
    InMux I__5130 (
            .O(N__23926),
            .I(N__23881));
    CascadeMux I__5129 (
            .O(N__23925),
            .I(N__23878));
    Span4Mux_v I__5128 (
            .O(N__23920),
            .I(N__23871));
    LocalMux I__5127 (
            .O(N__23917),
            .I(N__23871));
    LocalMux I__5126 (
            .O(N__23914),
            .I(N__23871));
    InMux I__5125 (
            .O(N__23911),
            .I(N__23868));
    InMux I__5124 (
            .O(N__23908),
            .I(N__23865));
    InMux I__5123 (
            .O(N__23905),
            .I(N__23862));
    Span4Mux_v I__5122 (
            .O(N__23902),
            .I(N__23855));
    LocalMux I__5121 (
            .O(N__23899),
            .I(N__23855));
    LocalMux I__5120 (
            .O(N__23896),
            .I(N__23855));
    InMux I__5119 (
            .O(N__23893),
            .I(N__23852));
    Span4Mux_v I__5118 (
            .O(N__23890),
            .I(N__23845));
    Span4Mux_h I__5117 (
            .O(N__23887),
            .I(N__23845));
    LocalMux I__5116 (
            .O(N__23884),
            .I(N__23845));
    LocalMux I__5115 (
            .O(N__23881),
            .I(N__23842));
    InMux I__5114 (
            .O(N__23878),
            .I(N__23839));
    Span4Mux_v I__5113 (
            .O(N__23871),
            .I(N__23832));
    LocalMux I__5112 (
            .O(N__23868),
            .I(N__23832));
    LocalMux I__5111 (
            .O(N__23865),
            .I(N__23832));
    LocalMux I__5110 (
            .O(N__23862),
            .I(N__23825));
    Span4Mux_v I__5109 (
            .O(N__23855),
            .I(N__23825));
    LocalMux I__5108 (
            .O(N__23852),
            .I(N__23825));
    Span4Mux_v I__5107 (
            .O(N__23845),
            .I(N__23819));
    Span4Mux_h I__5106 (
            .O(N__23842),
            .I(N__23819));
    LocalMux I__5105 (
            .O(N__23839),
            .I(N__23816));
    Span4Mux_v I__5104 (
            .O(N__23832),
            .I(N__23811));
    Span4Mux_v I__5103 (
            .O(N__23825),
            .I(N__23811));
    InMux I__5102 (
            .O(N__23824),
            .I(N__23808));
    Span4Mux_h I__5101 (
            .O(N__23819),
            .I(N__23805));
    Span4Mux_h I__5100 (
            .O(N__23816),
            .I(N__23802));
    Span4Mux_h I__5099 (
            .O(N__23811),
            .I(N__23796));
    LocalMux I__5098 (
            .O(N__23808),
            .I(N__23796));
    Span4Mux_h I__5097 (
            .O(N__23805),
            .I(N__23793));
    Span4Mux_h I__5096 (
            .O(N__23802),
            .I(N__23790));
    InMux I__5095 (
            .O(N__23801),
            .I(N__23787));
    Span4Mux_h I__5094 (
            .O(N__23796),
            .I(N__23784));
    Odrv4 I__5093 (
            .O(N__23793),
            .I(M_this_sprites_address_qZ0Z_0));
    Odrv4 I__5092 (
            .O(N__23790),
            .I(M_this_sprites_address_qZ0Z_0));
    LocalMux I__5091 (
            .O(N__23787),
            .I(M_this_sprites_address_qZ0Z_0));
    Odrv4 I__5090 (
            .O(N__23784),
            .I(M_this_sprites_address_qZ0Z_0));
    CascadeMux I__5089 (
            .O(N__23775),
            .I(N__23771));
    InMux I__5088 (
            .O(N__23774),
            .I(N__23768));
    InMux I__5087 (
            .O(N__23771),
            .I(N__23765));
    LocalMux I__5086 (
            .O(N__23768),
            .I(N_443_i));
    LocalMux I__5085 (
            .O(N__23765),
            .I(N_443_i));
    InMux I__5084 (
            .O(N__23760),
            .I(N__23757));
    LocalMux I__5083 (
            .O(N__23757),
            .I(N__23754));
    Span4Mux_v I__5082 (
            .O(N__23754),
            .I(N__23751));
    Span4Mux_h I__5081 (
            .O(N__23751),
            .I(N__23748));
    Odrv4 I__5080 (
            .O(N__23748),
            .I(M_this_sprites_address_q_RNO_0Z0Z_0));
    InMux I__5079 (
            .O(N__23745),
            .I(un1_M_this_sprites_address_q_cry_0));
    InMux I__5078 (
            .O(N__23742),
            .I(un1_M_this_sprites_address_q_cry_1));
    InMux I__5077 (
            .O(N__23739),
            .I(un1_M_this_sprites_address_q_cry_2));
    InMux I__5076 (
            .O(N__23736),
            .I(bfn_20_20_0_));
    CascadeMux I__5075 (
            .O(N__23733),
            .I(N__23730));
    InMux I__5074 (
            .O(N__23730),
            .I(N__23727));
    LocalMux I__5073 (
            .O(N__23727),
            .I(\this_ppu.un1_M_vaddress_q_cry_7_THRU_CO ));
    CascadeMux I__5072 (
            .O(N__23724),
            .I(N__23721));
    InMux I__5071 (
            .O(N__23721),
            .I(N__23718));
    LocalMux I__5070 (
            .O(N__23718),
            .I(N__23715));
    Span4Mux_h I__5069 (
            .O(N__23715),
            .I(N__23712));
    Span4Mux_v I__5068 (
            .O(N__23712),
            .I(N__23709));
    Span4Mux_h I__5067 (
            .O(N__23709),
            .I(N__23706));
    Span4Mux_h I__5066 (
            .O(N__23706),
            .I(N__23703));
    Odrv4 I__5065 (
            .O(N__23703),
            .I(M_this_map_ram_read_data_5));
    CascadeMux I__5064 (
            .O(N__23700),
            .I(N__23692));
    InMux I__5063 (
            .O(N__23699),
            .I(N__23688));
    InMux I__5062 (
            .O(N__23698),
            .I(N__23685));
    InMux I__5061 (
            .O(N__23697),
            .I(N__23682));
    InMux I__5060 (
            .O(N__23696),
            .I(N__23678));
    InMux I__5059 (
            .O(N__23695),
            .I(N__23675));
    InMux I__5058 (
            .O(N__23692),
            .I(N__23670));
    InMux I__5057 (
            .O(N__23691),
            .I(N__23670));
    LocalMux I__5056 (
            .O(N__23688),
            .I(N__23663));
    LocalMux I__5055 (
            .O(N__23685),
            .I(N__23663));
    LocalMux I__5054 (
            .O(N__23682),
            .I(N__23663));
    InMux I__5053 (
            .O(N__23681),
            .I(N__23660));
    LocalMux I__5052 (
            .O(N__23678),
            .I(N__23653));
    LocalMux I__5051 (
            .O(N__23675),
            .I(N__23653));
    LocalMux I__5050 (
            .O(N__23670),
            .I(N__23653));
    Sp12to4 I__5049 (
            .O(N__23663),
            .I(N__23646));
    LocalMux I__5048 (
            .O(N__23660),
            .I(N__23646));
    Sp12to4 I__5047 (
            .O(N__23653),
            .I(N__23646));
    Odrv12 I__5046 (
            .O(N__23646),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    InMux I__5045 (
            .O(N__23643),
            .I(N__23640));
    LocalMux I__5044 (
            .O(N__23640),
            .I(N__23635));
    InMux I__5043 (
            .O(N__23639),
            .I(N__23632));
    CascadeMux I__5042 (
            .O(N__23638),
            .I(N__23629));
    Span4Mux_v I__5041 (
            .O(N__23635),
            .I(N__23624));
    LocalMux I__5040 (
            .O(N__23632),
            .I(N__23624));
    InMux I__5039 (
            .O(N__23629),
            .I(N__23621));
    Span4Mux_v I__5038 (
            .O(N__23624),
            .I(N__23612));
    LocalMux I__5037 (
            .O(N__23621),
            .I(N__23612));
    CascadeMux I__5036 (
            .O(N__23620),
            .I(N__23609));
    InMux I__5035 (
            .O(N__23619),
            .I(N__23601));
    InMux I__5034 (
            .O(N__23618),
            .I(N__23601));
    InMux I__5033 (
            .O(N__23617),
            .I(N__23601));
    Span4Mux_v I__5032 (
            .O(N__23612),
            .I(N__23598));
    InMux I__5031 (
            .O(N__23609),
            .I(N__23595));
    InMux I__5030 (
            .O(N__23608),
            .I(N__23592));
    LocalMux I__5029 (
            .O(N__23601),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__5028 (
            .O(N__23598),
            .I(M_this_state_qZ0Z_13));
    LocalMux I__5027 (
            .O(N__23595),
            .I(M_this_state_qZ0Z_13));
    LocalMux I__5026 (
            .O(N__23592),
            .I(M_this_state_qZ0Z_13));
    InMux I__5025 (
            .O(N__23583),
            .I(N__23571));
    InMux I__5024 (
            .O(N__23582),
            .I(N__23571));
    InMux I__5023 (
            .O(N__23581),
            .I(N__23571));
    InMux I__5022 (
            .O(N__23580),
            .I(N__23571));
    LocalMux I__5021 (
            .O(N__23571),
            .I(M_this_delay_clk_out_0));
    InMux I__5020 (
            .O(N__23568),
            .I(N__23564));
    InMux I__5019 (
            .O(N__23567),
            .I(N__23561));
    LocalMux I__5018 (
            .O(N__23564),
            .I(N__23558));
    LocalMux I__5017 (
            .O(N__23561),
            .I(\this_ppu.M_this_ppu_vram_addr_i_7 ));
    Odrv4 I__5016 (
            .O(N__23558),
            .I(\this_ppu.M_this_ppu_vram_addr_i_7 ));
    InMux I__5015 (
            .O(N__23553),
            .I(N__23549));
    InMux I__5014 (
            .O(N__23552),
            .I(N__23546));
    LocalMux I__5013 (
            .O(N__23549),
            .I(N__23543));
    LocalMux I__5012 (
            .O(N__23546),
            .I(\this_ppu.M_vaddress_q_i_1 ));
    Odrv4 I__5011 (
            .O(N__23543),
            .I(\this_ppu.M_vaddress_q_i_1 ));
    InMux I__5010 (
            .O(N__23538),
            .I(N__23534));
    InMux I__5009 (
            .O(N__23537),
            .I(N__23531));
    LocalMux I__5008 (
            .O(N__23534),
            .I(N__23528));
    LocalMux I__5007 (
            .O(N__23531),
            .I(\this_ppu.M_vaddress_q_i_2 ));
    Odrv4 I__5006 (
            .O(N__23528),
            .I(\this_ppu.M_vaddress_q_i_2 ));
    CascadeMux I__5005 (
            .O(N__23523),
            .I(N__23520));
    InMux I__5004 (
            .O(N__23520),
            .I(N__23516));
    InMux I__5003 (
            .O(N__23519),
            .I(N__23513));
    LocalMux I__5002 (
            .O(N__23516),
            .I(N__23510));
    LocalMux I__5001 (
            .O(N__23513),
            .I(\this_ppu.M_this_ppu_map_addr_i_5 ));
    Odrv4 I__5000 (
            .O(N__23510),
            .I(\this_ppu.M_this_ppu_map_addr_i_5 ));
    CascadeMux I__4999 (
            .O(N__23505),
            .I(N__23502));
    InMux I__4998 (
            .O(N__23502),
            .I(N__23498));
    InMux I__4997 (
            .O(N__23501),
            .I(N__23495));
    LocalMux I__4996 (
            .O(N__23498),
            .I(N__23492));
    LocalMux I__4995 (
            .O(N__23495),
            .I(\this_ppu.M_this_ppu_map_addr_i_6 ));
    Odrv4 I__4994 (
            .O(N__23492),
            .I(\this_ppu.M_this_ppu_map_addr_i_6 ));
    CascadeMux I__4993 (
            .O(N__23487),
            .I(N__23484));
    InMux I__4992 (
            .O(N__23484),
            .I(N__23480));
    InMux I__4991 (
            .O(N__23483),
            .I(N__23477));
    LocalMux I__4990 (
            .O(N__23480),
            .I(N__23474));
    LocalMux I__4989 (
            .O(N__23477),
            .I(\this_ppu.M_this_ppu_map_addr_i_7 ));
    Odrv4 I__4988 (
            .O(N__23474),
            .I(\this_ppu.M_this_ppu_map_addr_i_7 ));
    CascadeMux I__4987 (
            .O(N__23469),
            .I(N__23466));
    InMux I__4986 (
            .O(N__23466),
            .I(N__23462));
    InMux I__4985 (
            .O(N__23465),
            .I(N__23459));
    LocalMux I__4984 (
            .O(N__23462),
            .I(N__23456));
    LocalMux I__4983 (
            .O(N__23459),
            .I(\this_ppu.M_this_ppu_map_addr_i_8 ));
    Odrv4 I__4982 (
            .O(N__23456),
            .I(\this_ppu.M_this_ppu_map_addr_i_8 ));
    CascadeMux I__4981 (
            .O(N__23451),
            .I(N__23447));
    InMux I__4980 (
            .O(N__23450),
            .I(N__23444));
    InMux I__4979 (
            .O(N__23447),
            .I(N__23441));
    LocalMux I__4978 (
            .O(N__23444),
            .I(N__23438));
    LocalMux I__4977 (
            .O(N__23441),
            .I(\this_ppu.M_this_ppu_map_addr_i_9 ));
    Odrv4 I__4976 (
            .O(N__23438),
            .I(\this_ppu.M_this_ppu_map_addr_i_9 ));
    CascadeMux I__4975 (
            .O(N__23433),
            .I(N__23425));
    InMux I__4974 (
            .O(N__23432),
            .I(N__23422));
    InMux I__4973 (
            .O(N__23431),
            .I(N__23419));
    InMux I__4972 (
            .O(N__23430),
            .I(N__23416));
    InMux I__4971 (
            .O(N__23429),
            .I(N__23411));
    InMux I__4970 (
            .O(N__23428),
            .I(N__23411));
    InMux I__4969 (
            .O(N__23425),
            .I(N__23408));
    LocalMux I__4968 (
            .O(N__23422),
            .I(N__23405));
    LocalMux I__4967 (
            .O(N__23419),
            .I(N__23398));
    LocalMux I__4966 (
            .O(N__23416),
            .I(N__23398));
    LocalMux I__4965 (
            .O(N__23411),
            .I(N__23398));
    LocalMux I__4964 (
            .O(N__23408),
            .I(N__23395));
    Span4Mux_h I__4963 (
            .O(N__23405),
            .I(N__23392));
    Span4Mux_h I__4962 (
            .O(N__23398),
            .I(N__23389));
    Odrv12 I__4961 (
            .O(N__23395),
            .I(N_775_0));
    Odrv4 I__4960 (
            .O(N__23392),
            .I(N_775_0));
    Odrv4 I__4959 (
            .O(N__23389),
            .I(N_775_0));
    CascadeMux I__4958 (
            .O(N__23382),
            .I(N_775_0_cascade_));
    InMux I__4957 (
            .O(N__23379),
            .I(N__23376));
    LocalMux I__4956 (
            .O(N__23376),
            .I(N__23373));
    Span4Mux_h I__4955 (
            .O(N__23373),
            .I(N__23370));
    Span4Mux_v I__4954 (
            .O(N__23370),
            .I(N__23367));
    Sp12to4 I__4953 (
            .O(N__23367),
            .I(N__23364));
    Odrv12 I__4952 (
            .O(N__23364),
            .I(port_address_in_5));
    InMux I__4951 (
            .O(N__23361),
            .I(N__23355));
    InMux I__4950 (
            .O(N__23360),
            .I(N__23355));
    LocalMux I__4949 (
            .O(N__23355),
            .I(N__23352));
    Odrv12 I__4948 (
            .O(N__23352),
            .I(\this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0Z0Z_0 ));
    CascadeMux I__4947 (
            .O(N__23349),
            .I(N_87_0_cascade_));
    CascadeMux I__4946 (
            .O(N__23346),
            .I(N__23339));
    CascadeMux I__4945 (
            .O(N__23345),
            .I(N__23336));
    CascadeMux I__4944 (
            .O(N__23344),
            .I(N__23333));
    CascadeMux I__4943 (
            .O(N__23343),
            .I(N__23330));
    InMux I__4942 (
            .O(N__23342),
            .I(N__23327));
    InMux I__4941 (
            .O(N__23339),
            .I(N__23324));
    InMux I__4940 (
            .O(N__23336),
            .I(N__23321));
    InMux I__4939 (
            .O(N__23333),
            .I(N__23316));
    InMux I__4938 (
            .O(N__23330),
            .I(N__23316));
    LocalMux I__4937 (
            .O(N__23327),
            .I(N__23312));
    LocalMux I__4936 (
            .O(N__23324),
            .I(N__23309));
    LocalMux I__4935 (
            .O(N__23321),
            .I(N__23304));
    LocalMux I__4934 (
            .O(N__23316),
            .I(N__23304));
    InMux I__4933 (
            .O(N__23315),
            .I(N__23301));
    Span4Mux_v I__4932 (
            .O(N__23312),
            .I(N__23294));
    Span4Mux_h I__4931 (
            .O(N__23309),
            .I(N__23294));
    Span4Mux_v I__4930 (
            .O(N__23304),
            .I(N__23294));
    LocalMux I__4929 (
            .O(N__23301),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__4928 (
            .O(N__23294),
            .I(M_this_state_qZ0Z_6));
    CascadeMux I__4927 (
            .O(N__23289),
            .I(N__23286));
    InMux I__4926 (
            .O(N__23286),
            .I(N__23274));
    InMux I__4925 (
            .O(N__23285),
            .I(N__23274));
    InMux I__4924 (
            .O(N__23284),
            .I(N__23274));
    InMux I__4923 (
            .O(N__23283),
            .I(N__23274));
    LocalMux I__4922 (
            .O(N__23274),
            .I(N__23271));
    Span4Mux_v I__4921 (
            .O(N__23271),
            .I(N__23268));
    Span4Mux_h I__4920 (
            .O(N__23268),
            .I(N__23265));
    Span4Mux_h I__4919 (
            .O(N__23265),
            .I(N__23262));
    Sp12to4 I__4918 (
            .O(N__23262),
            .I(N__23259));
    Span12Mux_h I__4917 (
            .O(N__23259),
            .I(N__23256));
    Odrv12 I__4916 (
            .O(N__23256),
            .I(port_enb_c));
    InMux I__4915 (
            .O(N__23253),
            .I(N__23250));
    LocalMux I__4914 (
            .O(N__23250),
            .I(N__23247));
    Span4Mux_v I__4913 (
            .O(N__23247),
            .I(N__23241));
    InMux I__4912 (
            .O(N__23246),
            .I(N__23234));
    InMux I__4911 (
            .O(N__23245),
            .I(N__23234));
    InMux I__4910 (
            .O(N__23244),
            .I(N__23234));
    Odrv4 I__4909 (
            .O(N__23241),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__4908 (
            .O(N__23234),
            .I(this_start_data_delay_M_last_q));
    InMux I__4907 (
            .O(N__23229),
            .I(N__23226));
    LocalMux I__4906 (
            .O(N__23226),
            .I(\this_reset_cond.M_stage_qZ0Z_4 ));
    InMux I__4905 (
            .O(N__23223),
            .I(N__23218));
    InMux I__4904 (
            .O(N__23222),
            .I(N__23214));
    InMux I__4903 (
            .O(N__23221),
            .I(N__23211));
    LocalMux I__4902 (
            .O(N__23218),
            .I(N__23207));
    InMux I__4901 (
            .O(N__23217),
            .I(N__23204));
    LocalMux I__4900 (
            .O(N__23214),
            .I(N__23197));
    LocalMux I__4899 (
            .O(N__23211),
            .I(N__23197));
    InMux I__4898 (
            .O(N__23210),
            .I(N__23194));
    Span4Mux_v I__4897 (
            .O(N__23207),
            .I(N__23189));
    LocalMux I__4896 (
            .O(N__23204),
            .I(N__23189));
    InMux I__4895 (
            .O(N__23203),
            .I(N__23186));
    InMux I__4894 (
            .O(N__23202),
            .I(N__23183));
    Span4Mux_h I__4893 (
            .O(N__23197),
            .I(N__23180));
    LocalMux I__4892 (
            .O(N__23194),
            .I(N__23175));
    Span4Mux_h I__4891 (
            .O(N__23189),
            .I(N__23175));
    LocalMux I__4890 (
            .O(N__23186),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__4889 (
            .O(N__23183),
            .I(M_this_state_qZ0Z_11));
    Odrv4 I__4888 (
            .O(N__23180),
            .I(M_this_state_qZ0Z_11));
    Odrv4 I__4887 (
            .O(N__23175),
            .I(M_this_state_qZ0Z_11));
    InMux I__4886 (
            .O(N__23166),
            .I(N__23163));
    LocalMux I__4885 (
            .O(N__23163),
            .I(N__23160));
    Odrv12 I__4884 (
            .O(N__23160),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    CascadeMux I__4883 (
            .O(N__23157),
            .I(N__23154));
    InMux I__4882 (
            .O(N__23154),
            .I(N__23151));
    LocalMux I__4881 (
            .O(N__23151),
            .I(N_126));
    InMux I__4880 (
            .O(N__23148),
            .I(N__23145));
    LocalMux I__4879 (
            .O(N__23145),
            .I(N__23141));
    InMux I__4878 (
            .O(N__23144),
            .I(N__23134));
    Span4Mux_h I__4877 (
            .O(N__23141),
            .I(N__23131));
    InMux I__4876 (
            .O(N__23140),
            .I(N__23124));
    InMux I__4875 (
            .O(N__23139),
            .I(N__23124));
    InMux I__4874 (
            .O(N__23138),
            .I(N__23124));
    InMux I__4873 (
            .O(N__23137),
            .I(N__23121));
    LocalMux I__4872 (
            .O(N__23134),
            .I(N__23118));
    Odrv4 I__4871 (
            .O(N__23131),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__4870 (
            .O(N__23124),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__4869 (
            .O(N__23121),
            .I(M_this_state_qZ0Z_7));
    Odrv12 I__4868 (
            .O(N__23118),
            .I(M_this_state_qZ0Z_7));
    CascadeMux I__4867 (
            .O(N__23109),
            .I(port_dmab_ac0_1_3_cascade_));
    InMux I__4866 (
            .O(N__23106),
            .I(N__23103));
    LocalMux I__4865 (
            .O(N__23103),
            .I(port_dmab_ac0_1_4));
    InMux I__4864 (
            .O(N__23100),
            .I(N__23096));
    InMux I__4863 (
            .O(N__23099),
            .I(N__23092));
    LocalMux I__4862 (
            .O(N__23096),
            .I(N__23087));
    InMux I__4861 (
            .O(N__23095),
            .I(N__23084));
    LocalMux I__4860 (
            .O(N__23092),
            .I(N__23081));
    InMux I__4859 (
            .O(N__23091),
            .I(N__23078));
    InMux I__4858 (
            .O(N__23090),
            .I(N__23074));
    Span4Mux_h I__4857 (
            .O(N__23087),
            .I(N__23069));
    LocalMux I__4856 (
            .O(N__23084),
            .I(N__23066));
    Span4Mux_v I__4855 (
            .O(N__23081),
            .I(N__23061));
    LocalMux I__4854 (
            .O(N__23078),
            .I(N__23061));
    InMux I__4853 (
            .O(N__23077),
            .I(N__23058));
    LocalMux I__4852 (
            .O(N__23074),
            .I(N__23055));
    InMux I__4851 (
            .O(N__23073),
            .I(N__23052));
    InMux I__4850 (
            .O(N__23072),
            .I(N__23049));
    Span4Mux_v I__4849 (
            .O(N__23069),
            .I(N__23044));
    Span4Mux_h I__4848 (
            .O(N__23066),
            .I(N__23044));
    Span4Mux_v I__4847 (
            .O(N__23061),
            .I(N__23039));
    LocalMux I__4846 (
            .O(N__23058),
            .I(N__23039));
    Span4Mux_h I__4845 (
            .O(N__23055),
            .I(N__23036));
    LocalMux I__4844 (
            .O(N__23052),
            .I(N__23033));
    LocalMux I__4843 (
            .O(N__23049),
            .I(N__23030));
    Span4Mux_v I__4842 (
            .O(N__23044),
            .I(N__23027));
    Sp12to4 I__4841 (
            .O(N__23039),
            .I(N__23024));
    Span4Mux_v I__4840 (
            .O(N__23036),
            .I(N__23019));
    Span4Mux_h I__4839 (
            .O(N__23033),
            .I(N__23019));
    Span4Mux_h I__4838 (
            .O(N__23030),
            .I(N__23016));
    Span4Mux_h I__4837 (
            .O(N__23027),
            .I(N__23013));
    Span12Mux_v I__4836 (
            .O(N__23024),
            .I(N__23010));
    Span4Mux_h I__4835 (
            .O(N__23019),
            .I(N__23005));
    Span4Mux_h I__4834 (
            .O(N__23016),
            .I(N__23005));
    Odrv4 I__4833 (
            .O(N__23013),
            .I(N_15));
    Odrv12 I__4832 (
            .O(N__23010),
            .I(N_15));
    Odrv4 I__4831 (
            .O(N__23005),
            .I(N_15));
    CascadeMux I__4830 (
            .O(N__22998),
            .I(N_809_cascade_));
    InMux I__4829 (
            .O(N__22995),
            .I(N__22988));
    InMux I__4828 (
            .O(N__22994),
            .I(N__22985));
    InMux I__4827 (
            .O(N__22993),
            .I(N__22982));
    CascadeMux I__4826 (
            .O(N__22992),
            .I(N__22978));
    InMux I__4825 (
            .O(N__22991),
            .I(N__22975));
    LocalMux I__4824 (
            .O(N__22988),
            .I(N__22972));
    LocalMux I__4823 (
            .O(N__22985),
            .I(N__22969));
    LocalMux I__4822 (
            .O(N__22982),
            .I(N__22966));
    InMux I__4821 (
            .O(N__22981),
            .I(N__22963));
    InMux I__4820 (
            .O(N__22978),
            .I(N__22960));
    LocalMux I__4819 (
            .O(N__22975),
            .I(N__22957));
    Span12Mux_h I__4818 (
            .O(N__22972),
            .I(N__22954));
    Span4Mux_h I__4817 (
            .O(N__22969),
            .I(N__22949));
    Span4Mux_h I__4816 (
            .O(N__22966),
            .I(N__22949));
    LocalMux I__4815 (
            .O(N__22963),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__4814 (
            .O(N__22960),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__4813 (
            .O(N__22957),
            .I(M_this_state_qZ0Z_5));
    Odrv12 I__4812 (
            .O(N__22954),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__4811 (
            .O(N__22949),
            .I(M_this_state_qZ0Z_5));
    InMux I__4810 (
            .O(N__22938),
            .I(N__22934));
    InMux I__4809 (
            .O(N__22937),
            .I(N__22931));
    LocalMux I__4808 (
            .O(N__22934),
            .I(N__22925));
    LocalMux I__4807 (
            .O(N__22931),
            .I(N__22922));
    InMux I__4806 (
            .O(N__22930),
            .I(N__22919));
    InMux I__4805 (
            .O(N__22929),
            .I(N__22916));
    InMux I__4804 (
            .O(N__22928),
            .I(N__22913));
    Span4Mux_h I__4803 (
            .O(N__22925),
            .I(N__22910));
    Span4Mux_h I__4802 (
            .O(N__22922),
            .I(N__22907));
    LocalMux I__4801 (
            .O(N__22919),
            .I(N__22902));
    LocalMux I__4800 (
            .O(N__22916),
            .I(N__22902));
    LocalMux I__4799 (
            .O(N__22913),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__4798 (
            .O(N__22910),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__4797 (
            .O(N__22907),
            .I(M_this_state_qZ0Z_8));
    Odrv12 I__4796 (
            .O(N__22902),
            .I(M_this_state_qZ0Z_8));
    InMux I__4795 (
            .O(N__22893),
            .I(N__22889));
    InMux I__4794 (
            .O(N__22892),
            .I(N__22886));
    LocalMux I__4793 (
            .O(N__22889),
            .I(N__22883));
    LocalMux I__4792 (
            .O(N__22886),
            .I(N__22878));
    Span4Mux_h I__4791 (
            .O(N__22883),
            .I(N__22875));
    InMux I__4790 (
            .O(N__22882),
            .I(N__22870));
    InMux I__4789 (
            .O(N__22881),
            .I(N__22870));
    Odrv12 I__4788 (
            .O(N__22878),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__4787 (
            .O(N__22875),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__4786 (
            .O(N__22870),
            .I(M_this_state_qZ0Z_1));
    CascadeMux I__4785 (
            .O(N__22863),
            .I(N__22860));
    InMux I__4784 (
            .O(N__22860),
            .I(N__22857));
    LocalMux I__4783 (
            .O(N__22857),
            .I(N_792));
    InMux I__4782 (
            .O(N__22854),
            .I(N__22851));
    LocalMux I__4781 (
            .O(N__22851),
            .I(M_this_sprites_address_qc_0_0_0));
    CascadeMux I__4780 (
            .O(N__22848),
            .I(N__22845));
    InMux I__4779 (
            .O(N__22845),
            .I(N__22842));
    LocalMux I__4778 (
            .O(N__22842),
            .I(N_795));
    CascadeMux I__4777 (
            .O(N__22839),
            .I(N__22836));
    InMux I__4776 (
            .O(N__22836),
            .I(N__22833));
    LocalMux I__4775 (
            .O(N__22833),
            .I(N__22830));
    Odrv4 I__4774 (
            .O(N__22830),
            .I(N_773_0));
    CascadeMux I__4773 (
            .O(N__22827),
            .I(N_773_0_cascade_));
    InMux I__4772 (
            .O(N__22824),
            .I(N__22821));
    LocalMux I__4771 (
            .O(N__22821),
            .I(\this_vga_signals.N_485 ));
    InMux I__4770 (
            .O(N__22818),
            .I(N__22814));
    InMux I__4769 (
            .O(N__22817),
            .I(N__22808));
    LocalMux I__4768 (
            .O(N__22814),
            .I(N__22804));
    InMux I__4767 (
            .O(N__22813),
            .I(N__22801));
    InMux I__4766 (
            .O(N__22812),
            .I(N__22797));
    InMux I__4765 (
            .O(N__22811),
            .I(N__22794));
    LocalMux I__4764 (
            .O(N__22808),
            .I(N__22790));
    InMux I__4763 (
            .O(N__22807),
            .I(N__22787));
    Span4Mux_v I__4762 (
            .O(N__22804),
            .I(N__22782));
    LocalMux I__4761 (
            .O(N__22801),
            .I(N__22782));
    InMux I__4760 (
            .O(N__22800),
            .I(N__22779));
    LocalMux I__4759 (
            .O(N__22797),
            .I(N__22776));
    LocalMux I__4758 (
            .O(N__22794),
            .I(N__22773));
    InMux I__4757 (
            .O(N__22793),
            .I(N__22770));
    Sp12to4 I__4756 (
            .O(N__22790),
            .I(N__22765));
    LocalMux I__4755 (
            .O(N__22787),
            .I(N__22765));
    Span4Mux_v I__4754 (
            .O(N__22782),
            .I(N__22760));
    LocalMux I__4753 (
            .O(N__22779),
            .I(N__22760));
    Span4Mux_h I__4752 (
            .O(N__22776),
            .I(N__22757));
    Span4Mux_h I__4751 (
            .O(N__22773),
            .I(N__22754));
    LocalMux I__4750 (
            .O(N__22770),
            .I(N__22751));
    Span12Mux_v I__4749 (
            .O(N__22765),
            .I(N__22748));
    Span4Mux_v I__4748 (
            .O(N__22760),
            .I(N__22745));
    Span4Mux_v I__4747 (
            .O(N__22757),
            .I(N__22738));
    Span4Mux_v I__4746 (
            .O(N__22754),
            .I(N__22738));
    Span4Mux_h I__4745 (
            .O(N__22751),
            .I(N__22738));
    Span12Mux_h I__4744 (
            .O(N__22748),
            .I(N__22735));
    Span4Mux_h I__4743 (
            .O(N__22745),
            .I(N__22732));
    Span4Mux_h I__4742 (
            .O(N__22738),
            .I(N__22729));
    Odrv12 I__4741 (
            .O(N__22735),
            .I(N_17));
    Odrv4 I__4740 (
            .O(N__22732),
            .I(N_17));
    Odrv4 I__4739 (
            .O(N__22729),
            .I(N_17));
    InMux I__4738 (
            .O(N__22722),
            .I(N__22719));
    LocalMux I__4737 (
            .O(N__22719),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ));
    CascadeMux I__4736 (
            .O(N__22716),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ));
    InMux I__4735 (
            .O(N__22713),
            .I(N__22710));
    LocalMux I__4734 (
            .O(N__22710),
            .I(N__22707));
    Span12Mux_s9_v I__4733 (
            .O(N__22707),
            .I(N__22704));
    Span12Mux_h I__4732 (
            .O(N__22704),
            .I(N__22700));
    InMux I__4731 (
            .O(N__22703),
            .I(N__22697));
    Odrv12 I__4730 (
            .O(N__22700),
            .I(M_this_ppu_vram_data_1));
    LocalMux I__4729 (
            .O(N__22697),
            .I(M_this_ppu_vram_data_1));
    InMux I__4728 (
            .O(N__22692),
            .I(N__22689));
    LocalMux I__4727 (
            .O(N__22689),
            .I(N__22686));
    Span4Mux_v I__4726 (
            .O(N__22686),
            .I(N__22683));
    Span4Mux_v I__4725 (
            .O(N__22683),
            .I(N__22680));
    Span4Mux_h I__4724 (
            .O(N__22680),
            .I(N__22677));
    Odrv4 I__4723 (
            .O(N__22677),
            .I(\this_sprites_ram.mem_out_bus7_2 ));
    InMux I__4722 (
            .O(N__22674),
            .I(N__22671));
    LocalMux I__4721 (
            .O(N__22671),
            .I(N__22668));
    Span4Mux_v I__4720 (
            .O(N__22668),
            .I(N__22665));
    Sp12to4 I__4719 (
            .O(N__22665),
            .I(N__22662));
    Odrv12 I__4718 (
            .O(N__22662),
            .I(\this_sprites_ram.mem_out_bus3_2 ));
    InMux I__4717 (
            .O(N__22659),
            .I(N__22656));
    LocalMux I__4716 (
            .O(N__22656),
            .I(N__22653));
    Span12Mux_v I__4715 (
            .O(N__22653),
            .I(N__22650));
    Odrv12 I__4714 (
            .O(N__22650),
            .I(\this_sprites_ram.mem_out_bus4_2 ));
    InMux I__4713 (
            .O(N__22647),
            .I(N__22644));
    LocalMux I__4712 (
            .O(N__22644),
            .I(N__22641));
    Span4Mux_v I__4711 (
            .O(N__22641),
            .I(N__22638));
    Span4Mux_h I__4710 (
            .O(N__22638),
            .I(N__22635));
    Odrv4 I__4709 (
            .O(N__22635),
            .I(\this_sprites_ram.mem_out_bus0_2 ));
    CascadeMux I__4708 (
            .O(N__22632),
            .I(N__22629));
    InMux I__4707 (
            .O(N__22629),
            .I(N__22625));
    CascadeMux I__4706 (
            .O(N__22628),
            .I(N__22621));
    LocalMux I__4705 (
            .O(N__22625),
            .I(N__22617));
    InMux I__4704 (
            .O(N__22624),
            .I(N__22614));
    InMux I__4703 (
            .O(N__22621),
            .I(N__22611));
    InMux I__4702 (
            .O(N__22620),
            .I(N__22608));
    Span4Mux_v I__4701 (
            .O(N__22617),
            .I(N__22605));
    LocalMux I__4700 (
            .O(N__22614),
            .I(N__22602));
    LocalMux I__4699 (
            .O(N__22611),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    LocalMux I__4698 (
            .O(N__22608),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv4 I__4697 (
            .O(N__22605),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv4 I__4696 (
            .O(N__22602),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    CascadeMux I__4695 (
            .O(N__22593),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ));
    InMux I__4694 (
            .O(N__22590),
            .I(N__22587));
    LocalMux I__4693 (
            .O(N__22587),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ));
    CascadeMux I__4692 (
            .O(N__22584),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ));
    InMux I__4691 (
            .O(N__22581),
            .I(N__22578));
    LocalMux I__4690 (
            .O(N__22578),
            .I(N__22575));
    Span12Mux_s9_v I__4689 (
            .O(N__22575),
            .I(N__22572));
    Span12Mux_h I__4688 (
            .O(N__22572),
            .I(N__22568));
    InMux I__4687 (
            .O(N__22571),
            .I(N__22565));
    Odrv12 I__4686 (
            .O(N__22568),
            .I(M_this_ppu_vram_data_2));
    LocalMux I__4685 (
            .O(N__22565),
            .I(M_this_ppu_vram_data_2));
    InMux I__4684 (
            .O(N__22560),
            .I(N__22557));
    LocalMux I__4683 (
            .O(N__22557),
            .I(N__22554));
    Span4Mux_v I__4682 (
            .O(N__22554),
            .I(N__22551));
    Span4Mux_v I__4681 (
            .O(N__22551),
            .I(N__22548));
    Sp12to4 I__4680 (
            .O(N__22548),
            .I(N__22545));
    Span12Mux_v I__4679 (
            .O(N__22545),
            .I(N__22542));
    Span12Mux_h I__4678 (
            .O(N__22542),
            .I(N__22539));
    Odrv12 I__4677 (
            .O(N__22539),
            .I(M_this_map_ram_read_data_0));
    CascadeMux I__4676 (
            .O(N__22536),
            .I(N__22532));
    CascadeMux I__4675 (
            .O(N__22535),
            .I(N__22521));
    InMux I__4674 (
            .O(N__22532),
            .I(N__22518));
    CascadeMux I__4673 (
            .O(N__22531),
            .I(N__22515));
    CascadeMux I__4672 (
            .O(N__22530),
            .I(N__22512));
    CascadeMux I__4671 (
            .O(N__22529),
            .I(N__22508));
    CascadeMux I__4670 (
            .O(N__22528),
            .I(N__22503));
    CascadeMux I__4669 (
            .O(N__22527),
            .I(N__22500));
    CascadeMux I__4668 (
            .O(N__22526),
            .I(N__22497));
    CascadeMux I__4667 (
            .O(N__22525),
            .I(N__22494));
    CascadeMux I__4666 (
            .O(N__22524),
            .I(N__22491));
    InMux I__4665 (
            .O(N__22521),
            .I(N__22488));
    LocalMux I__4664 (
            .O(N__22518),
            .I(N__22484));
    InMux I__4663 (
            .O(N__22515),
            .I(N__22481));
    InMux I__4662 (
            .O(N__22512),
            .I(N__22477));
    CascadeMux I__4661 (
            .O(N__22511),
            .I(N__22474));
    InMux I__4660 (
            .O(N__22508),
            .I(N__22471));
    CascadeMux I__4659 (
            .O(N__22507),
            .I(N__22468));
    CascadeMux I__4658 (
            .O(N__22506),
            .I(N__22465));
    InMux I__4657 (
            .O(N__22503),
            .I(N__22461));
    InMux I__4656 (
            .O(N__22500),
            .I(N__22458));
    InMux I__4655 (
            .O(N__22497),
            .I(N__22455));
    InMux I__4654 (
            .O(N__22494),
            .I(N__22452));
    InMux I__4653 (
            .O(N__22491),
            .I(N__22449));
    LocalMux I__4652 (
            .O(N__22488),
            .I(N__22446));
    CascadeMux I__4651 (
            .O(N__22487),
            .I(N__22443));
    Span4Mux_v I__4650 (
            .O(N__22484),
            .I(N__22438));
    LocalMux I__4649 (
            .O(N__22481),
            .I(N__22438));
    CascadeMux I__4648 (
            .O(N__22480),
            .I(N__22435));
    LocalMux I__4647 (
            .O(N__22477),
            .I(N__22432));
    InMux I__4646 (
            .O(N__22474),
            .I(N__22429));
    LocalMux I__4645 (
            .O(N__22471),
            .I(N__22426));
    InMux I__4644 (
            .O(N__22468),
            .I(N__22423));
    InMux I__4643 (
            .O(N__22465),
            .I(N__22420));
    CascadeMux I__4642 (
            .O(N__22464),
            .I(N__22417));
    LocalMux I__4641 (
            .O(N__22461),
            .I(N__22414));
    LocalMux I__4640 (
            .O(N__22458),
            .I(N__22405));
    LocalMux I__4639 (
            .O(N__22455),
            .I(N__22405));
    LocalMux I__4638 (
            .O(N__22452),
            .I(N__22405));
    LocalMux I__4637 (
            .O(N__22449),
            .I(N__22405));
    Span4Mux_s2_v I__4636 (
            .O(N__22446),
            .I(N__22402));
    InMux I__4635 (
            .O(N__22443),
            .I(N__22399));
    Span4Mux_v I__4634 (
            .O(N__22438),
            .I(N__22396));
    InMux I__4633 (
            .O(N__22435),
            .I(N__22393));
    Span4Mux_h I__4632 (
            .O(N__22432),
            .I(N__22390));
    LocalMux I__4631 (
            .O(N__22429),
            .I(N__22387));
    Span4Mux_h I__4630 (
            .O(N__22426),
            .I(N__22384));
    LocalMux I__4629 (
            .O(N__22423),
            .I(N__22381));
    LocalMux I__4628 (
            .O(N__22420),
            .I(N__22378));
    InMux I__4627 (
            .O(N__22417),
            .I(N__22375));
    Span4Mux_h I__4626 (
            .O(N__22414),
            .I(N__22372));
    Span12Mux_v I__4625 (
            .O(N__22405),
            .I(N__22369));
    Sp12to4 I__4624 (
            .O(N__22402),
            .I(N__22364));
    LocalMux I__4623 (
            .O(N__22399),
            .I(N__22364));
    Sp12to4 I__4622 (
            .O(N__22396),
            .I(N__22359));
    LocalMux I__4621 (
            .O(N__22393),
            .I(N__22359));
    Span4Mux_v I__4620 (
            .O(N__22390),
            .I(N__22354));
    Span4Mux_h I__4619 (
            .O(N__22387),
            .I(N__22354));
    Span4Mux_v I__4618 (
            .O(N__22384),
            .I(N__22349));
    Span4Mux_h I__4617 (
            .O(N__22381),
            .I(N__22349));
    Span4Mux_h I__4616 (
            .O(N__22378),
            .I(N__22346));
    LocalMux I__4615 (
            .O(N__22375),
            .I(N__22343));
    Sp12to4 I__4614 (
            .O(N__22372),
            .I(N__22340));
    Span12Mux_h I__4613 (
            .O(N__22369),
            .I(N__22333));
    Span12Mux_h I__4612 (
            .O(N__22364),
            .I(N__22333));
    Span12Mux_h I__4611 (
            .O(N__22359),
            .I(N__22333));
    Span4Mux_h I__4610 (
            .O(N__22354),
            .I(N__22328));
    Span4Mux_h I__4609 (
            .O(N__22349),
            .I(N__22328));
    Span4Mux_v I__4608 (
            .O(N__22346),
            .I(N__22323));
    Span4Mux_h I__4607 (
            .O(N__22343),
            .I(N__22323));
    Odrv12 I__4606 (
            .O(N__22340),
            .I(M_this_ppu_sprites_addr_6));
    Odrv12 I__4605 (
            .O(N__22333),
            .I(M_this_ppu_sprites_addr_6));
    Odrv4 I__4604 (
            .O(N__22328),
            .I(M_this_ppu_sprites_addr_6));
    Odrv4 I__4603 (
            .O(N__22323),
            .I(M_this_ppu_sprites_addr_6));
    InMux I__4602 (
            .O(N__22314),
            .I(N__22311));
    LocalMux I__4601 (
            .O(N__22311),
            .I(N__22308));
    Span4Mux_v I__4600 (
            .O(N__22308),
            .I(N__22305));
    Span4Mux_h I__4599 (
            .O(N__22305),
            .I(N__22302));
    Odrv4 I__4598 (
            .O(N__22302),
            .I(\this_sprites_ram.mem_out_bus6_2 ));
    InMux I__4597 (
            .O(N__22299),
            .I(N__22296));
    LocalMux I__4596 (
            .O(N__22296),
            .I(N__22293));
    Span12Mux_v I__4595 (
            .O(N__22293),
            .I(N__22290));
    Odrv12 I__4594 (
            .O(N__22290),
            .I(\this_sprites_ram.mem_out_bus2_2 ));
    InMux I__4593 (
            .O(N__22287),
            .I(N__22284));
    LocalMux I__4592 (
            .O(N__22284),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ));
    InMux I__4591 (
            .O(N__22281),
            .I(N__22277));
    InMux I__4590 (
            .O(N__22280),
            .I(N__22274));
    LocalMux I__4589 (
            .O(N__22277),
            .I(\this_ppu.M_this_ppu_map_addr_i_3 ));
    LocalMux I__4588 (
            .O(N__22274),
            .I(\this_ppu.M_this_ppu_map_addr_i_3 ));
    CascadeMux I__4587 (
            .O(N__22269),
            .I(N__22266));
    InMux I__4586 (
            .O(N__22266),
            .I(N__22262));
    InMux I__4585 (
            .O(N__22265),
            .I(N__22259));
    LocalMux I__4584 (
            .O(N__22262),
            .I(\this_ppu.M_this_ppu_map_addr_i_4 ));
    LocalMux I__4583 (
            .O(N__22259),
            .I(\this_ppu.M_this_ppu_map_addr_i_4 ));
    InMux I__4582 (
            .O(N__22254),
            .I(bfn_19_20_0_));
    InMux I__4581 (
            .O(N__22251),
            .I(N__22248));
    LocalMux I__4580 (
            .O(N__22248),
            .I(\this_ppu.vscroll8_1 ));
    CascadeMux I__4579 (
            .O(N__22245),
            .I(N__22242));
    InMux I__4578 (
            .O(N__22242),
            .I(N__22239));
    LocalMux I__4577 (
            .O(N__22239),
            .I(N__22236));
    Span4Mux_v I__4576 (
            .O(N__22236),
            .I(N__22233));
    Span4Mux_v I__4575 (
            .O(N__22233),
            .I(N__22230));
    Odrv4 I__4574 (
            .O(N__22230),
            .I(\this_ppu.un1_M_vaddress_q_3_4 ));
    InMux I__4573 (
            .O(N__22227),
            .I(N__22224));
    LocalMux I__4572 (
            .O(N__22224),
            .I(N__22221));
    Span12Mux_v I__4571 (
            .O(N__22221),
            .I(N__22218));
    Span12Mux_h I__4570 (
            .O(N__22218),
            .I(N__22215));
    Odrv12 I__4569 (
            .O(N__22215),
            .I(\this_sprites_ram.mem_out_bus4_1 ));
    InMux I__4568 (
            .O(N__22212),
            .I(N__22209));
    LocalMux I__4567 (
            .O(N__22209),
            .I(N__22206));
    Span4Mux_v I__4566 (
            .O(N__22206),
            .I(N__22203));
    Span4Mux_h I__4565 (
            .O(N__22203),
            .I(N__22200));
    Span4Mux_v I__4564 (
            .O(N__22200),
            .I(N__22197));
    Odrv4 I__4563 (
            .O(N__22197),
            .I(\this_sprites_ram.mem_out_bus0_1 ));
    InMux I__4562 (
            .O(N__22194),
            .I(N__22191));
    LocalMux I__4561 (
            .O(N__22191),
            .I(N__22188));
    Span4Mux_v I__4560 (
            .O(N__22188),
            .I(N__22185));
    Span4Mux_v I__4559 (
            .O(N__22185),
            .I(N__22182));
    Span4Mux_h I__4558 (
            .O(N__22182),
            .I(N__22179));
    Odrv4 I__4557 (
            .O(N__22179),
            .I(\this_sprites_ram.mem_out_bus7_1 ));
    InMux I__4556 (
            .O(N__22176),
            .I(N__22173));
    LocalMux I__4555 (
            .O(N__22173),
            .I(N__22170));
    Sp12to4 I__4554 (
            .O(N__22170),
            .I(N__22167));
    Odrv12 I__4553 (
            .O(N__22167),
            .I(\this_sprites_ram.mem_out_bus3_1 ));
    CascadeMux I__4552 (
            .O(N__22164),
            .I(N__22161));
    InMux I__4551 (
            .O(N__22161),
            .I(N__22158));
    LocalMux I__4550 (
            .O(N__22158),
            .I(N__22155));
    Span12Mux_v I__4549 (
            .O(N__22155),
            .I(N__22152));
    Span12Mux_h I__4548 (
            .O(N__22152),
            .I(N__22149));
    Odrv12 I__4547 (
            .O(N__22149),
            .I(M_this_map_ram_read_data_6));
    InMux I__4546 (
            .O(N__22146),
            .I(N__22143));
    LocalMux I__4545 (
            .O(N__22143),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ));
    CascadeMux I__4544 (
            .O(N__22140),
            .I(N__22137));
    CascadeBuf I__4543 (
            .O(N__22137),
            .I(N__22134));
    CascadeMux I__4542 (
            .O(N__22134),
            .I(N__22131));
    InMux I__4541 (
            .O(N__22131),
            .I(N__22128));
    LocalMux I__4540 (
            .O(N__22128),
            .I(N__22125));
    Sp12to4 I__4539 (
            .O(N__22125),
            .I(N__22120));
    InMux I__4538 (
            .O(N__22124),
            .I(N__22117));
    InMux I__4537 (
            .O(N__22123),
            .I(N__22114));
    Span12Mux_v I__4536 (
            .O(N__22120),
            .I(N__22111));
    LocalMux I__4535 (
            .O(N__22117),
            .I(M_this_ppu_map_addr_9));
    LocalMux I__4534 (
            .O(N__22114),
            .I(M_this_ppu_map_addr_9));
    Odrv12 I__4533 (
            .O(N__22111),
            .I(M_this_ppu_map_addr_9));
    InMux I__4532 (
            .O(N__22104),
            .I(bfn_19_18_0_));
    InMux I__4531 (
            .O(N__22101),
            .I(N__22098));
    LocalMux I__4530 (
            .O(N__22098),
            .I(N__22095));
    Odrv4 I__4529 (
            .O(N__22095),
            .I(\this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO ));
    InMux I__4528 (
            .O(N__22092),
            .I(N__22089));
    LocalMux I__4527 (
            .O(N__22089),
            .I(N__22086));
    Span4Mux_h I__4526 (
            .O(N__22086),
            .I(N__22083));
    Odrv4 I__4525 (
            .O(N__22083),
            .I(\this_reset_cond.M_stage_qZ0Z_3 ));
    InMux I__4524 (
            .O(N__22080),
            .I(N__22076));
    InMux I__4523 (
            .O(N__22079),
            .I(N__22073));
    LocalMux I__4522 (
            .O(N__22076),
            .I(\this_ppu.M_this_ppu_vram_addr_i_0 ));
    LocalMux I__4521 (
            .O(N__22073),
            .I(\this_ppu.M_this_ppu_vram_addr_i_0 ));
    InMux I__4520 (
            .O(N__22068),
            .I(N__22064));
    InMux I__4519 (
            .O(N__22067),
            .I(N__22061));
    LocalMux I__4518 (
            .O(N__22064),
            .I(\this_ppu.M_this_ppu_vram_addr_i_1 ));
    LocalMux I__4517 (
            .O(N__22061),
            .I(\this_ppu.M_this_ppu_vram_addr_i_1 ));
    CascadeMux I__4516 (
            .O(N__22056),
            .I(N__22053));
    InMux I__4515 (
            .O(N__22053),
            .I(N__22050));
    LocalMux I__4514 (
            .O(N__22050),
            .I(N__22046));
    InMux I__4513 (
            .O(N__22049),
            .I(N__22043));
    Odrv4 I__4512 (
            .O(N__22046),
            .I(\this_ppu.M_this_ppu_vram_addr_i_2 ));
    LocalMux I__4511 (
            .O(N__22043),
            .I(\this_ppu.M_this_ppu_vram_addr_i_2 ));
    CascadeMux I__4510 (
            .O(N__22038),
            .I(N__22034));
    InMux I__4509 (
            .O(N__22037),
            .I(N__22031));
    InMux I__4508 (
            .O(N__22034),
            .I(N__22028));
    LocalMux I__4507 (
            .O(N__22031),
            .I(\this_ppu.M_this_ppu_map_addr_i_0 ));
    LocalMux I__4506 (
            .O(N__22028),
            .I(\this_ppu.M_this_ppu_map_addr_i_0 ));
    CascadeMux I__4505 (
            .O(N__22023),
            .I(N__22019));
    InMux I__4504 (
            .O(N__22022),
            .I(N__22016));
    InMux I__4503 (
            .O(N__22019),
            .I(N__22013));
    LocalMux I__4502 (
            .O(N__22016),
            .I(\this_ppu.M_this_ppu_map_addr_i_1 ));
    LocalMux I__4501 (
            .O(N__22013),
            .I(\this_ppu.M_this_ppu_map_addr_i_1 ));
    CascadeMux I__4500 (
            .O(N__22008),
            .I(N__22004));
    InMux I__4499 (
            .O(N__22007),
            .I(N__22001));
    InMux I__4498 (
            .O(N__22004),
            .I(N__21998));
    LocalMux I__4497 (
            .O(N__22001),
            .I(\this_ppu.M_this_ppu_map_addr_i_2 ));
    LocalMux I__4496 (
            .O(N__21998),
            .I(\this_ppu.M_this_ppu_map_addr_i_2 ));
    InMux I__4495 (
            .O(N__21993),
            .I(N__21987));
    InMux I__4494 (
            .O(N__21992),
            .I(N__21987));
    LocalMux I__4493 (
            .O(N__21987),
            .I(N__21984));
    Odrv4 I__4492 (
            .O(N__21984),
            .I(\this_ppu.un1_M_vaddress_q_2_c2 ));
    SRMux I__4491 (
            .O(N__21981),
            .I(N__21978));
    LocalMux I__4490 (
            .O(N__21978),
            .I(N__21975));
    Span4Mux_v I__4489 (
            .O(N__21975),
            .I(N__21971));
    SRMux I__4488 (
            .O(N__21974),
            .I(N__21968));
    Span4Mux_h I__4487 (
            .O(N__21971),
            .I(N__21963));
    LocalMux I__4486 (
            .O(N__21968),
            .I(N__21963));
    Span4Mux_h I__4485 (
            .O(N__21963),
            .I(N__21960));
    Odrv4 I__4484 (
            .O(N__21960),
            .I(\this_ppu.M_state_q_RNILG0GDZ0Z_0 ));
    CascadeMux I__4483 (
            .O(N__21957),
            .I(N__21954));
    CascadeBuf I__4482 (
            .O(N__21954),
            .I(N__21951));
    CascadeMux I__4481 (
            .O(N__21951),
            .I(N__21948));
    InMux I__4480 (
            .O(N__21948),
            .I(N__21945));
    LocalMux I__4479 (
            .O(N__21945),
            .I(N__21942));
    Sp12to4 I__4478 (
            .O(N__21942),
            .I(N__21938));
    CascadeMux I__4477 (
            .O(N__21941),
            .I(N__21935));
    Span12Mux_s4_v I__4476 (
            .O(N__21938),
            .I(N__21929));
    InMux I__4475 (
            .O(N__21935),
            .I(N__21924));
    InMux I__4474 (
            .O(N__21934),
            .I(N__21924));
    InMux I__4473 (
            .O(N__21933),
            .I(N__21921));
    InMux I__4472 (
            .O(N__21932),
            .I(N__21918));
    Span12Mux_v I__4471 (
            .O(N__21929),
            .I(N__21915));
    LocalMux I__4470 (
            .O(N__21924),
            .I(M_this_ppu_map_addr_5));
    LocalMux I__4469 (
            .O(N__21921),
            .I(M_this_ppu_map_addr_5));
    LocalMux I__4468 (
            .O(N__21918),
            .I(M_this_ppu_map_addr_5));
    Odrv12 I__4467 (
            .O(N__21915),
            .I(M_this_ppu_map_addr_5));
    CascadeMux I__4466 (
            .O(N__21906),
            .I(N__21903));
    CascadeBuf I__4465 (
            .O(N__21903),
            .I(N__21900));
    CascadeMux I__4464 (
            .O(N__21900),
            .I(N__21897));
    InMux I__4463 (
            .O(N__21897),
            .I(N__21894));
    LocalMux I__4462 (
            .O(N__21894),
            .I(N__21888));
    InMux I__4461 (
            .O(N__21893),
            .I(N__21885));
    InMux I__4460 (
            .O(N__21892),
            .I(N__21882));
    InMux I__4459 (
            .O(N__21891),
            .I(N__21879));
    Span12Mux_v I__4458 (
            .O(N__21888),
            .I(N__21876));
    LocalMux I__4457 (
            .O(N__21885),
            .I(M_this_ppu_map_addr_6));
    LocalMux I__4456 (
            .O(N__21882),
            .I(M_this_ppu_map_addr_6));
    LocalMux I__4455 (
            .O(N__21879),
            .I(M_this_ppu_map_addr_6));
    Odrv12 I__4454 (
            .O(N__21876),
            .I(M_this_ppu_map_addr_6));
    CascadeMux I__4453 (
            .O(N__21867),
            .I(N__21864));
    CascadeBuf I__4452 (
            .O(N__21864),
            .I(N__21861));
    CascadeMux I__4451 (
            .O(N__21861),
            .I(N__21858));
    InMux I__4450 (
            .O(N__21858),
            .I(N__21855));
    LocalMux I__4449 (
            .O(N__21855),
            .I(N__21852));
    Span4Mux_v I__4448 (
            .O(N__21852),
            .I(N__21849));
    Span4Mux_v I__4447 (
            .O(N__21849),
            .I(N__21846));
    Span4Mux_v I__4446 (
            .O(N__21846),
            .I(N__21839));
    InMux I__4445 (
            .O(N__21845),
            .I(N__21832));
    InMux I__4444 (
            .O(N__21844),
            .I(N__21832));
    InMux I__4443 (
            .O(N__21843),
            .I(N__21832));
    InMux I__4442 (
            .O(N__21842),
            .I(N__21829));
    Sp12to4 I__4441 (
            .O(N__21839),
            .I(N__21826));
    LocalMux I__4440 (
            .O(N__21832),
            .I(M_this_ppu_map_addr_7));
    LocalMux I__4439 (
            .O(N__21829),
            .I(M_this_ppu_map_addr_7));
    Odrv12 I__4438 (
            .O(N__21826),
            .I(M_this_ppu_map_addr_7));
    CascadeMux I__4437 (
            .O(N__21819),
            .I(N__21816));
    CascadeBuf I__4436 (
            .O(N__21816),
            .I(N__21813));
    CascadeMux I__4435 (
            .O(N__21813),
            .I(N__21810));
    InMux I__4434 (
            .O(N__21810),
            .I(N__21806));
    CascadeMux I__4433 (
            .O(N__21809),
            .I(N__21803));
    LocalMux I__4432 (
            .O(N__21806),
            .I(N__21798));
    InMux I__4431 (
            .O(N__21803),
            .I(N__21793));
    InMux I__4430 (
            .O(N__21802),
            .I(N__21793));
    InMux I__4429 (
            .O(N__21801),
            .I(N__21790));
    Span12Mux_v I__4428 (
            .O(N__21798),
            .I(N__21787));
    LocalMux I__4427 (
            .O(N__21793),
            .I(M_this_ppu_map_addr_8));
    LocalMux I__4426 (
            .O(N__21790),
            .I(M_this_ppu_map_addr_8));
    Odrv12 I__4425 (
            .O(N__21787),
            .I(M_this_ppu_map_addr_8));
    CascadeMux I__4424 (
            .O(N__21780),
            .I(\this_vga_signals.M_this_state_q_srsts_i_a3_0_7_cascade_ ));
    CascadeMux I__4423 (
            .O(N__21777),
            .I(\this_vga_signals.M_this_state_q_srsts_i_0Z0Z_7_cascade_ ));
    InMux I__4422 (
            .O(N__21774),
            .I(N__21771));
    LocalMux I__4421 (
            .O(N__21771),
            .I(N__21768));
    Odrv4 I__4420 (
            .O(N__21768),
            .I(M_this_state_q_RNI6Q0SZ0Z_5));
    CascadeMux I__4419 (
            .O(N__21765),
            .I(N__21762));
    InMux I__4418 (
            .O(N__21762),
            .I(N__21759));
    LocalMux I__4417 (
            .O(N__21759),
            .I(N__21753));
    InMux I__4416 (
            .O(N__21758),
            .I(N__21750));
    InMux I__4415 (
            .O(N__21757),
            .I(N__21747));
    InMux I__4414 (
            .O(N__21756),
            .I(N__21744));
    Span4Mux_v I__4413 (
            .O(N__21753),
            .I(N__21741));
    LocalMux I__4412 (
            .O(N__21750),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__4411 (
            .O(N__21747),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__4410 (
            .O(N__21744),
            .I(M_this_state_qZ0Z_12));
    Odrv4 I__4409 (
            .O(N__21741),
            .I(M_this_state_qZ0Z_12));
    InMux I__4408 (
            .O(N__21732),
            .I(N__21723));
    InMux I__4407 (
            .O(N__21731),
            .I(N__21723));
    InMux I__4406 (
            .O(N__21730),
            .I(N__21717));
    InMux I__4405 (
            .O(N__21729),
            .I(N__21714));
    InMux I__4404 (
            .O(N__21728),
            .I(N__21711));
    LocalMux I__4403 (
            .O(N__21723),
            .I(N__21708));
    InMux I__4402 (
            .O(N__21722),
            .I(N__21703));
    InMux I__4401 (
            .O(N__21721),
            .I(N__21703));
    InMux I__4400 (
            .O(N__21720),
            .I(N__21700));
    LocalMux I__4399 (
            .O(N__21717),
            .I(N_848));
    LocalMux I__4398 (
            .O(N__21714),
            .I(N_848));
    LocalMux I__4397 (
            .O(N__21711),
            .I(N_848));
    Odrv4 I__4396 (
            .O(N__21708),
            .I(N_848));
    LocalMux I__4395 (
            .O(N__21703),
            .I(N_848));
    LocalMux I__4394 (
            .O(N__21700),
            .I(N_848));
    InMux I__4393 (
            .O(N__21687),
            .I(N__21681));
    InMux I__4392 (
            .O(N__21686),
            .I(N__21681));
    LocalMux I__4391 (
            .O(N__21681),
            .I(\this_vga_signals.N_93_0 ));
    InMux I__4390 (
            .O(N__21678),
            .I(N__21675));
    LocalMux I__4389 (
            .O(N__21675),
            .I(N__21670));
    InMux I__4388 (
            .O(N__21674),
            .I(N__21667));
    CascadeMux I__4387 (
            .O(N__21673),
            .I(N__21664));
    Span4Mux_v I__4386 (
            .O(N__21670),
            .I(N__21658));
    LocalMux I__4385 (
            .O(N__21667),
            .I(N__21655));
    InMux I__4384 (
            .O(N__21664),
            .I(N__21648));
    InMux I__4383 (
            .O(N__21663),
            .I(N__21648));
    InMux I__4382 (
            .O(N__21662),
            .I(N__21648));
    InMux I__4381 (
            .O(N__21661),
            .I(N__21645));
    Odrv4 I__4380 (
            .O(N__21658),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv4 I__4379 (
            .O(N__21655),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__4378 (
            .O(N__21648),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__4377 (
            .O(N__21645),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    InMux I__4376 (
            .O(N__21636),
            .I(N__21633));
    LocalMux I__4375 (
            .O(N__21633),
            .I(N__21630));
    Span4Mux_v I__4374 (
            .O(N__21630),
            .I(N__21624));
    InMux I__4373 (
            .O(N__21629),
            .I(N__21617));
    InMux I__4372 (
            .O(N__21628),
            .I(N__21617));
    InMux I__4371 (
            .O(N__21627),
            .I(N__21617));
    Span4Mux_h I__4370 (
            .O(N__21624),
            .I(N__21611));
    LocalMux I__4369 (
            .O(N__21617),
            .I(N__21611));
    InMux I__4368 (
            .O(N__21616),
            .I(N__21608));
    Odrv4 I__4367 (
            .O(N__21611),
            .I(M_this_vga_signals_line_clk_0));
    LocalMux I__4366 (
            .O(N__21608),
            .I(M_this_vga_signals_line_clk_0));
    CascadeMux I__4365 (
            .O(N__21603),
            .I(N__21599));
    CascadeMux I__4364 (
            .O(N__21602),
            .I(N__21596));
    InMux I__4363 (
            .O(N__21599),
            .I(N__21593));
    InMux I__4362 (
            .O(N__21596),
            .I(N__21588));
    LocalMux I__4361 (
            .O(N__21593),
            .I(N__21585));
    InMux I__4360 (
            .O(N__21592),
            .I(N__21580));
    InMux I__4359 (
            .O(N__21591),
            .I(N__21580));
    LocalMux I__4358 (
            .O(N__21588),
            .I(N__21577));
    Span12Mux_v I__4357 (
            .O(N__21585),
            .I(N__21572));
    LocalMux I__4356 (
            .O(N__21580),
            .I(N__21567));
    Span4Mux_h I__4355 (
            .O(N__21577),
            .I(N__21567));
    InMux I__4354 (
            .O(N__21576),
            .I(N__21564));
    InMux I__4353 (
            .O(N__21575),
            .I(N__21561));
    Odrv12 I__4352 (
            .O(N__21572),
            .I(\this_ppu.M_last_q ));
    Odrv4 I__4351 (
            .O(N__21567),
            .I(\this_ppu.M_last_q ));
    LocalMux I__4350 (
            .O(N__21564),
            .I(\this_ppu.M_last_q ));
    LocalMux I__4349 (
            .O(N__21561),
            .I(\this_ppu.M_last_q ));
    InMux I__4348 (
            .O(N__21552),
            .I(N__21543));
    InMux I__4347 (
            .O(N__21551),
            .I(N__21543));
    InMux I__4346 (
            .O(N__21550),
            .I(N__21538));
    InMux I__4345 (
            .O(N__21549),
            .I(N__21538));
    InMux I__4344 (
            .O(N__21548),
            .I(N__21535));
    LocalMux I__4343 (
            .O(N__21543),
            .I(N__21528));
    LocalMux I__4342 (
            .O(N__21538),
            .I(N__21528));
    LocalMux I__4341 (
            .O(N__21535),
            .I(N__21524));
    InMux I__4340 (
            .O(N__21534),
            .I(N__21521));
    InMux I__4339 (
            .O(N__21533),
            .I(N__21518));
    Span4Mux_v I__4338 (
            .O(N__21528),
            .I(N__21515));
    InMux I__4337 (
            .O(N__21527),
            .I(N__21512));
    Span4Mux_v I__4336 (
            .O(N__21524),
            .I(N__21509));
    LocalMux I__4335 (
            .O(N__21521),
            .I(N__21502));
    LocalMux I__4334 (
            .O(N__21518),
            .I(N__21502));
    Span4Mux_h I__4333 (
            .O(N__21515),
            .I(N__21502));
    LocalMux I__4332 (
            .O(N__21512),
            .I(\this_ppu.N_132_0 ));
    Odrv4 I__4331 (
            .O(N__21509),
            .I(\this_ppu.N_132_0 ));
    Odrv4 I__4330 (
            .O(N__21502),
            .I(\this_ppu.N_132_0 ));
    CascadeMux I__4329 (
            .O(N__21495),
            .I(M_this_state_q_RNIH92SZ0Z_10_cascade_));
    InMux I__4328 (
            .O(N__21492),
            .I(N__21488));
    CascadeMux I__4327 (
            .O(N__21491),
            .I(N__21485));
    LocalMux I__4326 (
            .O(N__21488),
            .I(N__21480));
    InMux I__4325 (
            .O(N__21485),
            .I(N__21477));
    InMux I__4324 (
            .O(N__21484),
            .I(N__21471));
    InMux I__4323 (
            .O(N__21483),
            .I(N__21471));
    Span4Mux_v I__4322 (
            .O(N__21480),
            .I(N__21464));
    LocalMux I__4321 (
            .O(N__21477),
            .I(N__21464));
    InMux I__4320 (
            .O(N__21476),
            .I(N__21461));
    LocalMux I__4319 (
            .O(N__21471),
            .I(N__21458));
    InMux I__4318 (
            .O(N__21470),
            .I(N__21453));
    InMux I__4317 (
            .O(N__21469),
            .I(N__21453));
    Odrv4 I__4316 (
            .O(N__21464),
            .I(\this_vga_signals.N_83 ));
    LocalMux I__4315 (
            .O(N__21461),
            .I(\this_vga_signals.N_83 ));
    Odrv12 I__4314 (
            .O(N__21458),
            .I(\this_vga_signals.N_83 ));
    LocalMux I__4313 (
            .O(N__21453),
            .I(\this_vga_signals.N_83 ));
    CascadeMux I__4312 (
            .O(N__21444),
            .I(N__21441));
    InMux I__4311 (
            .O(N__21441),
            .I(N__21438));
    LocalMux I__4310 (
            .O(N__21438),
            .I(N__21435));
    Span4Mux_h I__4309 (
            .O(N__21435),
            .I(N__21432));
    Odrv4 I__4308 (
            .O(N__21432),
            .I(\this_vga_signals.N_94_0 ));
    CascadeMux I__4307 (
            .O(N__21429),
            .I(\this_vga_signals.N_94_0_cascade_ ));
    InMux I__4306 (
            .O(N__21426),
            .I(N__21423));
    LocalMux I__4305 (
            .O(N__21423),
            .I(\this_vga_signals.M_this_state_q_srsts_i_i_0Z0Z_12 ));
    InMux I__4304 (
            .O(N__21420),
            .I(N__21417));
    LocalMux I__4303 (
            .O(N__21417),
            .I(N__21414));
    Odrv4 I__4302 (
            .O(N__21414),
            .I(M_this_state_q_RNI373A1Z0Z_8));
    CascadeMux I__4301 (
            .O(N__21411),
            .I(this_vga_signals_un21_i_a3_1_1_cascade_));
    InMux I__4300 (
            .O(N__21408),
            .I(N__21405));
    LocalMux I__4299 (
            .O(N__21405),
            .I(N__21401));
    InMux I__4298 (
            .O(N__21404),
            .I(N__21397));
    Span4Mux_h I__4297 (
            .O(N__21401),
            .I(N__21394));
    IoInMux I__4296 (
            .O(N__21400),
            .I(N__21391));
    LocalMux I__4295 (
            .O(N__21397),
            .I(N__21388));
    Span4Mux_v I__4294 (
            .O(N__21394),
            .I(N__21385));
    LocalMux I__4293 (
            .O(N__21391),
            .I(N__21381));
    Sp12to4 I__4292 (
            .O(N__21388),
            .I(N__21378));
    Span4Mux_h I__4291 (
            .O(N__21385),
            .I(N__21375));
    InMux I__4290 (
            .O(N__21384),
            .I(N__21372));
    Span12Mux_s6_h I__4289 (
            .O(N__21381),
            .I(N__21368));
    Span12Mux_v I__4288 (
            .O(N__21378),
            .I(N__21365));
    Span4Mux_h I__4287 (
            .O(N__21375),
            .I(N__21362));
    LocalMux I__4286 (
            .O(N__21372),
            .I(N__21359));
    InMux I__4285 (
            .O(N__21371),
            .I(N__21356));
    Span12Mux_h I__4284 (
            .O(N__21368),
            .I(N__21353));
    Span12Mux_h I__4283 (
            .O(N__21365),
            .I(N__21350));
    Span4Mux_h I__4282 (
            .O(N__21362),
            .I(N__21345));
    Span4Mux_v I__4281 (
            .O(N__21359),
            .I(N__21345));
    LocalMux I__4280 (
            .O(N__21356),
            .I(N__21342));
    Odrv12 I__4279 (
            .O(N__21353),
            .I(port_dmab_c));
    Odrv12 I__4278 (
            .O(N__21350),
            .I(port_dmab_c));
    Odrv4 I__4277 (
            .O(N__21345),
            .I(port_dmab_c));
    Odrv4 I__4276 (
            .O(N__21342),
            .I(port_dmab_c));
    InMux I__4275 (
            .O(N__21333),
            .I(N__21329));
    InMux I__4274 (
            .O(N__21332),
            .I(N__21325));
    LocalMux I__4273 (
            .O(N__21329),
            .I(N__21322));
    InMux I__4272 (
            .O(N__21328),
            .I(N__21319));
    LocalMux I__4271 (
            .O(N__21325),
            .I(M_this_data_count_qZ0Z_8));
    Odrv4 I__4270 (
            .O(N__21322),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__4269 (
            .O(N__21319),
            .I(M_this_data_count_qZ0Z_8));
    CascadeMux I__4268 (
            .O(N__21312),
            .I(N__21309));
    InMux I__4267 (
            .O(N__21309),
            .I(N__21305));
    InMux I__4266 (
            .O(N__21308),
            .I(N__21302));
    LocalMux I__4265 (
            .O(N__21305),
            .I(N__21296));
    LocalMux I__4264 (
            .O(N__21302),
            .I(N__21296));
    InMux I__4263 (
            .O(N__21301),
            .I(N__21293));
    Span4Mux_h I__4262 (
            .O(N__21296),
            .I(N__21290));
    LocalMux I__4261 (
            .O(N__21293),
            .I(M_this_data_count_qZ0Z_5));
    Odrv4 I__4260 (
            .O(N__21290),
            .I(M_this_data_count_qZ0Z_5));
    CascadeMux I__4259 (
            .O(N__21285),
            .I(N__21282));
    InMux I__4258 (
            .O(N__21282),
            .I(N__21277));
    CascadeMux I__4257 (
            .O(N__21281),
            .I(N__21274));
    InMux I__4256 (
            .O(N__21280),
            .I(N__21271));
    LocalMux I__4255 (
            .O(N__21277),
            .I(N__21268));
    InMux I__4254 (
            .O(N__21274),
            .I(N__21265));
    LocalMux I__4253 (
            .O(N__21271),
            .I(M_this_data_count_qZ0Z_9));
    Odrv4 I__4252 (
            .O(N__21268),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__4251 (
            .O(N__21265),
            .I(M_this_data_count_qZ0Z_9));
    InMux I__4250 (
            .O(N__21258),
            .I(N__21253));
    InMux I__4249 (
            .O(N__21257),
            .I(N__21250));
    InMux I__4248 (
            .O(N__21256),
            .I(N__21247));
    LocalMux I__4247 (
            .O(N__21253),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__4246 (
            .O(N__21250),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__4245 (
            .O(N__21247),
            .I(M_this_data_count_qZ0Z_4));
    InMux I__4244 (
            .O(N__21240),
            .I(N__21237));
    LocalMux I__4243 (
            .O(N__21237),
            .I(N__21234));
    Odrv4 I__4242 (
            .O(N__21234),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_8 ));
    CascadeMux I__4241 (
            .O(N__21231),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_ ));
    InMux I__4240 (
            .O(N__21228),
            .I(N__21225));
    LocalMux I__4239 (
            .O(N__21225),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ));
    CascadeMux I__4238 (
            .O(N__21222),
            .I(N__21219));
    InMux I__4237 (
            .O(N__21219),
            .I(N__21216));
    LocalMux I__4236 (
            .O(N__21216),
            .I(N__21213));
    Span4Mux_v I__4235 (
            .O(N__21213),
            .I(N__21210));
    Sp12to4 I__4234 (
            .O(N__21210),
            .I(N__21207));
    Span12Mux_v I__4233 (
            .O(N__21207),
            .I(N__21204));
    Span12Mux_h I__4232 (
            .O(N__21204),
            .I(N__21201));
    Odrv12 I__4231 (
            .O(N__21201),
            .I(M_this_map_ram_read_data_7));
    InMux I__4230 (
            .O(N__21198),
            .I(N__21195));
    LocalMux I__4229 (
            .O(N__21195),
            .I(N__21192));
    Span4Mux_h I__4228 (
            .O(N__21192),
            .I(N__21189));
    Span4Mux_v I__4227 (
            .O(N__21189),
            .I(N__21186));
    Span4Mux_v I__4226 (
            .O(N__21186),
            .I(N__21183));
    Span4Mux_h I__4225 (
            .O(N__21183),
            .I(N__21180));
    Odrv4 I__4224 (
            .O(N__21180),
            .I(\this_sprites_ram.mem_out_bus7_3 ));
    InMux I__4223 (
            .O(N__21177),
            .I(N__21174));
    LocalMux I__4222 (
            .O(N__21174),
            .I(N__21171));
    Span4Mux_v I__4221 (
            .O(N__21171),
            .I(N__21168));
    Span4Mux_h I__4220 (
            .O(N__21168),
            .I(N__21165));
    Span4Mux_h I__4219 (
            .O(N__21165),
            .I(N__21162));
    Odrv4 I__4218 (
            .O(N__21162),
            .I(\this_sprites_ram.mem_out_bus3_3 ));
    InMux I__4217 (
            .O(N__21159),
            .I(N__21156));
    LocalMux I__4216 (
            .O(N__21156),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ));
    InMux I__4215 (
            .O(N__21153),
            .I(N__21150));
    LocalMux I__4214 (
            .O(N__21150),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ));
    InMux I__4213 (
            .O(N__21147),
            .I(N__21144));
    LocalMux I__4212 (
            .O(N__21144),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ));
    CascadeMux I__4211 (
            .O(N__21141),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ));
    InMux I__4210 (
            .O(N__21138),
            .I(N__21135));
    LocalMux I__4209 (
            .O(N__21135),
            .I(N__21132));
    Span4Mux_v I__4208 (
            .O(N__21132),
            .I(N__21129));
    Sp12to4 I__4207 (
            .O(N__21129),
            .I(N__21126));
    Span12Mux_h I__4206 (
            .O(N__21126),
            .I(N__21122));
    InMux I__4205 (
            .O(N__21125),
            .I(N__21119));
    Odrv12 I__4204 (
            .O(N__21122),
            .I(M_this_ppu_vram_data_3));
    LocalMux I__4203 (
            .O(N__21119),
            .I(M_this_ppu_vram_data_3));
    InMux I__4202 (
            .O(N__21114),
            .I(N__21111));
    LocalMux I__4201 (
            .O(N__21111),
            .I(N__21106));
    InMux I__4200 (
            .O(N__21110),
            .I(N__21103));
    InMux I__4199 (
            .O(N__21109),
            .I(N__21100));
    Odrv12 I__4198 (
            .O(N__21106),
            .I(\this_ppu.N_156 ));
    LocalMux I__4197 (
            .O(N__21103),
            .I(\this_ppu.N_156 ));
    LocalMux I__4196 (
            .O(N__21100),
            .I(\this_ppu.N_156 ));
    InMux I__4195 (
            .O(N__21093),
            .I(N__21090));
    LocalMux I__4194 (
            .O(N__21090),
            .I(\this_ppu.N_150 ));
    CascadeMux I__4193 (
            .O(N__21087),
            .I(N__21083));
    CascadeMux I__4192 (
            .O(N__21086),
            .I(N__21080));
    InMux I__4191 (
            .O(N__21083),
            .I(N__21074));
    InMux I__4190 (
            .O(N__21080),
            .I(N__21069));
    InMux I__4189 (
            .O(N__21079),
            .I(N__21069));
    InMux I__4188 (
            .O(N__21078),
            .I(N__21066));
    InMux I__4187 (
            .O(N__21077),
            .I(N__21063));
    LocalMux I__4186 (
            .O(N__21074),
            .I(N__21060));
    LocalMux I__4185 (
            .O(N__21069),
            .I(N__21057));
    LocalMux I__4184 (
            .O(N__21066),
            .I(N__21054));
    LocalMux I__4183 (
            .O(N__21063),
            .I(N__21051));
    Span4Mux_h I__4182 (
            .O(N__21060),
            .I(N__21048));
    Span4Mux_v I__4181 (
            .O(N__21057),
            .I(N__21045));
    Span4Mux_h I__4180 (
            .O(N__21054),
            .I(N__21040));
    Span4Mux_h I__4179 (
            .O(N__21051),
            .I(N__21040));
    Span4Mux_v I__4178 (
            .O(N__21048),
            .I(N__21037));
    Span4Mux_v I__4177 (
            .O(N__21045),
            .I(N__21034));
    Span4Mux_v I__4176 (
            .O(N__21040),
            .I(N__21031));
    Odrv4 I__4175 (
            .O(N__21037),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    Odrv4 I__4174 (
            .O(N__21034),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    Odrv4 I__4173 (
            .O(N__21031),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    CascadeMux I__4172 (
            .O(N__21024),
            .I(N__21021));
    InMux I__4171 (
            .O(N__21021),
            .I(N__21017));
    CascadeMux I__4170 (
            .O(N__21020),
            .I(N__21013));
    LocalMux I__4169 (
            .O(N__21017),
            .I(N__21008));
    InMux I__4168 (
            .O(N__21016),
            .I(N__21005));
    InMux I__4167 (
            .O(N__21013),
            .I(N__21002));
    InMux I__4166 (
            .O(N__21012),
            .I(N__20999));
    InMux I__4165 (
            .O(N__21011),
            .I(N__20996));
    Span4Mux_h I__4164 (
            .O(N__21008),
            .I(N__20990));
    LocalMux I__4163 (
            .O(N__21005),
            .I(N__20990));
    LocalMux I__4162 (
            .O(N__21002),
            .I(N__20985));
    LocalMux I__4161 (
            .O(N__20999),
            .I(N__20985));
    LocalMux I__4160 (
            .O(N__20996),
            .I(N__20982));
    CascadeMux I__4159 (
            .O(N__20995),
            .I(N__20979));
    Span4Mux_v I__4158 (
            .O(N__20990),
            .I(N__20974));
    Span4Mux_v I__4157 (
            .O(N__20985),
            .I(N__20971));
    Span4Mux_h I__4156 (
            .O(N__20982),
            .I(N__20968));
    InMux I__4155 (
            .O(N__20979),
            .I(N__20965));
    InMux I__4154 (
            .O(N__20978),
            .I(N__20960));
    InMux I__4153 (
            .O(N__20977),
            .I(N__20960));
    Span4Mux_v I__4152 (
            .O(N__20974),
            .I(N__20957));
    Span4Mux_h I__4151 (
            .O(N__20971),
            .I(N__20952));
    Span4Mux_v I__4150 (
            .O(N__20968),
            .I(N__20952));
    LocalMux I__4149 (
            .O(N__20965),
            .I(N__20947));
    LocalMux I__4148 (
            .O(N__20960),
            .I(N__20947));
    Odrv4 I__4147 (
            .O(N__20957),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    Odrv4 I__4146 (
            .O(N__20952),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    Odrv12 I__4145 (
            .O(N__20947),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    InMux I__4144 (
            .O(N__20940),
            .I(N__20937));
    LocalMux I__4143 (
            .O(N__20937),
            .I(N__20934));
    Span4Mux_h I__4142 (
            .O(N__20934),
            .I(N__20931));
    Span4Mux_h I__4141 (
            .O(N__20931),
            .I(N__20928));
    Odrv4 I__4140 (
            .O(N__20928),
            .I(\this_sprites_ram.mem_out_bus5_3 ));
    InMux I__4139 (
            .O(N__20925),
            .I(N__20922));
    LocalMux I__4138 (
            .O(N__20922),
            .I(N__20919));
    Span4Mux_v I__4137 (
            .O(N__20919),
            .I(N__20916));
    Span4Mux_h I__4136 (
            .O(N__20916),
            .I(N__20913));
    Span4Mux_v I__4135 (
            .O(N__20913),
            .I(N__20910));
    Odrv4 I__4134 (
            .O(N__20910),
            .I(\this_sprites_ram.mem_out_bus1_3 ));
    InMux I__4133 (
            .O(N__20907),
            .I(N__20904));
    LocalMux I__4132 (
            .O(N__20904),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ));
    InMux I__4131 (
            .O(N__20901),
            .I(N__20895));
    InMux I__4130 (
            .O(N__20900),
            .I(N__20892));
    InMux I__4129 (
            .O(N__20899),
            .I(N__20889));
    InMux I__4128 (
            .O(N__20898),
            .I(N__20886));
    LocalMux I__4127 (
            .O(N__20895),
            .I(N__20883));
    LocalMux I__4126 (
            .O(N__20892),
            .I(N__20880));
    LocalMux I__4125 (
            .O(N__20889),
            .I(N__20875));
    LocalMux I__4124 (
            .O(N__20886),
            .I(N__20875));
    Odrv12 I__4123 (
            .O(N__20883),
            .I(M_this_state_qZ0Z_10));
    Odrv4 I__4122 (
            .O(N__20880),
            .I(M_this_state_qZ0Z_10));
    Odrv4 I__4121 (
            .O(N__20875),
            .I(M_this_state_qZ0Z_10));
    InMux I__4120 (
            .O(N__20868),
            .I(N__20865));
    LocalMux I__4119 (
            .O(N__20865),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    CascadeMux I__4118 (
            .O(N__20862),
            .I(N__20859));
    CascadeBuf I__4117 (
            .O(N__20859),
            .I(N__20856));
    CascadeMux I__4116 (
            .O(N__20856),
            .I(N__20853));
    InMux I__4115 (
            .O(N__20853),
            .I(N__20850));
    LocalMux I__4114 (
            .O(N__20850),
            .I(N__20847));
    Span4Mux_v I__4113 (
            .O(N__20847),
            .I(N__20843));
    CascadeMux I__4112 (
            .O(N__20846),
            .I(N__20839));
    Span4Mux_h I__4111 (
            .O(N__20843),
            .I(N__20834));
    InMux I__4110 (
            .O(N__20842),
            .I(N__20831));
    InMux I__4109 (
            .O(N__20839),
            .I(N__20826));
    InMux I__4108 (
            .O(N__20838),
            .I(N__20826));
    InMux I__4107 (
            .O(N__20837),
            .I(N__20823));
    Span4Mux_h I__4106 (
            .O(N__20834),
            .I(N__20820));
    LocalMux I__4105 (
            .O(N__20831),
            .I(M_this_ppu_oam_addr_3));
    LocalMux I__4104 (
            .O(N__20826),
            .I(M_this_ppu_oam_addr_3));
    LocalMux I__4103 (
            .O(N__20823),
            .I(M_this_ppu_oam_addr_3));
    Odrv4 I__4102 (
            .O(N__20820),
            .I(M_this_ppu_oam_addr_3));
    InMux I__4101 (
            .O(N__20811),
            .I(N__20807));
    InMux I__4100 (
            .O(N__20810),
            .I(N__20804));
    LocalMux I__4099 (
            .O(N__20807),
            .I(\this_ppu.N_144_4 ));
    LocalMux I__4098 (
            .O(N__20804),
            .I(\this_ppu.N_144_4 ));
    CascadeMux I__4097 (
            .O(N__20799),
            .I(N__20795));
    CascadeMux I__4096 (
            .O(N__20798),
            .I(N__20792));
    InMux I__4095 (
            .O(N__20795),
            .I(N__20789));
    InMux I__4094 (
            .O(N__20792),
            .I(N__20786));
    LocalMux I__4093 (
            .O(N__20789),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    LocalMux I__4092 (
            .O(N__20786),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    InMux I__4091 (
            .O(N__20781),
            .I(N__20778));
    LocalMux I__4090 (
            .O(N__20778),
            .I(N__20775));
    Sp12to4 I__4089 (
            .O(N__20775),
            .I(N__20772));
    Odrv12 I__4088 (
            .O(N__20772),
            .I(\this_ppu.N_144 ));
    InMux I__4087 (
            .O(N__20769),
            .I(N__20766));
    LocalMux I__4086 (
            .O(N__20766),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ));
    InMux I__4085 (
            .O(N__20763),
            .I(N__20760));
    LocalMux I__4084 (
            .O(N__20760),
            .I(N__20757));
    Span4Mux_v I__4083 (
            .O(N__20757),
            .I(N__20754));
    Span4Mux_h I__4082 (
            .O(N__20754),
            .I(N__20751));
    Span4Mux_h I__4081 (
            .O(N__20751),
            .I(N__20748));
    Span4Mux_h I__4080 (
            .O(N__20748),
            .I(N__20745));
    Odrv4 I__4079 (
            .O(N__20745),
            .I(M_this_ppu_vram_data_0));
    CascadeMux I__4078 (
            .O(N__20742),
            .I(M_this_ppu_vram_data_0_cascade_));
    CascadeMux I__4077 (
            .O(N__20739),
            .I(\this_ppu.N_156_cascade_ ));
    CEMux I__4076 (
            .O(N__20736),
            .I(N__20733));
    LocalMux I__4075 (
            .O(N__20733),
            .I(N__20730));
    Span4Mux_v I__4074 (
            .O(N__20730),
            .I(N__20727));
    Span4Mux_v I__4073 (
            .O(N__20727),
            .I(N__20724));
    Span4Mux_h I__4072 (
            .O(N__20724),
            .I(N__20719));
    InMux I__4071 (
            .O(N__20723),
            .I(N__20716));
    InMux I__4070 (
            .O(N__20722),
            .I(N__20712));
    Span4Mux_h I__4069 (
            .O(N__20719),
            .I(N__20707));
    LocalMux I__4068 (
            .O(N__20716),
            .I(N__20707));
    InMux I__4067 (
            .O(N__20715),
            .I(N__20704));
    LocalMux I__4066 (
            .O(N__20712),
            .I(M_this_ppu_vram_en_0));
    Odrv4 I__4065 (
            .O(N__20707),
            .I(M_this_ppu_vram_en_0));
    LocalMux I__4064 (
            .O(N__20704),
            .I(M_this_ppu_vram_en_0));
    InMux I__4063 (
            .O(N__20697),
            .I(N__20694));
    LocalMux I__4062 (
            .O(N__20694),
            .I(N__20691));
    Span4Mux_h I__4061 (
            .O(N__20691),
            .I(N__20688));
    Span4Mux_v I__4060 (
            .O(N__20688),
            .I(N__20685));
    Span4Mux_h I__4059 (
            .O(N__20685),
            .I(N__20682));
    Odrv4 I__4058 (
            .O(N__20682),
            .I(\this_sprites_ram.mem_out_bus6_3 ));
    InMux I__4057 (
            .O(N__20679),
            .I(N__20676));
    LocalMux I__4056 (
            .O(N__20676),
            .I(N__20673));
    Span12Mux_h I__4055 (
            .O(N__20673),
            .I(N__20670));
    Odrv12 I__4054 (
            .O(N__20670),
            .I(\this_sprites_ram.mem_out_bus2_3 ));
    InMux I__4053 (
            .O(N__20667),
            .I(N__20664));
    LocalMux I__4052 (
            .O(N__20664),
            .I(N__20661));
    Span4Mux_v I__4051 (
            .O(N__20661),
            .I(N__20658));
    Sp12to4 I__4050 (
            .O(N__20658),
            .I(N__20655));
    Odrv12 I__4049 (
            .O(N__20655),
            .I(\this_sprites_ram.mem_out_bus4_0 ));
    InMux I__4048 (
            .O(N__20652),
            .I(N__20649));
    LocalMux I__4047 (
            .O(N__20649),
            .I(N__20646));
    Span4Mux_v I__4046 (
            .O(N__20646),
            .I(N__20643));
    Span4Mux_h I__4045 (
            .O(N__20643),
            .I(N__20640));
    Span4Mux_v I__4044 (
            .O(N__20640),
            .I(N__20637));
    Span4Mux_v I__4043 (
            .O(N__20637),
            .I(N__20634));
    Odrv4 I__4042 (
            .O(N__20634),
            .I(\this_sprites_ram.mem_out_bus0_0 ));
    CascadeMux I__4041 (
            .O(N__20631),
            .I(N__20628));
    CascadeBuf I__4040 (
            .O(N__20628),
            .I(N__20625));
    CascadeMux I__4039 (
            .O(N__20625),
            .I(N__20622));
    InMux I__4038 (
            .O(N__20622),
            .I(N__20619));
    LocalMux I__4037 (
            .O(N__20619),
            .I(N__20615));
    CascadeMux I__4036 (
            .O(N__20618),
            .I(N__20611));
    Span4Mux_h I__4035 (
            .O(N__20615),
            .I(N__20608));
    InMux I__4034 (
            .O(N__20614),
            .I(N__20605));
    InMux I__4033 (
            .O(N__20611),
            .I(N__20602));
    Sp12to4 I__4032 (
            .O(N__20608),
            .I(N__20599));
    LocalMux I__4031 (
            .O(N__20605),
            .I(N__20594));
    LocalMux I__4030 (
            .O(N__20602),
            .I(N__20591));
    Span12Mux_v I__4029 (
            .O(N__20599),
            .I(N__20588));
    InMux I__4028 (
            .O(N__20598),
            .I(N__20585));
    InMux I__4027 (
            .O(N__20597),
            .I(N__20582));
    Span12Mux_v I__4026 (
            .O(N__20594),
            .I(N__20575));
    Span12Mux_h I__4025 (
            .O(N__20591),
            .I(N__20575));
    Span12Mux_h I__4024 (
            .O(N__20588),
            .I(N__20575));
    LocalMux I__4023 (
            .O(N__20585),
            .I(M_this_ppu_map_addr_1));
    LocalMux I__4022 (
            .O(N__20582),
            .I(M_this_ppu_map_addr_1));
    Odrv12 I__4021 (
            .O(N__20575),
            .I(M_this_ppu_map_addr_1));
    CascadeMux I__4020 (
            .O(N__20568),
            .I(N__20565));
    CascadeBuf I__4019 (
            .O(N__20565),
            .I(N__20562));
    CascadeMux I__4018 (
            .O(N__20562),
            .I(N__20558));
    CascadeMux I__4017 (
            .O(N__20561),
            .I(N__20555));
    InMux I__4016 (
            .O(N__20558),
            .I(N__20552));
    InMux I__4015 (
            .O(N__20555),
            .I(N__20549));
    LocalMux I__4014 (
            .O(N__20552),
            .I(N__20546));
    LocalMux I__4013 (
            .O(N__20549),
            .I(N__20542));
    Span4Mux_h I__4012 (
            .O(N__20546),
            .I(N__20539));
    InMux I__4011 (
            .O(N__20545),
            .I(N__20536));
    Span4Mux_h I__4010 (
            .O(N__20542),
            .I(N__20533));
    Span4Mux_v I__4009 (
            .O(N__20539),
            .I(N__20530));
    LocalMux I__4008 (
            .O(N__20536),
            .I(N__20524));
    Span4Mux_v I__4007 (
            .O(N__20533),
            .I(N__20521));
    Sp12to4 I__4006 (
            .O(N__20530),
            .I(N__20518));
    InMux I__4005 (
            .O(N__20529),
            .I(N__20515));
    InMux I__4004 (
            .O(N__20528),
            .I(N__20512));
    InMux I__4003 (
            .O(N__20527),
            .I(N__20509));
    Span12Mux_h I__4002 (
            .O(N__20524),
            .I(N__20506));
    Sp12to4 I__4001 (
            .O(N__20521),
            .I(N__20501));
    Span12Mux_v I__4000 (
            .O(N__20518),
            .I(N__20501));
    LocalMux I__3999 (
            .O(N__20515),
            .I(M_this_ppu_map_addr_2));
    LocalMux I__3998 (
            .O(N__20512),
            .I(M_this_ppu_map_addr_2));
    LocalMux I__3997 (
            .O(N__20509),
            .I(M_this_ppu_map_addr_2));
    Odrv12 I__3996 (
            .O(N__20506),
            .I(M_this_ppu_map_addr_2));
    Odrv12 I__3995 (
            .O(N__20501),
            .I(M_this_ppu_map_addr_2));
    CascadeMux I__3994 (
            .O(N__20490),
            .I(N__20487));
    CascadeBuf I__3993 (
            .O(N__20487),
            .I(N__20484));
    CascadeMux I__3992 (
            .O(N__20484),
            .I(N__20481));
    InMux I__3991 (
            .O(N__20481),
            .I(N__20477));
    CascadeMux I__3990 (
            .O(N__20480),
            .I(N__20474));
    LocalMux I__3989 (
            .O(N__20477),
            .I(N__20471));
    InMux I__3988 (
            .O(N__20474),
            .I(N__20468));
    Span4Mux_v I__3987 (
            .O(N__20471),
            .I(N__20464));
    LocalMux I__3986 (
            .O(N__20468),
            .I(N__20461));
    InMux I__3985 (
            .O(N__20467),
            .I(N__20458));
    Sp12to4 I__3984 (
            .O(N__20464),
            .I(N__20455));
    Span4Mux_v I__3983 (
            .O(N__20461),
            .I(N__20450));
    LocalMux I__3982 (
            .O(N__20458),
            .I(N__20445));
    Span12Mux_h I__3981 (
            .O(N__20455),
            .I(N__20445));
    InMux I__3980 (
            .O(N__20454),
            .I(N__20442));
    InMux I__3979 (
            .O(N__20453),
            .I(N__20439));
    Sp12to4 I__3978 (
            .O(N__20450),
            .I(N__20436));
    Span12Mux_v I__3977 (
            .O(N__20445),
            .I(N__20433));
    LocalMux I__3976 (
            .O(N__20442),
            .I(M_this_ppu_map_addr_3));
    LocalMux I__3975 (
            .O(N__20439),
            .I(M_this_ppu_map_addr_3));
    Odrv12 I__3974 (
            .O(N__20436),
            .I(M_this_ppu_map_addr_3));
    Odrv12 I__3973 (
            .O(N__20433),
            .I(M_this_ppu_map_addr_3));
    CascadeMux I__3972 (
            .O(N__20424),
            .I(N__20421));
    CascadeBuf I__3971 (
            .O(N__20421),
            .I(N__20418));
    CascadeMux I__3970 (
            .O(N__20418),
            .I(N__20415));
    InMux I__3969 (
            .O(N__20415),
            .I(N__20412));
    LocalMux I__3968 (
            .O(N__20412),
            .I(N__20408));
    InMux I__3967 (
            .O(N__20411),
            .I(N__20405));
    Span4Mux_h I__3966 (
            .O(N__20408),
            .I(N__20402));
    LocalMux I__3965 (
            .O(N__20405),
            .I(N__20398));
    Sp12to4 I__3964 (
            .O(N__20402),
            .I(N__20395));
    CascadeMux I__3963 (
            .O(N__20401),
            .I(N__20392));
    Span4Mux_v I__3962 (
            .O(N__20398),
            .I(N__20389));
    Span12Mux_v I__3961 (
            .O(N__20395),
            .I(N__20386));
    InMux I__3960 (
            .O(N__20392),
            .I(N__20383));
    Span4Mux_v I__3959 (
            .O(N__20389),
            .I(N__20380));
    Span12Mux_h I__3958 (
            .O(N__20386),
            .I(N__20377));
    LocalMux I__3957 (
            .O(N__20383),
            .I(M_this_ppu_map_addr_4));
    Odrv4 I__3956 (
            .O(N__20380),
            .I(M_this_ppu_map_addr_4));
    Odrv12 I__3955 (
            .O(N__20377),
            .I(M_this_ppu_map_addr_4));
    InMux I__3954 (
            .O(N__20370),
            .I(bfn_18_20_0_));
    InMux I__3953 (
            .O(N__20367),
            .I(N__20363));
    InMux I__3952 (
            .O(N__20366),
            .I(N__20358));
    LocalMux I__3951 (
            .O(N__20363),
            .I(N__20355));
    InMux I__3950 (
            .O(N__20362),
            .I(N__20350));
    InMux I__3949 (
            .O(N__20361),
            .I(N__20350));
    LocalMux I__3948 (
            .O(N__20358),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__3947 (
            .O(N__20355),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    LocalMux I__3946 (
            .O(N__20350),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    CascadeMux I__3945 (
            .O(N__20343),
            .I(N__20340));
    InMux I__3944 (
            .O(N__20340),
            .I(N__20337));
    LocalMux I__3943 (
            .O(N__20337),
            .I(N__20334));
    Odrv4 I__3942 (
            .O(N__20334),
            .I(\this_ppu.un1_M_haddress_q_2_4 ));
    InMux I__3941 (
            .O(N__20331),
            .I(N__20328));
    LocalMux I__3940 (
            .O(N__20328),
            .I(\this_ppu.N_148 ));
    InMux I__3939 (
            .O(N__20325),
            .I(N__20320));
    InMux I__3938 (
            .O(N__20324),
            .I(N__20316));
    InMux I__3937 (
            .O(N__20323),
            .I(N__20313));
    LocalMux I__3936 (
            .O(N__20320),
            .I(N__20310));
    InMux I__3935 (
            .O(N__20319),
            .I(N__20307));
    LocalMux I__3934 (
            .O(N__20316),
            .I(\this_ppu.vscroll8 ));
    LocalMux I__3933 (
            .O(N__20313),
            .I(\this_ppu.vscroll8 ));
    Odrv4 I__3932 (
            .O(N__20310),
            .I(\this_ppu.vscroll8 ));
    LocalMux I__3931 (
            .O(N__20307),
            .I(\this_ppu.vscroll8 ));
    CascadeMux I__3930 (
            .O(N__20298),
            .I(N__20295));
    InMux I__3929 (
            .O(N__20295),
            .I(N__20292));
    LocalMux I__3928 (
            .O(N__20292),
            .I(N__20289));
    Odrv4 I__3927 (
            .O(N__20289),
            .I(\this_ppu.un1_M_haddress_q_2_5 ));
    CascadeMux I__3926 (
            .O(N__20286),
            .I(\this_ppu.un1_M_vaddress_q_2_c2_cascade_ ));
    InMux I__3925 (
            .O(N__20283),
            .I(N__20274));
    InMux I__3924 (
            .O(N__20282),
            .I(N__20274));
    InMux I__3923 (
            .O(N__20281),
            .I(N__20274));
    LocalMux I__3922 (
            .O(N__20274),
            .I(\this_ppu.un1_M_vaddress_q_2_c5 ));
    CascadeMux I__3921 (
            .O(N__20271),
            .I(N__20268));
    CascadeBuf I__3920 (
            .O(N__20268),
            .I(N__20265));
    CascadeMux I__3919 (
            .O(N__20265),
            .I(N__20261));
    CascadeMux I__3918 (
            .O(N__20264),
            .I(N__20258));
    InMux I__3917 (
            .O(N__20261),
            .I(N__20255));
    InMux I__3916 (
            .O(N__20258),
            .I(N__20252));
    LocalMux I__3915 (
            .O(N__20255),
            .I(N__20249));
    LocalMux I__3914 (
            .O(N__20252),
            .I(N__20245));
    Span4Mux_h I__3913 (
            .O(N__20249),
            .I(N__20242));
    InMux I__3912 (
            .O(N__20248),
            .I(N__20239));
    Span4Mux_v I__3911 (
            .O(N__20245),
            .I(N__20236));
    Sp12to4 I__3910 (
            .O(N__20242),
            .I(N__20233));
    LocalMux I__3909 (
            .O(N__20239),
            .I(N__20227));
    Sp12to4 I__3908 (
            .O(N__20236),
            .I(N__20224));
    Span12Mux_v I__3907 (
            .O(N__20233),
            .I(N__20221));
    InMux I__3906 (
            .O(N__20232),
            .I(N__20216));
    InMux I__3905 (
            .O(N__20231),
            .I(N__20216));
    InMux I__3904 (
            .O(N__20230),
            .I(N__20213));
    Span12Mux_v I__3903 (
            .O(N__20227),
            .I(N__20206));
    Span12Mux_h I__3902 (
            .O(N__20224),
            .I(N__20206));
    Span12Mux_h I__3901 (
            .O(N__20221),
            .I(N__20206));
    LocalMux I__3900 (
            .O(N__20216),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__3899 (
            .O(N__20213),
            .I(M_this_ppu_map_addr_0));
    Odrv12 I__3898 (
            .O(N__20206),
            .I(M_this_ppu_map_addr_0));
    InMux I__3897 (
            .O(N__20199),
            .I(M_this_data_count_q_cry_6));
    InMux I__3896 (
            .O(N__20196),
            .I(N__20193));
    LocalMux I__3895 (
            .O(N__20193),
            .I(N__20190));
    Odrv4 I__3894 (
            .O(N__20190),
            .I(M_this_data_count_q_cry_7_THRU_CO));
    InMux I__3893 (
            .O(N__20187),
            .I(bfn_18_16_0_));
    InMux I__3892 (
            .O(N__20184),
            .I(N__20181));
    LocalMux I__3891 (
            .O(N__20181),
            .I(N__20178));
    Odrv4 I__3890 (
            .O(N__20178),
            .I(M_this_data_count_q_cry_8_THRU_CO));
    InMux I__3889 (
            .O(N__20175),
            .I(M_this_data_count_q_cry_8));
    InMux I__3888 (
            .O(N__20172),
            .I(N__20168));
    InMux I__3887 (
            .O(N__20171),
            .I(N__20165));
    LocalMux I__3886 (
            .O(N__20168),
            .I(M_this_data_count_qZ0Z_10));
    LocalMux I__3885 (
            .O(N__20165),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__3884 (
            .O(N__20160),
            .I(N__20157));
    LocalMux I__3883 (
            .O(N__20157),
            .I(M_this_data_count_q_s_10));
    InMux I__3882 (
            .O(N__20154),
            .I(M_this_data_count_q_cry_9));
    CascadeMux I__3881 (
            .O(N__20151),
            .I(N__20148));
    InMux I__3880 (
            .O(N__20148),
            .I(N__20144));
    InMux I__3879 (
            .O(N__20147),
            .I(N__20140));
    LocalMux I__3878 (
            .O(N__20144),
            .I(N__20137));
    InMux I__3877 (
            .O(N__20143),
            .I(N__20134));
    LocalMux I__3876 (
            .O(N__20140),
            .I(M_this_data_count_qZ0Z_11));
    Odrv12 I__3875 (
            .O(N__20137),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__3874 (
            .O(N__20134),
            .I(M_this_data_count_qZ0Z_11));
    InMux I__3873 (
            .O(N__20127),
            .I(N__20124));
    LocalMux I__3872 (
            .O(N__20124),
            .I(N__20121));
    Odrv4 I__3871 (
            .O(N__20121),
            .I(M_this_data_count_q_cry_10_THRU_CO));
    InMux I__3870 (
            .O(N__20118),
            .I(M_this_data_count_q_cry_10));
    InMux I__3869 (
            .O(N__20115),
            .I(N__20110));
    InMux I__3868 (
            .O(N__20114),
            .I(N__20105));
    InMux I__3867 (
            .O(N__20113),
            .I(N__20105));
    LocalMux I__3866 (
            .O(N__20110),
            .I(M_this_data_count_qZ0Z_12));
    LocalMux I__3865 (
            .O(N__20105),
            .I(M_this_data_count_qZ0Z_12));
    SRMux I__3864 (
            .O(N__20100),
            .I(N__20093));
    SRMux I__3863 (
            .O(N__20099),
            .I(N__20088));
    SRMux I__3862 (
            .O(N__20098),
            .I(N__20077));
    SRMux I__3861 (
            .O(N__20097),
            .I(N__20072));
    SRMux I__3860 (
            .O(N__20096),
            .I(N__20069));
    LocalMux I__3859 (
            .O(N__20093),
            .I(N__20064));
    SRMux I__3858 (
            .O(N__20092),
            .I(N__20061));
    SRMux I__3857 (
            .O(N__20091),
            .I(N__20058));
    LocalMux I__3856 (
            .O(N__20088),
            .I(N__20053));
    SRMux I__3855 (
            .O(N__20087),
            .I(N__20050));
    SRMux I__3854 (
            .O(N__20086),
            .I(N__20047));
    SRMux I__3853 (
            .O(N__20085),
            .I(N__20043));
    CascadeMux I__3852 (
            .O(N__20084),
            .I(N__20038));
    CascadeMux I__3851 (
            .O(N__20083),
            .I(N__20035));
    CascadeMux I__3850 (
            .O(N__20082),
            .I(N__20031));
    CascadeMux I__3849 (
            .O(N__20081),
            .I(N__20027));
    SRMux I__3848 (
            .O(N__20080),
            .I(N__20024));
    LocalMux I__3847 (
            .O(N__20077),
            .I(N__20020));
    SRMux I__3846 (
            .O(N__20076),
            .I(N__20017));
    SRMux I__3845 (
            .O(N__20075),
            .I(N__20014));
    LocalMux I__3844 (
            .O(N__20072),
            .I(N__20007));
    LocalMux I__3843 (
            .O(N__20069),
            .I(N__20007));
    SRMux I__3842 (
            .O(N__20068),
            .I(N__20004));
    SRMux I__3841 (
            .O(N__20067),
            .I(N__20001));
    Span4Mux_s2_v I__3840 (
            .O(N__20064),
            .I(N__19994));
    LocalMux I__3839 (
            .O(N__20061),
            .I(N__19994));
    LocalMux I__3838 (
            .O(N__20058),
            .I(N__19994));
    SRMux I__3837 (
            .O(N__20057),
            .I(N__19991));
    SRMux I__3836 (
            .O(N__20056),
            .I(N__19988));
    Span4Mux_v I__3835 (
            .O(N__20053),
            .I(N__19979));
    LocalMux I__3834 (
            .O(N__20050),
            .I(N__19979));
    LocalMux I__3833 (
            .O(N__20047),
            .I(N__19979));
    SRMux I__3832 (
            .O(N__20046),
            .I(N__19976));
    LocalMux I__3831 (
            .O(N__20043),
            .I(N__19972));
    SRMux I__3830 (
            .O(N__20042),
            .I(N__19969));
    IoInMux I__3829 (
            .O(N__20041),
            .I(N__19965));
    InMux I__3828 (
            .O(N__20038),
            .I(N__19957));
    InMux I__3827 (
            .O(N__20035),
            .I(N__19957));
    InMux I__3826 (
            .O(N__20034),
            .I(N__19957));
    InMux I__3825 (
            .O(N__20031),
            .I(N__19950));
    InMux I__3824 (
            .O(N__20030),
            .I(N__19950));
    InMux I__3823 (
            .O(N__20027),
            .I(N__19950));
    LocalMux I__3822 (
            .O(N__20024),
            .I(N__19947));
    SRMux I__3821 (
            .O(N__20023),
            .I(N__19944));
    Span4Mux_v I__3820 (
            .O(N__20020),
            .I(N__19937));
    LocalMux I__3819 (
            .O(N__20017),
            .I(N__19937));
    LocalMux I__3818 (
            .O(N__20014),
            .I(N__19937));
    SRMux I__3817 (
            .O(N__20013),
            .I(N__19934));
    SRMux I__3816 (
            .O(N__20012),
            .I(N__19931));
    Span4Mux_v I__3815 (
            .O(N__20007),
            .I(N__19924));
    LocalMux I__3814 (
            .O(N__20004),
            .I(N__19924));
    LocalMux I__3813 (
            .O(N__20001),
            .I(N__19924));
    Span4Mux_v I__3812 (
            .O(N__19994),
            .I(N__19917));
    LocalMux I__3811 (
            .O(N__19991),
            .I(N__19917));
    LocalMux I__3810 (
            .O(N__19988),
            .I(N__19917));
    SRMux I__3809 (
            .O(N__19987),
            .I(N__19914));
    SRMux I__3808 (
            .O(N__19986),
            .I(N__19907));
    Span4Mux_v I__3807 (
            .O(N__19979),
            .I(N__19902));
    LocalMux I__3806 (
            .O(N__19976),
            .I(N__19902));
    SRMux I__3805 (
            .O(N__19975),
            .I(N__19899));
    Span4Mux_v I__3804 (
            .O(N__19972),
            .I(N__19894));
    LocalMux I__3803 (
            .O(N__19969),
            .I(N__19894));
    SRMux I__3802 (
            .O(N__19968),
            .I(N__19891));
    LocalMux I__3801 (
            .O(N__19965),
            .I(N__19888));
    SRMux I__3800 (
            .O(N__19964),
            .I(N__19884));
    LocalMux I__3799 (
            .O(N__19957),
            .I(N__19879));
    LocalMux I__3798 (
            .O(N__19950),
            .I(N__19879));
    Span4Mux_h I__3797 (
            .O(N__19947),
            .I(N__19874));
    LocalMux I__3796 (
            .O(N__19944),
            .I(N__19871));
    Span4Mux_v I__3795 (
            .O(N__19937),
            .I(N__19866));
    LocalMux I__3794 (
            .O(N__19934),
            .I(N__19866));
    LocalMux I__3793 (
            .O(N__19931),
            .I(N__19862));
    Span4Mux_v I__3792 (
            .O(N__19924),
            .I(N__19859));
    Span4Mux_v I__3791 (
            .O(N__19917),
            .I(N__19854));
    LocalMux I__3790 (
            .O(N__19914),
            .I(N__19854));
    SRMux I__3789 (
            .O(N__19913),
            .I(N__19851));
    CascadeMux I__3788 (
            .O(N__19912),
            .I(N__19846));
    CascadeMux I__3787 (
            .O(N__19911),
            .I(N__19842));
    CascadeMux I__3786 (
            .O(N__19910),
            .I(N__19838));
    LocalMux I__3785 (
            .O(N__19907),
            .I(N__19828));
    Span4Mux_h I__3784 (
            .O(N__19902),
            .I(N__19828));
    LocalMux I__3783 (
            .O(N__19899),
            .I(N__19828));
    Span4Mux_v I__3782 (
            .O(N__19894),
            .I(N__19823));
    LocalMux I__3781 (
            .O(N__19891),
            .I(N__19823));
    IoSpan4Mux I__3780 (
            .O(N__19888),
            .I(N__19819));
    SRMux I__3779 (
            .O(N__19887),
            .I(N__19816));
    LocalMux I__3778 (
            .O(N__19884),
            .I(N__19813));
    Span4Mux_h I__3777 (
            .O(N__19879),
            .I(N__19810));
    SRMux I__3776 (
            .O(N__19878),
            .I(N__19806));
    SRMux I__3775 (
            .O(N__19877),
            .I(N__19803));
    Span4Mux_v I__3774 (
            .O(N__19874),
            .I(N__19797));
    Span4Mux_h I__3773 (
            .O(N__19871),
            .I(N__19797));
    Span4Mux_v I__3772 (
            .O(N__19866),
            .I(N__19794));
    SRMux I__3771 (
            .O(N__19865),
            .I(N__19791));
    Span4Mux_s2_v I__3770 (
            .O(N__19862),
            .I(N__19788));
    Span4Mux_v I__3769 (
            .O(N__19859),
            .I(N__19781));
    Span4Mux_v I__3768 (
            .O(N__19854),
            .I(N__19781));
    LocalMux I__3767 (
            .O(N__19851),
            .I(N__19781));
    InMux I__3766 (
            .O(N__19850),
            .I(N__19766));
    InMux I__3765 (
            .O(N__19849),
            .I(N__19766));
    InMux I__3764 (
            .O(N__19846),
            .I(N__19766));
    InMux I__3763 (
            .O(N__19845),
            .I(N__19766));
    InMux I__3762 (
            .O(N__19842),
            .I(N__19766));
    InMux I__3761 (
            .O(N__19841),
            .I(N__19766));
    InMux I__3760 (
            .O(N__19838),
            .I(N__19766));
    CascadeMux I__3759 (
            .O(N__19837),
            .I(N__19762));
    CascadeMux I__3758 (
            .O(N__19836),
            .I(N__19759));
    CascadeMux I__3757 (
            .O(N__19835),
            .I(N__19755));
    Span4Mux_v I__3756 (
            .O(N__19828),
            .I(N__19750));
    Span4Mux_v I__3755 (
            .O(N__19823),
            .I(N__19750));
    SRMux I__3754 (
            .O(N__19822),
            .I(N__19747));
    Span4Mux_s2_h I__3753 (
            .O(N__19819),
            .I(N__19741));
    LocalMux I__3752 (
            .O(N__19816),
            .I(N__19738));
    Span4Mux_v I__3751 (
            .O(N__19813),
            .I(N__19733));
    Span4Mux_h I__3750 (
            .O(N__19810),
            .I(N__19733));
    SRMux I__3749 (
            .O(N__19809),
            .I(N__19730));
    LocalMux I__3748 (
            .O(N__19806),
            .I(N__19724));
    LocalMux I__3747 (
            .O(N__19803),
            .I(N__19724));
    SRMux I__3746 (
            .O(N__19802),
            .I(N__19721));
    Span4Mux_v I__3745 (
            .O(N__19797),
            .I(N__19714));
    Span4Mux_v I__3744 (
            .O(N__19794),
            .I(N__19714));
    LocalMux I__3743 (
            .O(N__19791),
            .I(N__19714));
    Span4Mux_h I__3742 (
            .O(N__19788),
            .I(N__19711));
    Span4Mux_h I__3741 (
            .O(N__19781),
            .I(N__19706));
    LocalMux I__3740 (
            .O(N__19766),
            .I(N__19706));
    InMux I__3739 (
            .O(N__19765),
            .I(N__19695));
    InMux I__3738 (
            .O(N__19762),
            .I(N__19695));
    InMux I__3737 (
            .O(N__19759),
            .I(N__19695));
    InMux I__3736 (
            .O(N__19758),
            .I(N__19695));
    InMux I__3735 (
            .O(N__19755),
            .I(N__19695));
    Span4Mux_v I__3734 (
            .O(N__19750),
            .I(N__19690));
    LocalMux I__3733 (
            .O(N__19747),
            .I(N__19690));
    SRMux I__3732 (
            .O(N__19746),
            .I(N__19687));
    SRMux I__3731 (
            .O(N__19745),
            .I(N__19684));
    SRMux I__3730 (
            .O(N__19744),
            .I(N__19681));
    Sp12to4 I__3729 (
            .O(N__19741),
            .I(N__19676));
    Sp12to4 I__3728 (
            .O(N__19738),
            .I(N__19676));
    Span4Mux_v I__3727 (
            .O(N__19733),
            .I(N__19671));
    LocalMux I__3726 (
            .O(N__19730),
            .I(N__19671));
    IoInMux I__3725 (
            .O(N__19729),
            .I(N__19668));
    Span4Mux_v I__3724 (
            .O(N__19724),
            .I(N__19662));
    LocalMux I__3723 (
            .O(N__19721),
            .I(N__19662));
    Span4Mux_h I__3722 (
            .O(N__19714),
            .I(N__19659));
    Sp12to4 I__3721 (
            .O(N__19711),
            .I(N__19655));
    Span4Mux_h I__3720 (
            .O(N__19706),
            .I(N__19650));
    LocalMux I__3719 (
            .O(N__19695),
            .I(N__19650));
    Span4Mux_h I__3718 (
            .O(N__19690),
            .I(N__19647));
    LocalMux I__3717 (
            .O(N__19687),
            .I(N__19642));
    LocalMux I__3716 (
            .O(N__19684),
            .I(N__19642));
    LocalMux I__3715 (
            .O(N__19681),
            .I(N__19639));
    Span12Mux_h I__3714 (
            .O(N__19676),
            .I(N__19636));
    Span4Mux_h I__3713 (
            .O(N__19671),
            .I(N__19633));
    LocalMux I__3712 (
            .O(N__19668),
            .I(N__19630));
    SRMux I__3711 (
            .O(N__19667),
            .I(N__19627));
    Span4Mux_v I__3710 (
            .O(N__19662),
            .I(N__19624));
    Span4Mux_v I__3709 (
            .O(N__19659),
            .I(N__19621));
    SRMux I__3708 (
            .O(N__19658),
            .I(N__19618));
    Span12Mux_v I__3707 (
            .O(N__19655),
            .I(N__19614));
    Span4Mux_v I__3706 (
            .O(N__19650),
            .I(N__19611));
    Span4Mux_v I__3705 (
            .O(N__19647),
            .I(N__19606));
    Span4Mux_v I__3704 (
            .O(N__19642),
            .I(N__19606));
    Span4Mux_v I__3703 (
            .O(N__19639),
            .I(N__19603));
    Span12Mux_h I__3702 (
            .O(N__19636),
            .I(N__19598));
    Sp12to4 I__3701 (
            .O(N__19633),
            .I(N__19598));
    IoSpan4Mux I__3700 (
            .O(N__19630),
            .I(N__19595));
    LocalMux I__3699 (
            .O(N__19627),
            .I(N__19592));
    Span4Mux_v I__3698 (
            .O(N__19624),
            .I(N__19585));
    Span4Mux_v I__3697 (
            .O(N__19621),
            .I(N__19585));
    LocalMux I__3696 (
            .O(N__19618),
            .I(N__19585));
    SRMux I__3695 (
            .O(N__19617),
            .I(N__19582));
    Span12Mux_h I__3694 (
            .O(N__19614),
            .I(N__19578));
    Sp12to4 I__3693 (
            .O(N__19611),
            .I(N__19575));
    Sp12to4 I__3692 (
            .O(N__19606),
            .I(N__19570));
    Sp12to4 I__3691 (
            .O(N__19603),
            .I(N__19570));
    Span12Mux_v I__3690 (
            .O(N__19598),
            .I(N__19567));
    IoSpan4Mux I__3689 (
            .O(N__19595),
            .I(N__19564));
    Span4Mux_v I__3688 (
            .O(N__19592),
            .I(N__19557));
    Span4Mux_v I__3687 (
            .O(N__19585),
            .I(N__19557));
    LocalMux I__3686 (
            .O(N__19582),
            .I(N__19557));
    SRMux I__3685 (
            .O(N__19581),
            .I(N__19554));
    Span12Mux_v I__3684 (
            .O(N__19578),
            .I(N__19551));
    Span12Mux_h I__3683 (
            .O(N__19575),
            .I(N__19548));
    Span12Mux_h I__3682 (
            .O(N__19570),
            .I(N__19543));
    Span12Mux_v I__3681 (
            .O(N__19567),
            .I(N__19543));
    Span4Mux_s2_h I__3680 (
            .O(N__19564),
            .I(N__19540));
    Span4Mux_v I__3679 (
            .O(N__19557),
            .I(N__19535));
    LocalMux I__3678 (
            .O(N__19554),
            .I(N__19535));
    Odrv12 I__3677 (
            .O(N__19551),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3676 (
            .O(N__19548),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3675 (
            .O(N__19543),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3674 (
            .O(N__19540),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3673 (
            .O(N__19535),
            .I(CONSTANT_ONE_NET));
    InMux I__3672 (
            .O(N__19524),
            .I(N__19521));
    LocalMux I__3671 (
            .O(N__19521),
            .I(M_this_data_count_q_cry_11_THRU_CO));
    InMux I__3670 (
            .O(N__19518),
            .I(M_this_data_count_q_cry_11));
    InMux I__3669 (
            .O(N__19515),
            .I(N__19511));
    CascadeMux I__3668 (
            .O(N__19514),
            .I(N__19508));
    LocalMux I__3667 (
            .O(N__19511),
            .I(N__19505));
    InMux I__3666 (
            .O(N__19508),
            .I(N__19502));
    Odrv4 I__3665 (
            .O(N__19505),
            .I(M_this_data_count_qZ0Z_13));
    LocalMux I__3664 (
            .O(N__19502),
            .I(M_this_data_count_qZ0Z_13));
    InMux I__3663 (
            .O(N__19497),
            .I(M_this_data_count_q_cry_12));
    InMux I__3662 (
            .O(N__19494),
            .I(N__19491));
    LocalMux I__3661 (
            .O(N__19491),
            .I(N__19488));
    Odrv4 I__3660 (
            .O(N__19488),
            .I(M_this_data_count_q_s_13));
    InMux I__3659 (
            .O(N__19485),
            .I(N__19482));
    LocalMux I__3658 (
            .O(N__19482),
            .I(N_49));
    CascadeMux I__3657 (
            .O(N__19479),
            .I(N__19476));
    InMux I__3656 (
            .O(N__19476),
            .I(N__19473));
    LocalMux I__3655 (
            .O(N__19473),
            .I(N__19470));
    Span4Mux_v I__3654 (
            .O(N__19470),
            .I(N__19467));
    Span4Mux_h I__3653 (
            .O(N__19467),
            .I(N__19464));
    Odrv4 I__3652 (
            .O(N__19464),
            .I(this_vga_signals_vvisibility_1));
    InMux I__3651 (
            .O(N__19461),
            .I(N__19458));
    LocalMux I__3650 (
            .O(N__19458),
            .I(N__19443));
    InMux I__3649 (
            .O(N__19457),
            .I(N__19440));
    InMux I__3648 (
            .O(N__19456),
            .I(N__19437));
    InMux I__3647 (
            .O(N__19455),
            .I(N__19428));
    InMux I__3646 (
            .O(N__19454),
            .I(N__19428));
    InMux I__3645 (
            .O(N__19453),
            .I(N__19428));
    InMux I__3644 (
            .O(N__19452),
            .I(N__19428));
    InMux I__3643 (
            .O(N__19451),
            .I(N__19417));
    InMux I__3642 (
            .O(N__19450),
            .I(N__19417));
    InMux I__3641 (
            .O(N__19449),
            .I(N__19417));
    InMux I__3640 (
            .O(N__19448),
            .I(N__19417));
    InMux I__3639 (
            .O(N__19447),
            .I(N__19417));
    InMux I__3638 (
            .O(N__19446),
            .I(N__19414));
    Odrv4 I__3637 (
            .O(N__19443),
            .I(N_686_i));
    LocalMux I__3636 (
            .O(N__19440),
            .I(N_686_i));
    LocalMux I__3635 (
            .O(N__19437),
            .I(N_686_i));
    LocalMux I__3634 (
            .O(N__19428),
            .I(N_686_i));
    LocalMux I__3633 (
            .O(N__19417),
            .I(N_686_i));
    LocalMux I__3632 (
            .O(N__19414),
            .I(N_686_i));
    CEMux I__3631 (
            .O(N__19401),
            .I(N__19398));
    LocalMux I__3630 (
            .O(N__19398),
            .I(N__19390));
    CEMux I__3629 (
            .O(N__19397),
            .I(N__19387));
    CEMux I__3628 (
            .O(N__19396),
            .I(N__19384));
    CEMux I__3627 (
            .O(N__19395),
            .I(N__19381));
    CEMux I__3626 (
            .O(N__19394),
            .I(N__19378));
    CEMux I__3625 (
            .O(N__19393),
            .I(N__19375));
    Odrv12 I__3624 (
            .O(N__19390),
            .I(M_this_data_count_qlde_i_i));
    LocalMux I__3623 (
            .O(N__19387),
            .I(M_this_data_count_qlde_i_i));
    LocalMux I__3622 (
            .O(N__19384),
            .I(M_this_data_count_qlde_i_i));
    LocalMux I__3621 (
            .O(N__19381),
            .I(M_this_data_count_qlde_i_i));
    LocalMux I__3620 (
            .O(N__19378),
            .I(M_this_data_count_qlde_i_i));
    LocalMux I__3619 (
            .O(N__19375),
            .I(M_this_data_count_qlde_i_i));
    InMux I__3618 (
            .O(N__19362),
            .I(N__19357));
    InMux I__3617 (
            .O(N__19361),
            .I(N__19352));
    InMux I__3616 (
            .O(N__19360),
            .I(N__19352));
    LocalMux I__3615 (
            .O(N__19357),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__3614 (
            .O(N__19352),
            .I(M_this_data_count_qZ0Z_0));
    CascadeMux I__3613 (
            .O(N__19347),
            .I(N__19344));
    InMux I__3612 (
            .O(N__19344),
            .I(N__19339));
    InMux I__3611 (
            .O(N__19343),
            .I(N__19334));
    InMux I__3610 (
            .O(N__19342),
            .I(N__19334));
    LocalMux I__3609 (
            .O(N__19339),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__3608 (
            .O(N__19334),
            .I(M_this_data_count_qZ0Z_1));
    InMux I__3607 (
            .O(N__19329),
            .I(N__19326));
    LocalMux I__3606 (
            .O(N__19326),
            .I(M_this_data_count_q_cry_0_THRU_CO));
    InMux I__3605 (
            .O(N__19323),
            .I(M_this_data_count_q_cry_0));
    InMux I__3604 (
            .O(N__19320),
            .I(N__19317));
    LocalMux I__3603 (
            .O(N__19317),
            .I(N__19312));
    InMux I__3602 (
            .O(N__19316),
            .I(N__19309));
    InMux I__3601 (
            .O(N__19315),
            .I(N__19306));
    Span4Mux_v I__3600 (
            .O(N__19312),
            .I(N__19303));
    LocalMux I__3599 (
            .O(N__19309),
            .I(N__19300));
    LocalMux I__3598 (
            .O(N__19306),
            .I(M_this_data_count_qZ0Z_2));
    Odrv4 I__3597 (
            .O(N__19303),
            .I(M_this_data_count_qZ0Z_2));
    Odrv4 I__3596 (
            .O(N__19300),
            .I(M_this_data_count_qZ0Z_2));
    InMux I__3595 (
            .O(N__19293),
            .I(N__19290));
    LocalMux I__3594 (
            .O(N__19290),
            .I(N__19287));
    Span4Mux_h I__3593 (
            .O(N__19287),
            .I(N__19284));
    Odrv4 I__3592 (
            .O(N__19284),
            .I(M_this_data_count_q_cry_1_THRU_CO));
    InMux I__3591 (
            .O(N__19281),
            .I(M_this_data_count_q_cry_1));
    CascadeMux I__3590 (
            .O(N__19278),
            .I(N__19275));
    InMux I__3589 (
            .O(N__19275),
            .I(N__19272));
    LocalMux I__3588 (
            .O(N__19272),
            .I(N__19267));
    CascadeMux I__3587 (
            .O(N__19271),
            .I(N__19264));
    InMux I__3586 (
            .O(N__19270),
            .I(N__19261));
    Span4Mux_h I__3585 (
            .O(N__19267),
            .I(N__19258));
    InMux I__3584 (
            .O(N__19264),
            .I(N__19255));
    LocalMux I__3583 (
            .O(N__19261),
            .I(M_this_data_count_qZ0Z_3));
    Odrv4 I__3582 (
            .O(N__19258),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__3581 (
            .O(N__19255),
            .I(M_this_data_count_qZ0Z_3));
    InMux I__3580 (
            .O(N__19248),
            .I(N__19245));
    LocalMux I__3579 (
            .O(N__19245),
            .I(N__19242));
    Odrv4 I__3578 (
            .O(N__19242),
            .I(M_this_data_count_q_cry_2_THRU_CO));
    InMux I__3577 (
            .O(N__19239),
            .I(M_this_data_count_q_cry_2));
    InMux I__3576 (
            .O(N__19236),
            .I(N__19233));
    LocalMux I__3575 (
            .O(N__19233),
            .I(M_this_data_count_q_cry_3_THRU_CO));
    InMux I__3574 (
            .O(N__19230),
            .I(M_this_data_count_q_cry_3));
    InMux I__3573 (
            .O(N__19227),
            .I(N__19224));
    LocalMux I__3572 (
            .O(N__19224),
            .I(N__19221));
    Span4Mux_h I__3571 (
            .O(N__19221),
            .I(N__19218));
    Odrv4 I__3570 (
            .O(N__19218),
            .I(M_this_data_count_q_cry_4_THRU_CO));
    InMux I__3569 (
            .O(N__19215),
            .I(M_this_data_count_q_cry_4));
    InMux I__3568 (
            .O(N__19212),
            .I(N__19208));
    InMux I__3567 (
            .O(N__19211),
            .I(N__19205));
    LocalMux I__3566 (
            .O(N__19208),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__3565 (
            .O(N__19205),
            .I(M_this_data_count_qZ0Z_6));
    InMux I__3564 (
            .O(N__19200),
            .I(N__19197));
    LocalMux I__3563 (
            .O(N__19197),
            .I(M_this_data_count_q_s_6));
    InMux I__3562 (
            .O(N__19194),
            .I(M_this_data_count_q_cry_5));
    CascadeMux I__3561 (
            .O(N__19191),
            .I(N__19188));
    InMux I__3560 (
            .O(N__19188),
            .I(N__19185));
    LocalMux I__3559 (
            .O(N__19185),
            .I(N__19180));
    InMux I__3558 (
            .O(N__19184),
            .I(N__19175));
    InMux I__3557 (
            .O(N__19183),
            .I(N__19175));
    Odrv4 I__3556 (
            .O(N__19180),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__3555 (
            .O(N__19175),
            .I(M_this_data_count_qZ0Z_7));
    InMux I__3554 (
            .O(N__19170),
            .I(N__19167));
    LocalMux I__3553 (
            .O(N__19167),
            .I(M_this_data_count_q_cry_6_THRU_CO));
    InMux I__3552 (
            .O(N__19164),
            .I(N__19158));
    InMux I__3551 (
            .O(N__19163),
            .I(N__19158));
    LocalMux I__3550 (
            .O(N__19158),
            .I(\this_ppu.un1_M_haddress_q_3_c2 ));
    SRMux I__3549 (
            .O(N__19155),
            .I(N__19151));
    SRMux I__3548 (
            .O(N__19154),
            .I(N__19148));
    LocalMux I__3547 (
            .O(N__19151),
            .I(N__19145));
    LocalMux I__3546 (
            .O(N__19148),
            .I(N__19142));
    Span4Mux_v I__3545 (
            .O(N__19145),
            .I(N__19134));
    Span4Mux_v I__3544 (
            .O(N__19142),
            .I(N__19134));
    SRMux I__3543 (
            .O(N__19141),
            .I(N__19131));
    SRMux I__3542 (
            .O(N__19140),
            .I(N__19128));
    SRMux I__3541 (
            .O(N__19139),
            .I(N__19125));
    Odrv4 I__3540 (
            .O(N__19134),
            .I(\this_ppu.M_state_q_RNIGL6V4Z0Z_0 ));
    LocalMux I__3539 (
            .O(N__19131),
            .I(\this_ppu.M_state_q_RNIGL6V4Z0Z_0 ));
    LocalMux I__3538 (
            .O(N__19128),
            .I(\this_ppu.M_state_q_RNIGL6V4Z0Z_0 ));
    LocalMux I__3537 (
            .O(N__19125),
            .I(\this_ppu.M_state_q_RNIGL6V4Z0Z_0 ));
    InMux I__3536 (
            .O(N__19116),
            .I(N__19113));
    LocalMux I__3535 (
            .O(N__19113),
            .I(N__19110));
    Span4Mux_v I__3534 (
            .O(N__19110),
            .I(N__19107));
    Sp12to4 I__3533 (
            .O(N__19107),
            .I(N__19104));
    Odrv12 I__3532 (
            .O(N__19104),
            .I(\this_sprites_ram.mem_out_bus4_3 ));
    InMux I__3531 (
            .O(N__19101),
            .I(N__19098));
    LocalMux I__3530 (
            .O(N__19098),
            .I(N__19095));
    Span4Mux_v I__3529 (
            .O(N__19095),
            .I(N__19092));
    Span4Mux_h I__3528 (
            .O(N__19092),
            .I(N__19089));
    Span4Mux_h I__3527 (
            .O(N__19089),
            .I(N__19086));
    Span4Mux_v I__3526 (
            .O(N__19086),
            .I(N__19083));
    Odrv4 I__3525 (
            .O(N__19083),
            .I(\this_sprites_ram.mem_out_bus0_3 ));
    CEMux I__3524 (
            .O(N__19080),
            .I(N__19077));
    LocalMux I__3523 (
            .O(N__19077),
            .I(N__19073));
    CEMux I__3522 (
            .O(N__19076),
            .I(N__19070));
    Span4Mux_v I__3521 (
            .O(N__19073),
            .I(N__19065));
    LocalMux I__3520 (
            .O(N__19070),
            .I(N__19065));
    Span4Mux_h I__3519 (
            .O(N__19065),
            .I(N__19062));
    Span4Mux_h I__3518 (
            .O(N__19062),
            .I(N__19059));
    Odrv4 I__3517 (
            .O(N__19059),
            .I(\this_sprites_ram.mem_WE_8 ));
    CascadeMux I__3516 (
            .O(N__19056),
            .I(N__19053));
    CascadeBuf I__3515 (
            .O(N__19053),
            .I(N__19050));
    CascadeMux I__3514 (
            .O(N__19050),
            .I(N__19047));
    InMux I__3513 (
            .O(N__19047),
            .I(N__19042));
    CascadeMux I__3512 (
            .O(N__19046),
            .I(N__19039));
    InMux I__3511 (
            .O(N__19045),
            .I(N__19035));
    LocalMux I__3510 (
            .O(N__19042),
            .I(N__19032));
    InMux I__3509 (
            .O(N__19039),
            .I(N__19029));
    InMux I__3508 (
            .O(N__19038),
            .I(N__19026));
    LocalMux I__3507 (
            .O(N__19035),
            .I(N__19023));
    Span12Mux_v I__3506 (
            .O(N__19032),
            .I(N__19020));
    LocalMux I__3505 (
            .O(N__19029),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__3504 (
            .O(N__19026),
            .I(M_this_ppu_oam_addr_2));
    Odrv4 I__3503 (
            .O(N__19023),
            .I(M_this_ppu_oam_addr_2));
    Odrv12 I__3502 (
            .O(N__19020),
            .I(M_this_ppu_oam_addr_2));
    CascadeMux I__3501 (
            .O(N__19011),
            .I(N__19008));
    CascadeBuf I__3500 (
            .O(N__19008),
            .I(N__19005));
    CascadeMux I__3499 (
            .O(N__19005),
            .I(N__19002));
    InMux I__3498 (
            .O(N__19002),
            .I(N__18999));
    LocalMux I__3497 (
            .O(N__18999),
            .I(N__18996));
    Sp12to4 I__3496 (
            .O(N__18996),
            .I(N__18989));
    InMux I__3495 (
            .O(N__18995),
            .I(N__18982));
    InMux I__3494 (
            .O(N__18994),
            .I(N__18982));
    InMux I__3493 (
            .O(N__18993),
            .I(N__18982));
    InMux I__3492 (
            .O(N__18992),
            .I(N__18979));
    Span12Mux_v I__3491 (
            .O(N__18989),
            .I(N__18976));
    LocalMux I__3490 (
            .O(N__18982),
            .I(M_this_ppu_oam_addr_1));
    LocalMux I__3489 (
            .O(N__18979),
            .I(M_this_ppu_oam_addr_1));
    Odrv12 I__3488 (
            .O(N__18976),
            .I(M_this_ppu_oam_addr_1));
    CascadeMux I__3487 (
            .O(N__18969),
            .I(N__18965));
    InMux I__3486 (
            .O(N__18968),
            .I(N__18962));
    InMux I__3485 (
            .O(N__18965),
            .I(N__18959));
    LocalMux I__3484 (
            .O(N__18962),
            .I(\this_ppu.M_oam_idx_qZ0Z_4 ));
    LocalMux I__3483 (
            .O(N__18959),
            .I(\this_ppu.M_oam_idx_qZ0Z_4 ));
    CascadeMux I__3482 (
            .O(N__18954),
            .I(N__18951));
    CascadeBuf I__3481 (
            .O(N__18951),
            .I(N__18948));
    CascadeMux I__3480 (
            .O(N__18948),
            .I(N__18945));
    InMux I__3479 (
            .O(N__18945),
            .I(N__18942));
    LocalMux I__3478 (
            .O(N__18942),
            .I(N__18938));
    CascadeMux I__3477 (
            .O(N__18941),
            .I(N__18934));
    Span4Mux_v I__3476 (
            .O(N__18938),
            .I(N__18930));
    InMux I__3475 (
            .O(N__18937),
            .I(N__18927));
    InMux I__3474 (
            .O(N__18934),
            .I(N__18922));
    InMux I__3473 (
            .O(N__18933),
            .I(N__18922));
    Span4Mux_h I__3472 (
            .O(N__18930),
            .I(N__18919));
    LocalMux I__3471 (
            .O(N__18927),
            .I(M_this_ppu_oam_addr_0));
    LocalMux I__3470 (
            .O(N__18922),
            .I(M_this_ppu_oam_addr_0));
    Odrv4 I__3469 (
            .O(N__18919),
            .I(M_this_ppu_oam_addr_0));
    CascadeMux I__3468 (
            .O(N__18912),
            .I(\this_ppu.un1_M_haddress_q_3_c2_cascade_ ));
    InMux I__3467 (
            .O(N__18909),
            .I(N__18904));
    InMux I__3466 (
            .O(N__18908),
            .I(N__18901));
    InMux I__3465 (
            .O(N__18907),
            .I(N__18898));
    LocalMux I__3464 (
            .O(N__18904),
            .I(\this_ppu.un1_M_haddress_q_3_c5 ));
    LocalMux I__3463 (
            .O(N__18901),
            .I(\this_ppu.un1_M_haddress_q_3_c5 ));
    LocalMux I__3462 (
            .O(N__18898),
            .I(\this_ppu.un1_M_haddress_q_3_c5 ));
    InMux I__3461 (
            .O(N__18891),
            .I(N__18888));
    LocalMux I__3460 (
            .O(N__18888),
            .I(N__18885));
    Span4Mux_h I__3459 (
            .O(N__18885),
            .I(N__18882));
    Span4Mux_h I__3458 (
            .O(N__18882),
            .I(N__18879));
    Sp12to4 I__3457 (
            .O(N__18879),
            .I(N__18876));
    Odrv12 I__3456 (
            .O(N__18876),
            .I(\this_sprites_ram.mem_out_bus7_0 ));
    InMux I__3455 (
            .O(N__18873),
            .I(N__18870));
    LocalMux I__3454 (
            .O(N__18870),
            .I(N__18867));
    Span12Mux_h I__3453 (
            .O(N__18867),
            .I(N__18864));
    Odrv12 I__3452 (
            .O(N__18864),
            .I(\this_sprites_ram.mem_out_bus3_0 ));
    CascadeMux I__3451 (
            .O(N__18861),
            .I(\this_ppu.un2_hscroll_axb_0_cascade_ ));
    CascadeMux I__3450 (
            .O(N__18858),
            .I(N__18855));
    InMux I__3449 (
            .O(N__18855),
            .I(N__18848));
    CascadeMux I__3448 (
            .O(N__18854),
            .I(N__18845));
    CascadeMux I__3447 (
            .O(N__18853),
            .I(N__18840));
    CascadeMux I__3446 (
            .O(N__18852),
            .I(N__18837));
    CascadeMux I__3445 (
            .O(N__18851),
            .I(N__18834));
    LocalMux I__3444 (
            .O(N__18848),
            .I(N__18826));
    InMux I__3443 (
            .O(N__18845),
            .I(N__18823));
    CascadeMux I__3442 (
            .O(N__18844),
            .I(N__18820));
    CascadeMux I__3441 (
            .O(N__18843),
            .I(N__18817));
    InMux I__3440 (
            .O(N__18840),
            .I(N__18813));
    InMux I__3439 (
            .O(N__18837),
            .I(N__18810));
    InMux I__3438 (
            .O(N__18834),
            .I(N__18807));
    CascadeMux I__3437 (
            .O(N__18833),
            .I(N__18804));
    CascadeMux I__3436 (
            .O(N__18832),
            .I(N__18800));
    CascadeMux I__3435 (
            .O(N__18831),
            .I(N__18797));
    CascadeMux I__3434 (
            .O(N__18830),
            .I(N__18794));
    CascadeMux I__3433 (
            .O(N__18829),
            .I(N__18791));
    Span4Mux_s0_v I__3432 (
            .O(N__18826),
            .I(N__18784));
    LocalMux I__3431 (
            .O(N__18823),
            .I(N__18784));
    InMux I__3430 (
            .O(N__18820),
            .I(N__18781));
    InMux I__3429 (
            .O(N__18817),
            .I(N__18778));
    CascadeMux I__3428 (
            .O(N__18816),
            .I(N__18775));
    LocalMux I__3427 (
            .O(N__18813),
            .I(N__18770));
    LocalMux I__3426 (
            .O(N__18810),
            .I(N__18770));
    LocalMux I__3425 (
            .O(N__18807),
            .I(N__18767));
    InMux I__3424 (
            .O(N__18804),
            .I(N__18764));
    CascadeMux I__3423 (
            .O(N__18803),
            .I(N__18761));
    InMux I__3422 (
            .O(N__18800),
            .I(N__18758));
    InMux I__3421 (
            .O(N__18797),
            .I(N__18755));
    InMux I__3420 (
            .O(N__18794),
            .I(N__18752));
    InMux I__3419 (
            .O(N__18791),
            .I(N__18749));
    CascadeMux I__3418 (
            .O(N__18790),
            .I(N__18746));
    CascadeMux I__3417 (
            .O(N__18789),
            .I(N__18743));
    Span4Mux_v I__3416 (
            .O(N__18784),
            .I(N__18738));
    LocalMux I__3415 (
            .O(N__18781),
            .I(N__18738));
    LocalMux I__3414 (
            .O(N__18778),
            .I(N__18735));
    InMux I__3413 (
            .O(N__18775),
            .I(N__18732));
    Span4Mux_v I__3412 (
            .O(N__18770),
            .I(N__18725));
    Span4Mux_h I__3411 (
            .O(N__18767),
            .I(N__18725));
    LocalMux I__3410 (
            .O(N__18764),
            .I(N__18725));
    InMux I__3409 (
            .O(N__18761),
            .I(N__18722));
    LocalMux I__3408 (
            .O(N__18758),
            .I(N__18719));
    LocalMux I__3407 (
            .O(N__18755),
            .I(N__18716));
    LocalMux I__3406 (
            .O(N__18752),
            .I(N__18711));
    LocalMux I__3405 (
            .O(N__18749),
            .I(N__18711));
    InMux I__3404 (
            .O(N__18746),
            .I(N__18708));
    InMux I__3403 (
            .O(N__18743),
            .I(N__18705));
    Span4Mux_h I__3402 (
            .O(N__18738),
            .I(N__18702));
    Span4Mux_v I__3401 (
            .O(N__18735),
            .I(N__18697));
    LocalMux I__3400 (
            .O(N__18732),
            .I(N__18697));
    Span4Mux_v I__3399 (
            .O(N__18725),
            .I(N__18692));
    LocalMux I__3398 (
            .O(N__18722),
            .I(N__18692));
    Span4Mux_h I__3397 (
            .O(N__18719),
            .I(N__18689));
    Span4Mux_v I__3396 (
            .O(N__18716),
            .I(N__18682));
    Span4Mux_v I__3395 (
            .O(N__18711),
            .I(N__18682));
    LocalMux I__3394 (
            .O(N__18708),
            .I(N__18682));
    LocalMux I__3393 (
            .O(N__18705),
            .I(N__18679));
    Span4Mux_v I__3392 (
            .O(N__18702),
            .I(N__18674));
    Span4Mux_h I__3391 (
            .O(N__18697),
            .I(N__18674));
    Span4Mux_h I__3390 (
            .O(N__18692),
            .I(N__18671));
    Span4Mux_v I__3389 (
            .O(N__18689),
            .I(N__18666));
    Span4Mux_h I__3388 (
            .O(N__18682),
            .I(N__18666));
    Span4Mux_h I__3387 (
            .O(N__18679),
            .I(N__18663));
    Span4Mux_h I__3386 (
            .O(N__18674),
            .I(N__18658));
    Span4Mux_h I__3385 (
            .O(N__18671),
            .I(N__18658));
    Span4Mux_h I__3384 (
            .O(N__18666),
            .I(N__18653));
    Span4Mux_h I__3383 (
            .O(N__18663),
            .I(N__18653));
    Odrv4 I__3382 (
            .O(N__18658),
            .I(M_this_ppu_sprites_addr_0));
    Odrv4 I__3381 (
            .O(N__18653),
            .I(M_this_ppu_sprites_addr_0));
    IoInMux I__3380 (
            .O(N__18648),
            .I(N__18644));
    IoInMux I__3379 (
            .O(N__18647),
            .I(N__18637));
    LocalMux I__3378 (
            .O(N__18644),
            .I(N__18633));
    IoInMux I__3377 (
            .O(N__18643),
            .I(N__18630));
    IoInMux I__3376 (
            .O(N__18642),
            .I(N__18627));
    IoInMux I__3375 (
            .O(N__18641),
            .I(N__18623));
    IoInMux I__3374 (
            .O(N__18640),
            .I(N__18620));
    LocalMux I__3373 (
            .O(N__18637),
            .I(N__18617));
    IoInMux I__3372 (
            .O(N__18636),
            .I(N__18614));
    IoSpan4Mux I__3371 (
            .O(N__18633),
            .I(N__18604));
    LocalMux I__3370 (
            .O(N__18630),
            .I(N__18604));
    LocalMux I__3369 (
            .O(N__18627),
            .I(N__18601));
    IoInMux I__3368 (
            .O(N__18626),
            .I(N__18598));
    LocalMux I__3367 (
            .O(N__18623),
            .I(N__18591));
    LocalMux I__3366 (
            .O(N__18620),
            .I(N__18591));
    IoSpan4Mux I__3365 (
            .O(N__18617),
            .I(N__18585));
    LocalMux I__3364 (
            .O(N__18614),
            .I(N__18585));
    IoInMux I__3363 (
            .O(N__18613),
            .I(N__18582));
    IoInMux I__3362 (
            .O(N__18612),
            .I(N__18579));
    IoInMux I__3361 (
            .O(N__18611),
            .I(N__18576));
    IoInMux I__3360 (
            .O(N__18610),
            .I(N__18573));
    IoInMux I__3359 (
            .O(N__18609),
            .I(N__18570));
    IoSpan4Mux I__3358 (
            .O(N__18604),
            .I(N__18563));
    IoSpan4Mux I__3357 (
            .O(N__18601),
            .I(N__18563));
    LocalMux I__3356 (
            .O(N__18598),
            .I(N__18563));
    IoInMux I__3355 (
            .O(N__18597),
            .I(N__18560));
    IoInMux I__3354 (
            .O(N__18596),
            .I(N__18557));
    IoSpan4Mux I__3353 (
            .O(N__18591),
            .I(N__18553));
    IoInMux I__3352 (
            .O(N__18590),
            .I(N__18550));
    IoSpan4Mux I__3351 (
            .O(N__18585),
            .I(N__18541));
    LocalMux I__3350 (
            .O(N__18582),
            .I(N__18541));
    LocalMux I__3349 (
            .O(N__18579),
            .I(N__18541));
    LocalMux I__3348 (
            .O(N__18576),
            .I(N__18541));
    LocalMux I__3347 (
            .O(N__18573),
            .I(N__18536));
    LocalMux I__3346 (
            .O(N__18570),
            .I(N__18536));
    IoSpan4Mux I__3345 (
            .O(N__18563),
            .I(N__18531));
    LocalMux I__3344 (
            .O(N__18560),
            .I(N__18531));
    LocalMux I__3343 (
            .O(N__18557),
            .I(N__18528));
    IoInMux I__3342 (
            .O(N__18556),
            .I(N__18525));
    Sp12to4 I__3341 (
            .O(N__18553),
            .I(N__18522));
    LocalMux I__3340 (
            .O(N__18550),
            .I(N__18519));
    IoSpan4Mux I__3339 (
            .O(N__18541),
            .I(N__18514));
    IoSpan4Mux I__3338 (
            .O(N__18536),
            .I(N__18514));
    IoSpan4Mux I__3337 (
            .O(N__18531),
            .I(N__18509));
    IoSpan4Mux I__3336 (
            .O(N__18528),
            .I(N__18509));
    LocalMux I__3335 (
            .O(N__18525),
            .I(N__18506));
    Span12Mux_s1_h I__3334 (
            .O(N__18522),
            .I(N__18503));
    IoSpan4Mux I__3333 (
            .O(N__18519),
            .I(N__18500));
    Span4Mux_s0_h I__3332 (
            .O(N__18514),
            .I(N__18497));
    Span4Mux_s2_v I__3331 (
            .O(N__18509),
            .I(N__18492));
    Span4Mux_s2_v I__3330 (
            .O(N__18506),
            .I(N__18492));
    Span12Mux_h I__3329 (
            .O(N__18503),
            .I(N__18489));
    Sp12to4 I__3328 (
            .O(N__18500),
            .I(N__18486));
    Span4Mux_h I__3327 (
            .O(N__18497),
            .I(N__18483));
    Span4Mux_v I__3326 (
            .O(N__18492),
            .I(N__18480));
    Span12Mux_v I__3325 (
            .O(N__18489),
            .I(N__18475));
    Span12Mux_s6_h I__3324 (
            .O(N__18486),
            .I(N__18475));
    Sp12to4 I__3323 (
            .O(N__18483),
            .I(N__18472));
    Span4Mux_v I__3322 (
            .O(N__18480),
            .I(N__18469));
    Odrv12 I__3321 (
            .O(N__18475),
            .I(port_dmab_c_i));
    Odrv12 I__3320 (
            .O(N__18472),
            .I(port_dmab_c_i));
    Odrv4 I__3319 (
            .O(N__18469),
            .I(port_dmab_c_i));
    CascadeMux I__3318 (
            .O(N__18462),
            .I(\this_ppu.un1_M_oam_idx_q_1_c1_cascade_ ));
    CascadeMux I__3317 (
            .O(N__18459),
            .I(\this_ppu.un1_M_oam_idx_q_1_c3_cascade_ ));
    InMux I__3316 (
            .O(N__18456),
            .I(N__18452));
    InMux I__3315 (
            .O(N__18455),
            .I(N__18449));
    LocalMux I__3314 (
            .O(N__18452),
            .I(N__18443));
    LocalMux I__3313 (
            .O(N__18449),
            .I(N__18443));
    InMux I__3312 (
            .O(N__18448),
            .I(N__18439));
    Span12Mux_v I__3311 (
            .O(N__18443),
            .I(N__18436));
    InMux I__3310 (
            .O(N__18442),
            .I(N__18433));
    LocalMux I__3309 (
            .O(N__18439),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_7 ));
    Odrv12 I__3308 (
            .O(N__18436),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_7 ));
    LocalMux I__3307 (
            .O(N__18433),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_7 ));
    InMux I__3306 (
            .O(N__18426),
            .I(N__18423));
    LocalMux I__3305 (
            .O(N__18423),
            .I(\this_ppu.un1_M_oam_idx_q_1_c3 ));
    InMux I__3304 (
            .O(N__18420),
            .I(N__18414));
    InMux I__3303 (
            .O(N__18419),
            .I(N__18414));
    LocalMux I__3302 (
            .O(N__18414),
            .I(\this_ppu.un1_M_oam_idx_q_1_c1 ));
    InMux I__3301 (
            .O(N__18411),
            .I(N__18407));
    InMux I__3300 (
            .O(N__18410),
            .I(N__18401));
    LocalMux I__3299 (
            .O(N__18407),
            .I(N__18398));
    InMux I__3298 (
            .O(N__18406),
            .I(N__18391));
    InMux I__3297 (
            .O(N__18405),
            .I(N__18391));
    InMux I__3296 (
            .O(N__18404),
            .I(N__18391));
    LocalMux I__3295 (
            .O(N__18401),
            .I(\this_ppu.N_1156_0 ));
    Odrv4 I__3294 (
            .O(N__18398),
            .I(\this_ppu.N_1156_0 ));
    LocalMux I__3293 (
            .O(N__18391),
            .I(\this_ppu.N_1156_0 ));
    InMux I__3292 (
            .O(N__18384),
            .I(N__18381));
    LocalMux I__3291 (
            .O(N__18381),
            .I(N__18378));
    Span4Mux_v I__3290 (
            .O(N__18378),
            .I(N__18374));
    InMux I__3289 (
            .O(N__18377),
            .I(N__18371));
    Odrv4 I__3288 (
            .O(N__18374),
            .I(\this_vga_signals.N_97 ));
    LocalMux I__3287 (
            .O(N__18371),
            .I(\this_vga_signals.N_97 ));
    InMux I__3286 (
            .O(N__18366),
            .I(N__18363));
    LocalMux I__3285 (
            .O(N__18363),
            .I(\this_vga_signals.M_this_state_q_srsts_0_0_a2_0_2_0 ));
    InMux I__3284 (
            .O(N__18360),
            .I(N__18357));
    LocalMux I__3283 (
            .O(N__18357),
            .I(\this_vga_signals.N_154 ));
    CascadeMux I__3282 (
            .O(N__18354),
            .I(\this_vga_signals.N_62_cascade_ ));
    InMux I__3281 (
            .O(N__18351),
            .I(N__18348));
    LocalMux I__3280 (
            .O(N__18348),
            .I(\this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0 ));
    InMux I__3279 (
            .O(N__18345),
            .I(N__18342));
    LocalMux I__3278 (
            .O(N__18342),
            .I(N__18339));
    Span4Mux_v I__3277 (
            .O(N__18339),
            .I(N__18336));
    Sp12to4 I__3276 (
            .O(N__18336),
            .I(N__18333));
    Span12Mux_h I__3275 (
            .O(N__18333),
            .I(N__18330));
    Odrv12 I__3274 (
            .O(N__18330),
            .I(M_this_map_ram_read_data_2));
    CascadeMux I__3273 (
            .O(N__18327),
            .I(N__18322));
    CascadeMux I__3272 (
            .O(N__18326),
            .I(N__18318));
    CascadeMux I__3271 (
            .O(N__18325),
            .I(N__18314));
    InMux I__3270 (
            .O(N__18322),
            .I(N__18310));
    CascadeMux I__3269 (
            .O(N__18321),
            .I(N__18307));
    InMux I__3268 (
            .O(N__18318),
            .I(N__18303));
    CascadeMux I__3267 (
            .O(N__18317),
            .I(N__18300));
    InMux I__3266 (
            .O(N__18314),
            .I(N__18296));
    CascadeMux I__3265 (
            .O(N__18313),
            .I(N__18293));
    LocalMux I__3264 (
            .O(N__18310),
            .I(N__18289));
    InMux I__3263 (
            .O(N__18307),
            .I(N__18286));
    CascadeMux I__3262 (
            .O(N__18306),
            .I(N__18283));
    LocalMux I__3261 (
            .O(N__18303),
            .I(N__18279));
    InMux I__3260 (
            .O(N__18300),
            .I(N__18276));
    CascadeMux I__3259 (
            .O(N__18299),
            .I(N__18273));
    LocalMux I__3258 (
            .O(N__18296),
            .I(N__18269));
    InMux I__3257 (
            .O(N__18293),
            .I(N__18266));
    CascadeMux I__3256 (
            .O(N__18292),
            .I(N__18263));
    Span4Mux_v I__3255 (
            .O(N__18289),
            .I(N__18256));
    LocalMux I__3254 (
            .O(N__18286),
            .I(N__18256));
    InMux I__3253 (
            .O(N__18283),
            .I(N__18253));
    CascadeMux I__3252 (
            .O(N__18282),
            .I(N__18250));
    Span4Mux_v I__3251 (
            .O(N__18279),
            .I(N__18243));
    LocalMux I__3250 (
            .O(N__18276),
            .I(N__18243));
    InMux I__3249 (
            .O(N__18273),
            .I(N__18240));
    CascadeMux I__3248 (
            .O(N__18272),
            .I(N__18237));
    Span4Mux_s0_v I__3247 (
            .O(N__18269),
            .I(N__18232));
    LocalMux I__3246 (
            .O(N__18266),
            .I(N__18232));
    InMux I__3245 (
            .O(N__18263),
            .I(N__18229));
    CascadeMux I__3244 (
            .O(N__18262),
            .I(N__18226));
    CascadeMux I__3243 (
            .O(N__18261),
            .I(N__18223));
    Span4Mux_h I__3242 (
            .O(N__18256),
            .I(N__18218));
    LocalMux I__3241 (
            .O(N__18253),
            .I(N__18218));
    InMux I__3240 (
            .O(N__18250),
            .I(N__18215));
    CascadeMux I__3239 (
            .O(N__18249),
            .I(N__18212));
    CascadeMux I__3238 (
            .O(N__18248),
            .I(N__18209));
    Span4Mux_v I__3237 (
            .O(N__18243),
            .I(N__18204));
    LocalMux I__3236 (
            .O(N__18240),
            .I(N__18204));
    InMux I__3235 (
            .O(N__18237),
            .I(N__18201));
    Span4Mux_v I__3234 (
            .O(N__18232),
            .I(N__18198));
    LocalMux I__3233 (
            .O(N__18229),
            .I(N__18195));
    InMux I__3232 (
            .O(N__18226),
            .I(N__18192));
    InMux I__3231 (
            .O(N__18223),
            .I(N__18189));
    Span4Mux_v I__3230 (
            .O(N__18218),
            .I(N__18184));
    LocalMux I__3229 (
            .O(N__18215),
            .I(N__18184));
    InMux I__3228 (
            .O(N__18212),
            .I(N__18181));
    InMux I__3227 (
            .O(N__18209),
            .I(N__18177));
    Span4Mux_h I__3226 (
            .O(N__18204),
            .I(N__18172));
    LocalMux I__3225 (
            .O(N__18201),
            .I(N__18172));
    Sp12to4 I__3224 (
            .O(N__18198),
            .I(N__18167));
    Sp12to4 I__3223 (
            .O(N__18195),
            .I(N__18167));
    LocalMux I__3222 (
            .O(N__18192),
            .I(N__18162));
    LocalMux I__3221 (
            .O(N__18189),
            .I(N__18162));
    Span4Mux_h I__3220 (
            .O(N__18184),
            .I(N__18157));
    LocalMux I__3219 (
            .O(N__18181),
            .I(N__18157));
    CascadeMux I__3218 (
            .O(N__18180),
            .I(N__18154));
    LocalMux I__3217 (
            .O(N__18177),
            .I(N__18151));
    Span4Mux_v I__3216 (
            .O(N__18172),
            .I(N__18148));
    Span12Mux_h I__3215 (
            .O(N__18167),
            .I(N__18145));
    Span4Mux_v I__3214 (
            .O(N__18162),
            .I(N__18140));
    Span4Mux_v I__3213 (
            .O(N__18157),
            .I(N__18140));
    InMux I__3212 (
            .O(N__18154),
            .I(N__18137));
    Span12Mux_h I__3211 (
            .O(N__18151),
            .I(N__18134));
    Sp12to4 I__3210 (
            .O(N__18148),
            .I(N__18131));
    Span12Mux_v I__3209 (
            .O(N__18145),
            .I(N__18124));
    Sp12to4 I__3208 (
            .O(N__18140),
            .I(N__18124));
    LocalMux I__3207 (
            .O(N__18137),
            .I(N__18124));
    Odrv12 I__3206 (
            .O(N__18134),
            .I(M_this_ppu_sprites_addr_8));
    Odrv12 I__3205 (
            .O(N__18131),
            .I(M_this_ppu_sprites_addr_8));
    Odrv12 I__3204 (
            .O(N__18124),
            .I(M_this_ppu_sprites_addr_8));
    InMux I__3203 (
            .O(N__18117),
            .I(N__18114));
    LocalMux I__3202 (
            .O(N__18114),
            .I(N__18111));
    Span4Mux_v I__3201 (
            .O(N__18111),
            .I(N__18108));
    Span4Mux_v I__3200 (
            .O(N__18108),
            .I(N__18105));
    Span4Mux_h I__3199 (
            .O(N__18105),
            .I(N__18102));
    Span4Mux_h I__3198 (
            .O(N__18102),
            .I(N__18099));
    Odrv4 I__3197 (
            .O(N__18099),
            .I(M_this_map_ram_read_data_1));
    CascadeMux I__3196 (
            .O(N__18096),
            .I(N__18093));
    InMux I__3195 (
            .O(N__18093),
            .I(N__18089));
    CascadeMux I__3194 (
            .O(N__18092),
            .I(N__18086));
    LocalMux I__3193 (
            .O(N__18089),
            .I(N__18082));
    InMux I__3192 (
            .O(N__18086),
            .I(N__18079));
    CascadeMux I__3191 (
            .O(N__18085),
            .I(N__18076));
    Span4Mux_h I__3190 (
            .O(N__18082),
            .I(N__18070));
    LocalMux I__3189 (
            .O(N__18079),
            .I(N__18070));
    InMux I__3188 (
            .O(N__18076),
            .I(N__18067));
    CascadeMux I__3187 (
            .O(N__18075),
            .I(N__18064));
    Span4Mux_v I__3186 (
            .O(N__18070),
            .I(N__18058));
    LocalMux I__3185 (
            .O(N__18067),
            .I(N__18058));
    InMux I__3184 (
            .O(N__18064),
            .I(N__18055));
    CascadeMux I__3183 (
            .O(N__18063),
            .I(N__18052));
    Span4Mux_h I__3182 (
            .O(N__18058),
            .I(N__18045));
    LocalMux I__3181 (
            .O(N__18055),
            .I(N__18045));
    InMux I__3180 (
            .O(N__18052),
            .I(N__18042));
    CascadeMux I__3179 (
            .O(N__18051),
            .I(N__18039));
    CascadeMux I__3178 (
            .O(N__18050),
            .I(N__18035));
    Span4Mux_v I__3177 (
            .O(N__18045),
            .I(N__18029));
    LocalMux I__3176 (
            .O(N__18042),
            .I(N__18029));
    InMux I__3175 (
            .O(N__18039),
            .I(N__18026));
    CascadeMux I__3174 (
            .O(N__18038),
            .I(N__18023));
    InMux I__3173 (
            .O(N__18035),
            .I(N__18014));
    CascadeMux I__3172 (
            .O(N__18034),
            .I(N__18011));
    Span4Mux_h I__3171 (
            .O(N__18029),
            .I(N__18006));
    LocalMux I__3170 (
            .O(N__18026),
            .I(N__18006));
    InMux I__3169 (
            .O(N__18023),
            .I(N__18003));
    CascadeMux I__3168 (
            .O(N__18022),
            .I(N__18000));
    CascadeMux I__3167 (
            .O(N__18021),
            .I(N__17996));
    CascadeMux I__3166 (
            .O(N__18020),
            .I(N__17993));
    CascadeMux I__3165 (
            .O(N__18019),
            .I(N__17990));
    CascadeMux I__3164 (
            .O(N__18018),
            .I(N__17987));
    CascadeMux I__3163 (
            .O(N__18017),
            .I(N__17984));
    LocalMux I__3162 (
            .O(N__18014),
            .I(N__17981));
    InMux I__3161 (
            .O(N__18011),
            .I(N__17978));
    Span4Mux_v I__3160 (
            .O(N__18006),
            .I(N__17973));
    LocalMux I__3159 (
            .O(N__18003),
            .I(N__17973));
    InMux I__3158 (
            .O(N__18000),
            .I(N__17970));
    CascadeMux I__3157 (
            .O(N__17999),
            .I(N__17967));
    InMux I__3156 (
            .O(N__17996),
            .I(N__17964));
    InMux I__3155 (
            .O(N__17993),
            .I(N__17961));
    InMux I__3154 (
            .O(N__17990),
            .I(N__17958));
    InMux I__3153 (
            .O(N__17987),
            .I(N__17955));
    InMux I__3152 (
            .O(N__17984),
            .I(N__17952));
    Span4Mux_h I__3151 (
            .O(N__17981),
            .I(N__17947));
    LocalMux I__3150 (
            .O(N__17978),
            .I(N__17947));
    Span4Mux_h I__3149 (
            .O(N__17973),
            .I(N__17942));
    LocalMux I__3148 (
            .O(N__17970),
            .I(N__17942));
    InMux I__3147 (
            .O(N__17967),
            .I(N__17939));
    LocalMux I__3146 (
            .O(N__17964),
            .I(N__17928));
    LocalMux I__3145 (
            .O(N__17961),
            .I(N__17928));
    LocalMux I__3144 (
            .O(N__17958),
            .I(N__17928));
    LocalMux I__3143 (
            .O(N__17955),
            .I(N__17928));
    LocalMux I__3142 (
            .O(N__17952),
            .I(N__17928));
    Span4Mux_v I__3141 (
            .O(N__17947),
            .I(N__17925));
    Span4Mux_v I__3140 (
            .O(N__17942),
            .I(N__17920));
    LocalMux I__3139 (
            .O(N__17939),
            .I(N__17920));
    Span12Mux_v I__3138 (
            .O(N__17928),
            .I(N__17917));
    Sp12to4 I__3137 (
            .O(N__17925),
            .I(N__17912));
    Sp12to4 I__3136 (
            .O(N__17920),
            .I(N__17912));
    Odrv12 I__3135 (
            .O(N__17917),
            .I(M_this_ppu_sprites_addr_7));
    Odrv12 I__3134 (
            .O(N__17912),
            .I(M_this_ppu_sprites_addr_7));
    InMux I__3133 (
            .O(N__17907),
            .I(N__17901));
    InMux I__3132 (
            .O(N__17906),
            .I(N__17901));
    LocalMux I__3131 (
            .O(N__17901),
            .I(N__17898));
    Span12Mux_h I__3130 (
            .O(N__17898),
            .I(N__17895));
    Span12Mux_v I__3129 (
            .O(N__17895),
            .I(N__17892));
    Odrv12 I__3128 (
            .O(N__17892),
            .I(port_address_in_7));
    IoInMux I__3127 (
            .O(N__17889),
            .I(N__17886));
    LocalMux I__3126 (
            .O(N__17886),
            .I(N__17883));
    Span12Mux_s3_h I__3125 (
            .O(N__17883),
            .I(N__17880));
    Span12Mux_h I__3124 (
            .O(N__17880),
            .I(N__17876));
    CascadeMux I__3123 (
            .O(N__17879),
            .I(N__17873));
    Span12Mux_v I__3122 (
            .O(N__17876),
            .I(N__17869));
    InMux I__3121 (
            .O(N__17873),
            .I(N__17864));
    InMux I__3120 (
            .O(N__17872),
            .I(N__17864));
    Odrv12 I__3119 (
            .O(N__17869),
            .I(led_c_1));
    LocalMux I__3118 (
            .O(N__17864),
            .I(led_c_1));
    InMux I__3117 (
            .O(N__17859),
            .I(N__17855));
    InMux I__3116 (
            .O(N__17858),
            .I(N__17852));
    LocalMux I__3115 (
            .O(N__17855),
            .I(N__17849));
    LocalMux I__3114 (
            .O(N__17852),
            .I(N__17846));
    Span4Mux_h I__3113 (
            .O(N__17849),
            .I(N__17843));
    Odrv4 I__3112 (
            .O(N__17846),
            .I(N_84));
    Odrv4 I__3111 (
            .O(N__17843),
            .I(N_84));
    CascadeMux I__3110 (
            .O(N__17838),
            .I(N__17833));
    InMux I__3109 (
            .O(N__17837),
            .I(N__17828));
    InMux I__3108 (
            .O(N__17836),
            .I(N__17823));
    InMux I__3107 (
            .O(N__17833),
            .I(N__17823));
    InMux I__3106 (
            .O(N__17832),
            .I(N__17819));
    InMux I__3105 (
            .O(N__17831),
            .I(N__17816));
    LocalMux I__3104 (
            .O(N__17828),
            .I(N__17810));
    LocalMux I__3103 (
            .O(N__17823),
            .I(N__17810));
    InMux I__3102 (
            .O(N__17822),
            .I(N__17807));
    LocalMux I__3101 (
            .O(N__17819),
            .I(N__17804));
    LocalMux I__3100 (
            .O(N__17816),
            .I(N__17801));
    InMux I__3099 (
            .O(N__17815),
            .I(N__17798));
    Span4Mux_v I__3098 (
            .O(N__17810),
            .I(N__17795));
    LocalMux I__3097 (
            .O(N__17807),
            .I(N__17792));
    Span4Mux_h I__3096 (
            .O(N__17804),
            .I(N__17785));
    Span4Mux_v I__3095 (
            .O(N__17801),
            .I(N__17785));
    LocalMux I__3094 (
            .O(N__17798),
            .I(N__17785));
    Span4Mux_v I__3093 (
            .O(N__17795),
            .I(N__17782));
    Span4Mux_v I__3092 (
            .O(N__17792),
            .I(N__17777));
    Span4Mux_v I__3091 (
            .O(N__17785),
            .I(N__17777));
    Sp12to4 I__3090 (
            .O(N__17782),
            .I(N__17772));
    Sp12to4 I__3089 (
            .O(N__17777),
            .I(N__17772));
    Span12Mux_h I__3088 (
            .O(N__17772),
            .I(N__17769));
    Odrv12 I__3087 (
            .O(N__17769),
            .I(port_address_in_1));
    CascadeMux I__3086 (
            .O(N__17766),
            .I(N__17762));
    InMux I__3085 (
            .O(N__17765),
            .I(N__17758));
    InMux I__3084 (
            .O(N__17762),
            .I(N__17750));
    InMux I__3083 (
            .O(N__17761),
            .I(N__17750));
    LocalMux I__3082 (
            .O(N__17758),
            .I(N__17747));
    InMux I__3081 (
            .O(N__17757),
            .I(N__17744));
    InMux I__3080 (
            .O(N__17756),
            .I(N__17741));
    InMux I__3079 (
            .O(N__17755),
            .I(N__17738));
    LocalMux I__3078 (
            .O(N__17750),
            .I(N__17734));
    Span4Mux_h I__3077 (
            .O(N__17747),
            .I(N__17727));
    LocalMux I__3076 (
            .O(N__17744),
            .I(N__17727));
    LocalMux I__3075 (
            .O(N__17741),
            .I(N__17727));
    LocalMux I__3074 (
            .O(N__17738),
            .I(N__17724));
    InMux I__3073 (
            .O(N__17737),
            .I(N__17721));
    Span4Mux_v I__3072 (
            .O(N__17734),
            .I(N__17718));
    Span4Mux_v I__3071 (
            .O(N__17727),
            .I(N__17715));
    Span4Mux_h I__3070 (
            .O(N__17724),
            .I(N__17710));
    LocalMux I__3069 (
            .O(N__17721),
            .I(N__17710));
    Span4Mux_v I__3068 (
            .O(N__17718),
            .I(N__17707));
    Span4Mux_v I__3067 (
            .O(N__17715),
            .I(N__17704));
    Sp12to4 I__3066 (
            .O(N__17710),
            .I(N__17701));
    Sp12to4 I__3065 (
            .O(N__17707),
            .I(N__17698));
    Sp12to4 I__3064 (
            .O(N__17704),
            .I(N__17693));
    Span12Mux_v I__3063 (
            .O(N__17701),
            .I(N__17693));
    Span12Mux_h I__3062 (
            .O(N__17698),
            .I(N__17690));
    Span12Mux_h I__3061 (
            .O(N__17693),
            .I(N__17687));
    Odrv12 I__3060 (
            .O(N__17690),
            .I(port_address_in_4));
    Odrv12 I__3059 (
            .O(N__17687),
            .I(port_address_in_4));
    InMux I__3058 (
            .O(N__17682),
            .I(N__17677));
    InMux I__3057 (
            .O(N__17681),
            .I(N__17672));
    InMux I__3056 (
            .O(N__17680),
            .I(N__17672));
    LocalMux I__3055 (
            .O(N__17677),
            .I(N__17665));
    LocalMux I__3054 (
            .O(N__17672),
            .I(N__17665));
    InMux I__3053 (
            .O(N__17671),
            .I(N__17662));
    InMux I__3052 (
            .O(N__17670),
            .I(N__17659));
    Span4Mux_v I__3051 (
            .O(N__17665),
            .I(N__17655));
    LocalMux I__3050 (
            .O(N__17662),
            .I(N__17652));
    LocalMux I__3049 (
            .O(N__17659),
            .I(N__17649));
    InMux I__3048 (
            .O(N__17658),
            .I(N__17646));
    Span4Mux_v I__3047 (
            .O(N__17655),
            .I(N__17642));
    Span4Mux_h I__3046 (
            .O(N__17652),
            .I(N__17635));
    Span4Mux_v I__3045 (
            .O(N__17649),
            .I(N__17635));
    LocalMux I__3044 (
            .O(N__17646),
            .I(N__17635));
    InMux I__3043 (
            .O(N__17645),
            .I(N__17632));
    Sp12to4 I__3042 (
            .O(N__17642),
            .I(N__17629));
    Span4Mux_v I__3041 (
            .O(N__17635),
            .I(N__17626));
    LocalMux I__3040 (
            .O(N__17632),
            .I(N__17623));
    Span12Mux_h I__3039 (
            .O(N__17629),
            .I(N__17618));
    Sp12to4 I__3038 (
            .O(N__17626),
            .I(N__17618));
    Span12Mux_v I__3037 (
            .O(N__17623),
            .I(N__17615));
    Odrv12 I__3036 (
            .O(N__17618),
            .I(port_address_in_0));
    Odrv12 I__3035 (
            .O(N__17615),
            .I(port_address_in_0));
    CascadeMux I__3034 (
            .O(N__17610),
            .I(N__17607));
    InMux I__3033 (
            .O(N__17607),
            .I(N__17603));
    InMux I__3032 (
            .O(N__17606),
            .I(N__17600));
    LocalMux I__3031 (
            .O(N__17603),
            .I(N__17597));
    LocalMux I__3030 (
            .O(N__17600),
            .I(N__17594));
    Span4Mux_v I__3029 (
            .O(N__17597),
            .I(N__17591));
    Span4Mux_h I__3028 (
            .O(N__17594),
            .I(N__17588));
    Odrv4 I__3027 (
            .O(N__17591),
            .I(N_36));
    Odrv4 I__3026 (
            .O(N__17588),
            .I(N_36));
    InMux I__3025 (
            .O(N__17583),
            .I(N__17569));
    InMux I__3024 (
            .O(N__17582),
            .I(N__17569));
    InMux I__3023 (
            .O(N__17581),
            .I(N__17560));
    InMux I__3022 (
            .O(N__17580),
            .I(N__17560));
    InMux I__3021 (
            .O(N__17579),
            .I(N__17560));
    InMux I__3020 (
            .O(N__17578),
            .I(N__17560));
    InMux I__3019 (
            .O(N__17577),
            .I(N__17551));
    InMux I__3018 (
            .O(N__17576),
            .I(N__17551));
    InMux I__3017 (
            .O(N__17575),
            .I(N__17551));
    InMux I__3016 (
            .O(N__17574),
            .I(N__17551));
    LocalMux I__3015 (
            .O(N__17569),
            .I(N__17547));
    LocalMux I__3014 (
            .O(N__17560),
            .I(N__17542));
    LocalMux I__3013 (
            .O(N__17551),
            .I(N__17542));
    CascadeMux I__3012 (
            .O(N__17550),
            .I(N__17539));
    Span4Mux_v I__3011 (
            .O(N__17547),
            .I(N__17534));
    Span4Mux_v I__3010 (
            .O(N__17542),
            .I(N__17534));
    InMux I__3009 (
            .O(N__17539),
            .I(N__17531));
    Sp12to4 I__3008 (
            .O(N__17534),
            .I(N__17528));
    LocalMux I__3007 (
            .O(N__17531),
            .I(N__17525));
    Span12Mux_h I__3006 (
            .O(N__17528),
            .I(N__17522));
    Odrv4 I__3005 (
            .O(N__17525),
            .I(N_164));
    Odrv12 I__3004 (
            .O(N__17522),
            .I(N_164));
    InMux I__3003 (
            .O(N__17517),
            .I(N__17514));
    LocalMux I__3002 (
            .O(N__17514),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_8 ));
    CascadeMux I__3001 (
            .O(N__17511),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_8_cascade_ ));
    InMux I__3000 (
            .O(N__17508),
            .I(N__17505));
    LocalMux I__2999 (
            .O(N__17505),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_8 ));
    InMux I__2998 (
            .O(N__17502),
            .I(N__17498));
    InMux I__2997 (
            .O(N__17501),
            .I(N__17495));
    LocalMux I__2996 (
            .O(N__17498),
            .I(N__17492));
    LocalMux I__2995 (
            .O(N__17495),
            .I(N__17489));
    Span4Mux_h I__2994 (
            .O(N__17492),
            .I(N__17486));
    Span4Mux_h I__2993 (
            .O(N__17489),
            .I(N__17483));
    Odrv4 I__2992 (
            .O(N__17486),
            .I(\this_vga_signals.N_124_0 ));
    Odrv4 I__2991 (
            .O(N__17483),
            .I(\this_vga_signals.N_124_0 ));
    CascadeMux I__2990 (
            .O(N__17478),
            .I(\this_vga_signals.N_154_cascade_ ));
    InMux I__2989 (
            .O(N__17475),
            .I(N__17472));
    LocalMux I__2988 (
            .O(N__17472),
            .I(N__17469));
    Span4Mux_h I__2987 (
            .O(N__17469),
            .I(N__17466));
    Odrv4 I__2986 (
            .O(N__17466),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    CascadeMux I__2985 (
            .O(N__17463),
            .I(\this_vga_signals.N_153_0_cascade_ ));
    CascadeMux I__2984 (
            .O(N__17460),
            .I(N_686_i_cascade_));
    CascadeMux I__2983 (
            .O(N__17457),
            .I(N__17454));
    InMux I__2982 (
            .O(N__17454),
            .I(N__17451));
    LocalMux I__2981 (
            .O(N__17451),
            .I(\this_vga_signals.M_this_state_q_srsts_i_1Z0Z_11 ));
    CascadeMux I__2980 (
            .O(N__17448),
            .I(N__17445));
    InMux I__2979 (
            .O(N__17445),
            .I(N__17442));
    LocalMux I__2978 (
            .O(N__17442),
            .I(N__17439));
    Odrv12 I__2977 (
            .O(N__17439),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0Z0Z_3 ));
    InMux I__2976 (
            .O(N__17436),
            .I(N__17429));
    CEMux I__2975 (
            .O(N__17435),
            .I(N__17424));
    CEMux I__2974 (
            .O(N__17434),
            .I(N__17421));
    CascadeMux I__2973 (
            .O(N__17433),
            .I(N__17418));
    InMux I__2972 (
            .O(N__17432),
            .I(N__17415));
    LocalMux I__2971 (
            .O(N__17429),
            .I(N__17412));
    InMux I__2970 (
            .O(N__17428),
            .I(N__17407));
    InMux I__2969 (
            .O(N__17427),
            .I(N__17407));
    LocalMux I__2968 (
            .O(N__17424),
            .I(N__17401));
    LocalMux I__2967 (
            .O(N__17421),
            .I(N__17401));
    InMux I__2966 (
            .O(N__17418),
            .I(N__17398));
    LocalMux I__2965 (
            .O(N__17415),
            .I(N__17394));
    Span4Mux_v I__2964 (
            .O(N__17412),
            .I(N__17389));
    LocalMux I__2963 (
            .O(N__17407),
            .I(N__17389));
    InMux I__2962 (
            .O(N__17406),
            .I(N__17386));
    Span4Mux_v I__2961 (
            .O(N__17401),
            .I(N__17379));
    LocalMux I__2960 (
            .O(N__17398),
            .I(N__17379));
    InMux I__2959 (
            .O(N__17397),
            .I(N__17376));
    Span4Mux_v I__2958 (
            .O(N__17394),
            .I(N__17368));
    Span4Mux_h I__2957 (
            .O(N__17389),
            .I(N__17368));
    LocalMux I__2956 (
            .O(N__17386),
            .I(N__17368));
    InMux I__2955 (
            .O(N__17385),
            .I(N__17363));
    InMux I__2954 (
            .O(N__17384),
            .I(N__17363));
    Span4Mux_v I__2953 (
            .O(N__17379),
            .I(N__17360));
    LocalMux I__2952 (
            .O(N__17376),
            .I(N__17357));
    InMux I__2951 (
            .O(N__17375),
            .I(N__17354));
    Span4Mux_h I__2950 (
            .O(N__17368),
            .I(N__17349));
    LocalMux I__2949 (
            .O(N__17363),
            .I(N__17349));
    Span4Mux_h I__2948 (
            .O(N__17360),
            .I(N__17346));
    Span12Mux_h I__2947 (
            .O(N__17357),
            .I(N__17341));
    LocalMux I__2946 (
            .O(N__17354),
            .I(N__17341));
    Span4Mux_v I__2945 (
            .O(N__17349),
            .I(N__17336));
    Span4Mux_h I__2944 (
            .O(N__17346),
            .I(N__17336));
    Odrv12 I__2943 (
            .O(N__17341),
            .I(M_this_state_d_0_sqmuxa_1));
    Odrv4 I__2942 (
            .O(N__17336),
            .I(M_this_state_d_0_sqmuxa_1));
    InMux I__2941 (
            .O(N__17331),
            .I(N__17328));
    LocalMux I__2940 (
            .O(N__17328),
            .I(N__17325));
    Span4Mux_h I__2939 (
            .O(N__17325),
            .I(N__17322));
    Span4Mux_h I__2938 (
            .O(N__17322),
            .I(N__17319));
    Odrv4 I__2937 (
            .O(N__17319),
            .I(M_this_map_ram_write_data_7));
    IoInMux I__2936 (
            .O(N__17316),
            .I(N__17313));
    LocalMux I__2935 (
            .O(N__17313),
            .I(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO));
    InMux I__2934 (
            .O(N__17310),
            .I(N__17302));
    InMux I__2933 (
            .O(N__17309),
            .I(N__17296));
    InMux I__2932 (
            .O(N__17308),
            .I(N__17289));
    InMux I__2931 (
            .O(N__17307),
            .I(N__17289));
    InMux I__2930 (
            .O(N__17306),
            .I(N__17289));
    CEMux I__2929 (
            .O(N__17305),
            .I(N__17279));
    LocalMux I__2928 (
            .O(N__17302),
            .I(N__17276));
    InMux I__2927 (
            .O(N__17301),
            .I(N__17273));
    InMux I__2926 (
            .O(N__17300),
            .I(N__17263));
    InMux I__2925 (
            .O(N__17299),
            .I(N__17263));
    LocalMux I__2924 (
            .O(N__17296),
            .I(N__17260));
    LocalMux I__2923 (
            .O(N__17289),
            .I(N__17257));
    InMux I__2922 (
            .O(N__17288),
            .I(N__17254));
    InMux I__2921 (
            .O(N__17287),
            .I(N__17248));
    InMux I__2920 (
            .O(N__17286),
            .I(N__17248));
    InMux I__2919 (
            .O(N__17285),
            .I(N__17243));
    InMux I__2918 (
            .O(N__17284),
            .I(N__17243));
    InMux I__2917 (
            .O(N__17283),
            .I(N__17240));
    InMux I__2916 (
            .O(N__17282),
            .I(N__17237));
    LocalMux I__2915 (
            .O(N__17279),
            .I(N__17234));
    Span4Mux_v I__2914 (
            .O(N__17276),
            .I(N__17229));
    LocalMux I__2913 (
            .O(N__17273),
            .I(N__17229));
    InMux I__2912 (
            .O(N__17272),
            .I(N__17226));
    InMux I__2911 (
            .O(N__17271),
            .I(N__17217));
    InMux I__2910 (
            .O(N__17270),
            .I(N__17217));
    InMux I__2909 (
            .O(N__17269),
            .I(N__17217));
    InMux I__2908 (
            .O(N__17268),
            .I(N__17217));
    LocalMux I__2907 (
            .O(N__17263),
            .I(N__17212));
    Span4Mux_h I__2906 (
            .O(N__17260),
            .I(N__17212));
    Span4Mux_h I__2905 (
            .O(N__17257),
            .I(N__17207));
    LocalMux I__2904 (
            .O(N__17254),
            .I(N__17207));
    InMux I__2903 (
            .O(N__17253),
            .I(N__17204));
    LocalMux I__2902 (
            .O(N__17248),
            .I(N__17195));
    LocalMux I__2901 (
            .O(N__17243),
            .I(N__17195));
    LocalMux I__2900 (
            .O(N__17240),
            .I(N__17195));
    LocalMux I__2899 (
            .O(N__17237),
            .I(N__17195));
    Span4Mux_h I__2898 (
            .O(N__17234),
            .I(N__17190));
    Span4Mux_h I__2897 (
            .O(N__17229),
            .I(N__17190));
    LocalMux I__2896 (
            .O(N__17226),
            .I(N__17187));
    LocalMux I__2895 (
            .O(N__17217),
            .I(N__17184));
    Span4Mux_v I__2894 (
            .O(N__17212),
            .I(N__17177));
    Span4Mux_v I__2893 (
            .O(N__17207),
            .I(N__17177));
    LocalMux I__2892 (
            .O(N__17204),
            .I(N__17177));
    Span4Mux_v I__2891 (
            .O(N__17195),
            .I(N__17174));
    Span4Mux_h I__2890 (
            .O(N__17190),
            .I(N__17169));
    Span4Mux_v I__2889 (
            .O(N__17187),
            .I(N__17169));
    Odrv12 I__2888 (
            .O(N__17184),
            .I(G_425));
    Odrv4 I__2887 (
            .O(N__17177),
            .I(G_425));
    Odrv4 I__2886 (
            .O(N__17174),
            .I(G_425));
    Odrv4 I__2885 (
            .O(N__17169),
            .I(G_425));
    IoInMux I__2884 (
            .O(N__17160),
            .I(N__17157));
    LocalMux I__2883 (
            .O(N__17157),
            .I(N__17154));
    Span12Mux_s1_v I__2882 (
            .O(N__17154),
            .I(N__17151));
    Odrv12 I__2881 (
            .O(N__17151),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ));
    InMux I__2880 (
            .O(N__17148),
            .I(N__17143));
    InMux I__2879 (
            .O(N__17147),
            .I(N__17138));
    InMux I__2878 (
            .O(N__17146),
            .I(N__17138));
    LocalMux I__2877 (
            .O(N__17143),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    LocalMux I__2876 (
            .O(N__17138),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    InMux I__2875 (
            .O(N__17133),
            .I(N__17129));
    InMux I__2874 (
            .O(N__17132),
            .I(N__17126));
    LocalMux I__2873 (
            .O(N__17129),
            .I(N__17123));
    LocalMux I__2872 (
            .O(N__17126),
            .I(\this_vga_signals.M_vcounter_d8 ));
    Odrv4 I__2871 (
            .O(N__17123),
            .I(\this_vga_signals.M_vcounter_d8 ));
    InMux I__2870 (
            .O(N__17118),
            .I(N__17112));
    CascadeMux I__2869 (
            .O(N__17117),
            .I(N__17109));
    InMux I__2868 (
            .O(N__17116),
            .I(N__17104));
    InMux I__2867 (
            .O(N__17115),
            .I(N__17101));
    LocalMux I__2866 (
            .O(N__17112),
            .I(N__17098));
    InMux I__2865 (
            .O(N__17109),
            .I(N__17095));
    InMux I__2864 (
            .O(N__17108),
            .I(N__17088));
    InMux I__2863 (
            .O(N__17107),
            .I(N__17088));
    LocalMux I__2862 (
            .O(N__17104),
            .I(N__17085));
    LocalMux I__2861 (
            .O(N__17101),
            .I(N__17078));
    Span4Mux_v I__2860 (
            .O(N__17098),
            .I(N__17078));
    LocalMux I__2859 (
            .O(N__17095),
            .I(N__17078));
    InMux I__2858 (
            .O(N__17094),
            .I(N__17075));
    InMux I__2857 (
            .O(N__17093),
            .I(N__17072));
    LocalMux I__2856 (
            .O(N__17088),
            .I(N__17068));
    Span4Mux_h I__2855 (
            .O(N__17085),
            .I(N__17062));
    Span4Mux_h I__2854 (
            .O(N__17078),
            .I(N__17062));
    LocalMux I__2853 (
            .O(N__17075),
            .I(N__17057));
    LocalMux I__2852 (
            .O(N__17072),
            .I(N__17057));
    InMux I__2851 (
            .O(N__17071),
            .I(N__17053));
    Span4Mux_h I__2850 (
            .O(N__17068),
            .I(N__17050));
    InMux I__2849 (
            .O(N__17067),
            .I(N__17047));
    Span4Mux_v I__2848 (
            .O(N__17062),
            .I(N__17044));
    Span12Mux_v I__2847 (
            .O(N__17057),
            .I(N__17041));
    InMux I__2846 (
            .O(N__17056),
            .I(N__17038));
    LocalMux I__2845 (
            .O(N__17053),
            .I(N__17035));
    Odrv4 I__2844 (
            .O(N__17050),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    LocalMux I__2843 (
            .O(N__17047),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__2842 (
            .O(N__17044),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv12 I__2841 (
            .O(N__17041),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    LocalMux I__2840 (
            .O(N__17038),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__2839 (
            .O(N__17035),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    CascadeMux I__2838 (
            .O(N__17022),
            .I(N__17019));
    InMux I__2837 (
            .O(N__17019),
            .I(N__17016));
    LocalMux I__2836 (
            .O(N__17016),
            .I(N__17012));
    CascadeMux I__2835 (
            .O(N__17015),
            .I(N__17009));
    Span4Mux_v I__2834 (
            .O(N__17012),
            .I(N__17006));
    InMux I__2833 (
            .O(N__17009),
            .I(N__17003));
    Span4Mux_h I__2832 (
            .O(N__17006),
            .I(N__16998));
    LocalMux I__2831 (
            .O(N__17003),
            .I(N__16998));
    Odrv4 I__2830 (
            .O(N__16998),
            .I(\this_vga_signals.un1_M_hcounter_d7_1_0 ));
    CEMux I__2829 (
            .O(N__16995),
            .I(N__16992));
    LocalMux I__2828 (
            .O(N__16992),
            .I(N__16988));
    CEMux I__2827 (
            .O(N__16991),
            .I(N__16985));
    Span4Mux_v I__2826 (
            .O(N__16988),
            .I(N__16980));
    LocalMux I__2825 (
            .O(N__16985),
            .I(N__16980));
    Span4Mux_h I__2824 (
            .O(N__16980),
            .I(N__16977));
    Span4Mux_h I__2823 (
            .O(N__16977),
            .I(N__16974));
    Odrv4 I__2822 (
            .O(N__16974),
            .I(\this_sprites_ram.mem_WE_6 ));
    InMux I__2821 (
            .O(N__16971),
            .I(N__16968));
    LocalMux I__2820 (
            .O(N__16968),
            .I(N__16965));
    Odrv4 I__2819 (
            .O(N__16965),
            .I(\this_vga_signals.M_this_state_q_srsts_i_i_1Z0Z_10 ));
    CEMux I__2818 (
            .O(N__16962),
            .I(N__16959));
    LocalMux I__2817 (
            .O(N__16959),
            .I(N__16956));
    Span4Mux_h I__2816 (
            .O(N__16956),
            .I(N__16952));
    CEMux I__2815 (
            .O(N__16955),
            .I(N__16949));
    Span4Mux_v I__2814 (
            .O(N__16952),
            .I(N__16946));
    LocalMux I__2813 (
            .O(N__16949),
            .I(N__16943));
    Span4Mux_h I__2812 (
            .O(N__16946),
            .I(N__16940));
    Span12Mux_v I__2811 (
            .O(N__16943),
            .I(N__16937));
    Odrv4 I__2810 (
            .O(N__16940),
            .I(\this_sprites_ram.mem_WE_10 ));
    Odrv12 I__2809 (
            .O(N__16937),
            .I(\this_sprites_ram.mem_WE_10 ));
    CascadeMux I__2808 (
            .O(N__16932),
            .I(N__16929));
    InMux I__2807 (
            .O(N__16929),
            .I(N__16925));
    InMux I__2806 (
            .O(N__16928),
            .I(N__16922));
    LocalMux I__2805 (
            .O(N__16925),
            .I(this_vga_signals_M_this_state_q_srsts_0_1_i_a2_0_0_1));
    LocalMux I__2804 (
            .O(N__16922),
            .I(this_vga_signals_M_this_state_q_srsts_0_1_i_a2_0_0_1));
    CascadeMux I__2803 (
            .O(N__16917),
            .I(N__16914));
    InMux I__2802 (
            .O(N__16914),
            .I(N__16911));
    LocalMux I__2801 (
            .O(N__16911),
            .I(N__16908));
    Span4Mux_h I__2800 (
            .O(N__16908),
            .I(N__16905));
    Odrv4 I__2799 (
            .O(N__16905),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_6 ));
    InMux I__2798 (
            .O(N__16902),
            .I(N__16893));
    InMux I__2797 (
            .O(N__16901),
            .I(N__16893));
    InMux I__2796 (
            .O(N__16900),
            .I(N__16888));
    InMux I__2795 (
            .O(N__16899),
            .I(N__16888));
    InMux I__2794 (
            .O(N__16898),
            .I(N__16885));
    LocalMux I__2793 (
            .O(N__16893),
            .I(\this_vga_signals.N_85 ));
    LocalMux I__2792 (
            .O(N__16888),
            .I(\this_vga_signals.N_85 ));
    LocalMux I__2791 (
            .O(N__16885),
            .I(\this_vga_signals.N_85 ));
    CascadeMux I__2790 (
            .O(N__16878),
            .I(N__16875));
    InMux I__2789 (
            .O(N__16875),
            .I(N__16872));
    LocalMux I__2788 (
            .O(N__16872),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_4 ));
    InMux I__2787 (
            .O(N__16869),
            .I(N__16865));
    InMux I__2786 (
            .O(N__16868),
            .I(N__16862));
    LocalMux I__2785 (
            .O(N__16865),
            .I(N__16856));
    LocalMux I__2784 (
            .O(N__16862),
            .I(N__16856));
    InMux I__2783 (
            .O(N__16861),
            .I(N__16853));
    Span4Mux_v I__2782 (
            .O(N__16856),
            .I(N__16850));
    LocalMux I__2781 (
            .O(N__16853),
            .I(N__16847));
    Span4Mux_h I__2780 (
            .O(N__16850),
            .I(N__16844));
    Odrv4 I__2779 (
            .O(N__16847),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    Odrv4 I__2778 (
            .O(N__16844),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    InMux I__2777 (
            .O(N__16839),
            .I(N__16836));
    LocalMux I__2776 (
            .O(N__16836),
            .I(N__16833));
    Odrv4 I__2775 (
            .O(N__16833),
            .I(\this_vga_signals.CO0 ));
    InMux I__2774 (
            .O(N__16830),
            .I(N__16824));
    InMux I__2773 (
            .O(N__16829),
            .I(N__16824));
    LocalMux I__2772 (
            .O(N__16824),
            .I(this_pixel_clk_M_counter_q_i_1));
    InMux I__2771 (
            .O(N__16821),
            .I(N__16816));
    InMux I__2770 (
            .O(N__16820),
            .I(N__16811));
    InMux I__2769 (
            .O(N__16819),
            .I(N__16811));
    LocalMux I__2768 (
            .O(N__16816),
            .I(this_pixel_clk_M_counter_q_0));
    LocalMux I__2767 (
            .O(N__16811),
            .I(this_pixel_clk_M_counter_q_0));
    CascadeMux I__2766 (
            .O(N__16806),
            .I(\this_vga_signals.N_152_0_cascade_ ));
    CascadeMux I__2765 (
            .O(N__16803),
            .I(N__16800));
    InMux I__2764 (
            .O(N__16800),
            .I(N__16797));
    LocalMux I__2763 (
            .O(N__16797),
            .I(N__16794));
    Odrv4 I__2762 (
            .O(N__16794),
            .I(\this_vga_signals.M_vcounter_d7lto8_1 ));
    InMux I__2761 (
            .O(N__16791),
            .I(N__16785));
    InMux I__2760 (
            .O(N__16790),
            .I(N__16785));
    LocalMux I__2759 (
            .O(N__16785),
            .I(\this_vga_signals.M_vcounter_d7lt8_0 ));
    CascadeMux I__2758 (
            .O(N__16782),
            .I(N__16772));
    InMux I__2757 (
            .O(N__16781),
            .I(N__16763));
    InMux I__2756 (
            .O(N__16780),
            .I(N__16763));
    InMux I__2755 (
            .O(N__16779),
            .I(N__16756));
    CascadeMux I__2754 (
            .O(N__16778),
            .I(N__16753));
    CascadeMux I__2753 (
            .O(N__16777),
            .I(N__16750));
    InMux I__2752 (
            .O(N__16776),
            .I(N__16747));
    InMux I__2751 (
            .O(N__16775),
            .I(N__16743));
    InMux I__2750 (
            .O(N__16772),
            .I(N__16738));
    InMux I__2749 (
            .O(N__16771),
            .I(N__16738));
    InMux I__2748 (
            .O(N__16770),
            .I(N__16731));
    InMux I__2747 (
            .O(N__16769),
            .I(N__16731));
    InMux I__2746 (
            .O(N__16768),
            .I(N__16731));
    LocalMux I__2745 (
            .O(N__16763),
            .I(N__16728));
    InMux I__2744 (
            .O(N__16762),
            .I(N__16723));
    InMux I__2743 (
            .O(N__16761),
            .I(N__16723));
    InMux I__2742 (
            .O(N__16760),
            .I(N__16718));
    InMux I__2741 (
            .O(N__16759),
            .I(N__16718));
    LocalMux I__2740 (
            .O(N__16756),
            .I(N__16712));
    InMux I__2739 (
            .O(N__16753),
            .I(N__16703));
    InMux I__2738 (
            .O(N__16750),
            .I(N__16703));
    LocalMux I__2737 (
            .O(N__16747),
            .I(N__16700));
    InMux I__2736 (
            .O(N__16746),
            .I(N__16697));
    LocalMux I__2735 (
            .O(N__16743),
            .I(N__16692));
    LocalMux I__2734 (
            .O(N__16738),
            .I(N__16692));
    LocalMux I__2733 (
            .O(N__16731),
            .I(N__16689));
    Span4Mux_v I__2732 (
            .O(N__16728),
            .I(N__16684));
    LocalMux I__2731 (
            .O(N__16723),
            .I(N__16684));
    LocalMux I__2730 (
            .O(N__16718),
            .I(N__16681));
    InMux I__2729 (
            .O(N__16717),
            .I(N__16676));
    InMux I__2728 (
            .O(N__16716),
            .I(N__16676));
    InMux I__2727 (
            .O(N__16715),
            .I(N__16673));
    Span4Mux_v I__2726 (
            .O(N__16712),
            .I(N__16670));
    InMux I__2725 (
            .O(N__16711),
            .I(N__16665));
    InMux I__2724 (
            .O(N__16710),
            .I(N__16665));
    InMux I__2723 (
            .O(N__16709),
            .I(N__16660));
    InMux I__2722 (
            .O(N__16708),
            .I(N__16660));
    LocalMux I__2721 (
            .O(N__16703),
            .I(N__16655));
    Span12Mux_s9_v I__2720 (
            .O(N__16700),
            .I(N__16655));
    LocalMux I__2719 (
            .O(N__16697),
            .I(N__16642));
    Span4Mux_v I__2718 (
            .O(N__16692),
            .I(N__16642));
    Span4Mux_h I__2717 (
            .O(N__16689),
            .I(N__16642));
    Span4Mux_h I__2716 (
            .O(N__16684),
            .I(N__16642));
    Span4Mux_v I__2715 (
            .O(N__16681),
            .I(N__16642));
    LocalMux I__2714 (
            .O(N__16676),
            .I(N__16642));
    LocalMux I__2713 (
            .O(N__16673),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2712 (
            .O(N__16670),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2711 (
            .O(N__16665),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2710 (
            .O(N__16660),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv12 I__2709 (
            .O(N__16655),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2708 (
            .O(N__16642),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    InMux I__2707 (
            .O(N__16629),
            .I(N__16624));
    InMux I__2706 (
            .O(N__16628),
            .I(N__16621));
    CascadeMux I__2705 (
            .O(N__16627),
            .I(N__16616));
    LocalMux I__2704 (
            .O(N__16624),
            .I(N__16611));
    LocalMux I__2703 (
            .O(N__16621),
            .I(N__16607));
    InMux I__2702 (
            .O(N__16620),
            .I(N__16604));
    CascadeMux I__2701 (
            .O(N__16619),
            .I(N__16599));
    InMux I__2700 (
            .O(N__16616),
            .I(N__16596));
    CascadeMux I__2699 (
            .O(N__16615),
            .I(N__16593));
    CascadeMux I__2698 (
            .O(N__16614),
            .I(N__16590));
    Span4Mux_h I__2697 (
            .O(N__16611),
            .I(N__16587));
    InMux I__2696 (
            .O(N__16610),
            .I(N__16584));
    Span4Mux_h I__2695 (
            .O(N__16607),
            .I(N__16581));
    LocalMux I__2694 (
            .O(N__16604),
            .I(N__16578));
    InMux I__2693 (
            .O(N__16603),
            .I(N__16573));
    InMux I__2692 (
            .O(N__16602),
            .I(N__16573));
    InMux I__2691 (
            .O(N__16599),
            .I(N__16570));
    LocalMux I__2690 (
            .O(N__16596),
            .I(N__16567));
    InMux I__2689 (
            .O(N__16593),
            .I(N__16564));
    InMux I__2688 (
            .O(N__16590),
            .I(N__16561));
    Odrv4 I__2687 (
            .O(N__16587),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2686 (
            .O(N__16584),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2685 (
            .O(N__16581),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2684 (
            .O(N__16578),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2683 (
            .O(N__16573),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2682 (
            .O(N__16570),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2681 (
            .O(N__16567),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2680 (
            .O(N__16564),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2679 (
            .O(N__16561),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    InMux I__2678 (
            .O(N__16542),
            .I(N__16533));
    InMux I__2677 (
            .O(N__16541),
            .I(N__16530));
    InMux I__2676 (
            .O(N__16540),
            .I(N__16523));
    InMux I__2675 (
            .O(N__16539),
            .I(N__16523));
    InMux I__2674 (
            .O(N__16538),
            .I(N__16523));
    InMux I__2673 (
            .O(N__16537),
            .I(N__16518));
    InMux I__2672 (
            .O(N__16536),
            .I(N__16518));
    LocalMux I__2671 (
            .O(N__16533),
            .I(N__16512));
    LocalMux I__2670 (
            .O(N__16530),
            .I(N__16503));
    LocalMux I__2669 (
            .O(N__16523),
            .I(N__16500));
    LocalMux I__2668 (
            .O(N__16518),
            .I(N__16497));
    InMux I__2667 (
            .O(N__16517),
            .I(N__16494));
    InMux I__2666 (
            .O(N__16516),
            .I(N__16491));
    InMux I__2665 (
            .O(N__16515),
            .I(N__16488));
    Span4Mux_v I__2664 (
            .O(N__16512),
            .I(N__16483));
    InMux I__2663 (
            .O(N__16511),
            .I(N__16478));
    InMux I__2662 (
            .O(N__16510),
            .I(N__16478));
    InMux I__2661 (
            .O(N__16509),
            .I(N__16475));
    InMux I__2660 (
            .O(N__16508),
            .I(N__16472));
    InMux I__2659 (
            .O(N__16507),
            .I(N__16467));
    InMux I__2658 (
            .O(N__16506),
            .I(N__16467));
    Span4Mux_v I__2657 (
            .O(N__16503),
            .I(N__16458));
    Span4Mux_v I__2656 (
            .O(N__16500),
            .I(N__16458));
    Span4Mux_v I__2655 (
            .O(N__16497),
            .I(N__16458));
    LocalMux I__2654 (
            .O(N__16494),
            .I(N__16458));
    LocalMux I__2653 (
            .O(N__16491),
            .I(N__16453));
    LocalMux I__2652 (
            .O(N__16488),
            .I(N__16453));
    InMux I__2651 (
            .O(N__16487),
            .I(N__16450));
    InMux I__2650 (
            .O(N__16486),
            .I(N__16447));
    Span4Mux_h I__2649 (
            .O(N__16483),
            .I(N__16442));
    LocalMux I__2648 (
            .O(N__16478),
            .I(N__16442));
    LocalMux I__2647 (
            .O(N__16475),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2646 (
            .O(N__16472),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2645 (
            .O(N__16467),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2644 (
            .O(N__16458),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv12 I__2643 (
            .O(N__16453),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2642 (
            .O(N__16450),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2641 (
            .O(N__16447),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2640 (
            .O(N__16442),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__2639 (
            .O(N__16425),
            .I(N__16420));
    InMux I__2638 (
            .O(N__16424),
            .I(N__16413));
    InMux I__2637 (
            .O(N__16423),
            .I(N__16413));
    LocalMux I__2636 (
            .O(N__16420),
            .I(N__16404));
    InMux I__2635 (
            .O(N__16419),
            .I(N__16399));
    InMux I__2634 (
            .O(N__16418),
            .I(N__16399));
    LocalMux I__2633 (
            .O(N__16413),
            .I(N__16396));
    InMux I__2632 (
            .O(N__16412),
            .I(N__16391));
    InMux I__2631 (
            .O(N__16411),
            .I(N__16391));
    InMux I__2630 (
            .O(N__16410),
            .I(N__16388));
    InMux I__2629 (
            .O(N__16409),
            .I(N__16383));
    InMux I__2628 (
            .O(N__16408),
            .I(N__16383));
    InMux I__2627 (
            .O(N__16407),
            .I(N__16380));
    Span4Mux_v I__2626 (
            .O(N__16404),
            .I(N__16371));
    LocalMux I__2625 (
            .O(N__16399),
            .I(N__16371));
    Span4Mux_v I__2624 (
            .O(N__16396),
            .I(N__16371));
    LocalMux I__2623 (
            .O(N__16391),
            .I(N__16371));
    LocalMux I__2622 (
            .O(N__16388),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2621 (
            .O(N__16383),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2620 (
            .O(N__16380),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__2619 (
            .O(N__16371),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    CascadeMux I__2618 (
            .O(N__16362),
            .I(\this_vga_signals.line_clk_1_cascade_ ));
    CascadeMux I__2617 (
            .O(N__16359),
            .I(M_this_vga_signals_line_clk_0_cascade_));
    InMux I__2616 (
            .O(N__16356),
            .I(N__16350));
    InMux I__2615 (
            .O(N__16355),
            .I(N__16350));
    LocalMux I__2614 (
            .O(N__16350),
            .I(\this_vga_signals.un4_lvisibility_1 ));
    InMux I__2613 (
            .O(N__16347),
            .I(N__16343));
    InMux I__2612 (
            .O(N__16346),
            .I(N__16338));
    LocalMux I__2611 (
            .O(N__16343),
            .I(N__16332));
    InMux I__2610 (
            .O(N__16342),
            .I(N__16327));
    InMux I__2609 (
            .O(N__16341),
            .I(N__16327));
    LocalMux I__2608 (
            .O(N__16338),
            .I(N__16324));
    CascadeMux I__2607 (
            .O(N__16337),
            .I(N__16321));
    InMux I__2606 (
            .O(N__16336),
            .I(N__16316));
    InMux I__2605 (
            .O(N__16335),
            .I(N__16313));
    Span4Mux_v I__2604 (
            .O(N__16332),
            .I(N__16306));
    LocalMux I__2603 (
            .O(N__16327),
            .I(N__16306));
    Span4Mux_v I__2602 (
            .O(N__16324),
            .I(N__16306));
    InMux I__2601 (
            .O(N__16321),
            .I(N__16301));
    InMux I__2600 (
            .O(N__16320),
            .I(N__16301));
    InMux I__2599 (
            .O(N__16319),
            .I(N__16298));
    LocalMux I__2598 (
            .O(N__16316),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2597 (
            .O(N__16313),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2596 (
            .O(N__16306),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2595 (
            .O(N__16301),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2594 (
            .O(N__16298),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    CascadeMux I__2593 (
            .O(N__16287),
            .I(N__16284));
    InMux I__2592 (
            .O(N__16284),
            .I(N__16281));
    LocalMux I__2591 (
            .O(N__16281),
            .I(\this_vga_signals.line_clk_1 ));
    InMux I__2590 (
            .O(N__16278),
            .I(N__16275));
    LocalMux I__2589 (
            .O(N__16275),
            .I(N__16263));
    InMux I__2588 (
            .O(N__16274),
            .I(N__16258));
    InMux I__2587 (
            .O(N__16273),
            .I(N__16258));
    InMux I__2586 (
            .O(N__16272),
            .I(N__16255));
    InMux I__2585 (
            .O(N__16271),
            .I(N__16250));
    InMux I__2584 (
            .O(N__16270),
            .I(N__16250));
    InMux I__2583 (
            .O(N__16269),
            .I(N__16245));
    InMux I__2582 (
            .O(N__16268),
            .I(N__16245));
    InMux I__2581 (
            .O(N__16267),
            .I(N__16242));
    InMux I__2580 (
            .O(N__16266),
            .I(N__16239));
    Span4Mux_v I__2579 (
            .O(N__16263),
            .I(N__16234));
    LocalMux I__2578 (
            .O(N__16258),
            .I(N__16234));
    LocalMux I__2577 (
            .O(N__16255),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2576 (
            .O(N__16250),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2575 (
            .O(N__16245),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2574 (
            .O(N__16242),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2573 (
            .O(N__16239),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2572 (
            .O(N__16234),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    CascadeMux I__2571 (
            .O(N__16221),
            .I(\this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0Z0Z_2_cascade_ ));
    InMux I__2570 (
            .O(N__16218),
            .I(N__16213));
    InMux I__2569 (
            .O(N__16217),
            .I(N__16208));
    InMux I__2568 (
            .O(N__16216),
            .I(N__16208));
    LocalMux I__2567 (
            .O(N__16213),
            .I(M_this_substate_qZ0));
    LocalMux I__2566 (
            .O(N__16208),
            .I(M_this_substate_qZ0));
    InMux I__2565 (
            .O(N__16203),
            .I(N__16200));
    LocalMux I__2564 (
            .O(N__16200),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    InMux I__2563 (
            .O(N__16197),
            .I(N__16194));
    LocalMux I__2562 (
            .O(N__16194),
            .I(N__16191));
    Span12Mux_s10_h I__2561 (
            .O(N__16191),
            .I(N__16188));
    Odrv12 I__2560 (
            .O(N__16188),
            .I(M_this_map_ram_write_data_3));
    InMux I__2559 (
            .O(N__16185),
            .I(N__16182));
    LocalMux I__2558 (
            .O(N__16182),
            .I(N__16179));
    Odrv12 I__2557 (
            .O(N__16179),
            .I(M_this_map_ram_write_data_2));
    InMux I__2556 (
            .O(N__16176),
            .I(N__16171));
    CascadeMux I__2555 (
            .O(N__16175),
            .I(N__16167));
    InMux I__2554 (
            .O(N__16174),
            .I(N__16164));
    LocalMux I__2553 (
            .O(N__16171),
            .I(N__16161));
    InMux I__2552 (
            .O(N__16170),
            .I(N__16156));
    InMux I__2551 (
            .O(N__16167),
            .I(N__16156));
    LocalMux I__2550 (
            .O(N__16164),
            .I(N__16152));
    Span4Mux_v I__2549 (
            .O(N__16161),
            .I(N__16148));
    LocalMux I__2548 (
            .O(N__16156),
            .I(N__16145));
    InMux I__2547 (
            .O(N__16155),
            .I(N__16142));
    Span4Mux_h I__2546 (
            .O(N__16152),
            .I(N__16138));
    InMux I__2545 (
            .O(N__16151),
            .I(N__16135));
    Sp12to4 I__2544 (
            .O(N__16148),
            .I(N__16128));
    Sp12to4 I__2543 (
            .O(N__16145),
            .I(N__16128));
    LocalMux I__2542 (
            .O(N__16142),
            .I(N__16128));
    InMux I__2541 (
            .O(N__16141),
            .I(N__16125));
    Odrv4 I__2540 (
            .O(N__16138),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2539 (
            .O(N__16135),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv12 I__2538 (
            .O(N__16128),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2537 (
            .O(N__16125),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    InMux I__2536 (
            .O(N__16116),
            .I(N__16112));
    InMux I__2535 (
            .O(N__16115),
            .I(N__16109));
    LocalMux I__2534 (
            .O(N__16112),
            .I(N__16106));
    LocalMux I__2533 (
            .O(N__16109),
            .I(N__16100));
    Span4Mux_h I__2532 (
            .O(N__16106),
            .I(N__16100));
    InMux I__2531 (
            .O(N__16105),
            .I(N__16097));
    Odrv4 I__2530 (
            .O(N__16100),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__2529 (
            .O(N__16097),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    CascadeMux I__2528 (
            .O(N__16092),
            .I(N__16086));
    CascadeMux I__2527 (
            .O(N__16091),
            .I(N__16080));
    CascadeMux I__2526 (
            .O(N__16090),
            .I(N__16075));
    InMux I__2525 (
            .O(N__16089),
            .I(N__16072));
    InMux I__2524 (
            .O(N__16086),
            .I(N__16068));
    InMux I__2523 (
            .O(N__16085),
            .I(N__16063));
    InMux I__2522 (
            .O(N__16084),
            .I(N__16063));
    InMux I__2521 (
            .O(N__16083),
            .I(N__16058));
    InMux I__2520 (
            .O(N__16080),
            .I(N__16058));
    InMux I__2519 (
            .O(N__16079),
            .I(N__16055));
    InMux I__2518 (
            .O(N__16078),
            .I(N__16052));
    InMux I__2517 (
            .O(N__16075),
            .I(N__16049));
    LocalMux I__2516 (
            .O(N__16072),
            .I(N__16044));
    InMux I__2515 (
            .O(N__16071),
            .I(N__16041));
    LocalMux I__2514 (
            .O(N__16068),
            .I(N__16036));
    LocalMux I__2513 (
            .O(N__16063),
            .I(N__16036));
    LocalMux I__2512 (
            .O(N__16058),
            .I(N__16027));
    LocalMux I__2511 (
            .O(N__16055),
            .I(N__16027));
    LocalMux I__2510 (
            .O(N__16052),
            .I(N__16027));
    LocalMux I__2509 (
            .O(N__16049),
            .I(N__16027));
    CascadeMux I__2508 (
            .O(N__16048),
            .I(N__16024));
    InMux I__2507 (
            .O(N__16047),
            .I(N__16021));
    Span4Mux_h I__2506 (
            .O(N__16044),
            .I(N__16018));
    LocalMux I__2505 (
            .O(N__16041),
            .I(N__16011));
    Span4Mux_h I__2504 (
            .O(N__16036),
            .I(N__16011));
    Span4Mux_v I__2503 (
            .O(N__16027),
            .I(N__16011));
    InMux I__2502 (
            .O(N__16024),
            .I(N__16008));
    LocalMux I__2501 (
            .O(N__16021),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2500 (
            .O(N__16018),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2499 (
            .O(N__16011),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__2498 (
            .O(N__16008),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    CascadeMux I__2497 (
            .O(N__15999),
            .I(N__15995));
    InMux I__2496 (
            .O(N__15998),
            .I(N__15976));
    InMux I__2495 (
            .O(N__15995),
            .I(N__15971));
    InMux I__2494 (
            .O(N__15994),
            .I(N__15971));
    InMux I__2493 (
            .O(N__15993),
            .I(N__15968));
    InMux I__2492 (
            .O(N__15992),
            .I(N__15965));
    InMux I__2491 (
            .O(N__15991),
            .I(N__15962));
    InMux I__2490 (
            .O(N__15990),
            .I(N__15953));
    InMux I__2489 (
            .O(N__15989),
            .I(N__15953));
    InMux I__2488 (
            .O(N__15988),
            .I(N__15953));
    InMux I__2487 (
            .O(N__15987),
            .I(N__15953));
    InMux I__2486 (
            .O(N__15986),
            .I(N__15950));
    InMux I__2485 (
            .O(N__15985),
            .I(N__15947));
    InMux I__2484 (
            .O(N__15984),
            .I(N__15942));
    InMux I__2483 (
            .O(N__15983),
            .I(N__15942));
    InMux I__2482 (
            .O(N__15982),
            .I(N__15936));
    InMux I__2481 (
            .O(N__15981),
            .I(N__15936));
    InMux I__2480 (
            .O(N__15980),
            .I(N__15931));
    InMux I__2479 (
            .O(N__15979),
            .I(N__15931));
    LocalMux I__2478 (
            .O(N__15976),
            .I(N__15926));
    LocalMux I__2477 (
            .O(N__15971),
            .I(N__15926));
    LocalMux I__2476 (
            .O(N__15968),
            .I(N__15915));
    LocalMux I__2475 (
            .O(N__15965),
            .I(N__15915));
    LocalMux I__2474 (
            .O(N__15962),
            .I(N__15915));
    LocalMux I__2473 (
            .O(N__15953),
            .I(N__15915));
    LocalMux I__2472 (
            .O(N__15950),
            .I(N__15915));
    LocalMux I__2471 (
            .O(N__15947),
            .I(N__15910));
    LocalMux I__2470 (
            .O(N__15942),
            .I(N__15910));
    InMux I__2469 (
            .O(N__15941),
            .I(N__15906));
    LocalMux I__2468 (
            .O(N__15936),
            .I(N__15903));
    LocalMux I__2467 (
            .O(N__15931),
            .I(N__15896));
    Span4Mux_v I__2466 (
            .O(N__15926),
            .I(N__15896));
    Span4Mux_v I__2465 (
            .O(N__15915),
            .I(N__15896));
    Span4Mux_h I__2464 (
            .O(N__15910),
            .I(N__15893));
    InMux I__2463 (
            .O(N__15909),
            .I(N__15890));
    LocalMux I__2462 (
            .O(N__15906),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv12 I__2461 (
            .O(N__15903),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2460 (
            .O(N__15896),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2459 (
            .O(N__15893),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2458 (
            .O(N__15890),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    InMux I__2457 (
            .O(N__15879),
            .I(N__15874));
    InMux I__2456 (
            .O(N__15878),
            .I(N__15869));
    InMux I__2455 (
            .O(N__15877),
            .I(N__15869));
    LocalMux I__2454 (
            .O(N__15874),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    LocalMux I__2453 (
            .O(N__15869),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    CascadeMux I__2452 (
            .O(N__15864),
            .I(N__15861));
    InMux I__2451 (
            .O(N__15861),
            .I(N__15856));
    InMux I__2450 (
            .O(N__15860),
            .I(N__15853));
    InMux I__2449 (
            .O(N__15859),
            .I(N__15850));
    LocalMux I__2448 (
            .O(N__15856),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    LocalMux I__2447 (
            .O(N__15853),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    LocalMux I__2446 (
            .O(N__15850),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    CascadeMux I__2445 (
            .O(N__15843),
            .I(N__15838));
    InMux I__2444 (
            .O(N__15842),
            .I(N__15835));
    InMux I__2443 (
            .O(N__15841),
            .I(N__15830));
    InMux I__2442 (
            .O(N__15838),
            .I(N__15830));
    LocalMux I__2441 (
            .O(N__15835),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    LocalMux I__2440 (
            .O(N__15830),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    CascadeMux I__2439 (
            .O(N__15825),
            .I(N__15821));
    InMux I__2438 (
            .O(N__15824),
            .I(N__15817));
    InMux I__2437 (
            .O(N__15821),
            .I(N__15814));
    InMux I__2436 (
            .O(N__15820),
            .I(N__15811));
    LocalMux I__2435 (
            .O(N__15817),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    LocalMux I__2434 (
            .O(N__15814),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    LocalMux I__2433 (
            .O(N__15811),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    InMux I__2432 (
            .O(N__15804),
            .I(N__15799));
    InMux I__2431 (
            .O(N__15803),
            .I(N__15794));
    InMux I__2430 (
            .O(N__15802),
            .I(N__15794));
    LocalMux I__2429 (
            .O(N__15799),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    LocalMux I__2428 (
            .O(N__15794),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    CascadeMux I__2427 (
            .O(N__15789),
            .I(\this_ppu.M_count_d_1_sqmuxa_1_i_a2_4_cascade_ ));
    InMux I__2426 (
            .O(N__15786),
            .I(N__15783));
    LocalMux I__2425 (
            .O(N__15783),
            .I(\this_ppu.M_count_d_1_sqmuxa_1_i_a2_3 ));
    CascadeMux I__2424 (
            .O(N__15780),
            .I(N__15776));
    CascadeMux I__2423 (
            .O(N__15779),
            .I(N__15773));
    InMux I__2422 (
            .O(N__15776),
            .I(N__15758));
    InMux I__2421 (
            .O(N__15773),
            .I(N__15758));
    InMux I__2420 (
            .O(N__15772),
            .I(N__15758));
    InMux I__2419 (
            .O(N__15771),
            .I(N__15758));
    InMux I__2418 (
            .O(N__15770),
            .I(N__15758));
    InMux I__2417 (
            .O(N__15769),
            .I(N__15755));
    LocalMux I__2416 (
            .O(N__15758),
            .I(\this_ppu.un16_0 ));
    LocalMux I__2415 (
            .O(N__15755),
            .I(\this_ppu.un16_0 ));
    CascadeMux I__2414 (
            .O(N__15750),
            .I(N__15747));
    InMux I__2413 (
            .O(N__15747),
            .I(N__15744));
    LocalMux I__2412 (
            .O(N__15744),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ));
    InMux I__2411 (
            .O(N__15741),
            .I(N__15726));
    InMux I__2410 (
            .O(N__15740),
            .I(N__15726));
    InMux I__2409 (
            .O(N__15739),
            .I(N__15726));
    InMux I__2408 (
            .O(N__15738),
            .I(N__15726));
    InMux I__2407 (
            .O(N__15737),
            .I(N__15726));
    LocalMux I__2406 (
            .O(N__15726),
            .I(\this_ppu.N_1195_0 ));
    InMux I__2405 (
            .O(N__15723),
            .I(N__15719));
    CascadeMux I__2404 (
            .O(N__15722),
            .I(N__15716));
    LocalMux I__2403 (
            .O(N__15719),
            .I(N__15712));
    InMux I__2402 (
            .O(N__15716),
            .I(N__15709));
    InMux I__2401 (
            .O(N__15715),
            .I(N__15706));
    Odrv4 I__2400 (
            .O(N__15712),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    LocalMux I__2399 (
            .O(N__15709),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    LocalMux I__2398 (
            .O(N__15706),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    InMux I__2397 (
            .O(N__15699),
            .I(N__15696));
    LocalMux I__2396 (
            .O(N__15696),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_7 ));
    CascadeMux I__2395 (
            .O(N__15693),
            .I(N__15690));
    InMux I__2394 (
            .O(N__15690),
            .I(N__15687));
    LocalMux I__2393 (
            .O(N__15687),
            .I(N__15683));
    InMux I__2392 (
            .O(N__15686),
            .I(N__15680));
    Odrv4 I__2391 (
            .O(N__15683),
            .I(\this_ppu.M_count_qZ0Z_7 ));
    LocalMux I__2390 (
            .O(N__15680),
            .I(\this_ppu.M_count_qZ0Z_7 ));
    CascadeMux I__2389 (
            .O(N__15675),
            .I(\this_vga_signals.N_85_cascade_ ));
    InMux I__2388 (
            .O(N__15672),
            .I(N__15669));
    LocalMux I__2387 (
            .O(N__15669),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_5 ));
    CascadeMux I__2386 (
            .O(N__15666),
            .I(\this_ppu.N_1195_0_cascade_ ));
    InMux I__2385 (
            .O(N__15663),
            .I(N__15660));
    LocalMux I__2384 (
            .O(N__15660),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ));
    InMux I__2383 (
            .O(N__15657),
            .I(N__15653));
    InMux I__2382 (
            .O(N__15656),
            .I(N__15650));
    LocalMux I__2381 (
            .O(N__15653),
            .I(\this_ppu.N_1195_0_1 ));
    LocalMux I__2380 (
            .O(N__15650),
            .I(\this_ppu.N_1195_0_1 ));
    InMux I__2379 (
            .O(N__15645),
            .I(N__15640));
    InMux I__2378 (
            .O(N__15644),
            .I(N__15637));
    InMux I__2377 (
            .O(N__15643),
            .I(N__15634));
    LocalMux I__2376 (
            .O(N__15640),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    LocalMux I__2375 (
            .O(N__15637),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    LocalMux I__2374 (
            .O(N__15634),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    CascadeMux I__2373 (
            .O(N__15627),
            .I(N__15624));
    InMux I__2372 (
            .O(N__15624),
            .I(N__15621));
    LocalMux I__2371 (
            .O(N__15621),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ));
    InMux I__2370 (
            .O(N__15618),
            .I(N__15615));
    LocalMux I__2369 (
            .O(N__15615),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ));
    InMux I__2368 (
            .O(N__15612),
            .I(N__15609));
    LocalMux I__2367 (
            .O(N__15609),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ));
    InMux I__2366 (
            .O(N__15606),
            .I(N__15603));
    LocalMux I__2365 (
            .O(N__15603),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ));
    InMux I__2364 (
            .O(N__15600),
            .I(N__15595));
    InMux I__2363 (
            .O(N__15599),
            .I(N__15592));
    InMux I__2362 (
            .O(N__15598),
            .I(N__15589));
    LocalMux I__2361 (
            .O(N__15595),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    LocalMux I__2360 (
            .O(N__15592),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    LocalMux I__2359 (
            .O(N__15589),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    InMux I__2358 (
            .O(N__15582),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__2357 (
            .O(N__15579),
            .I(N__15573));
    InMux I__2356 (
            .O(N__15578),
            .I(N__15573));
    LocalMux I__2355 (
            .O(N__15573),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    InMux I__2354 (
            .O(N__15570),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__2353 (
            .O(N__15567),
            .I(N__15562));
    InMux I__2352 (
            .O(N__15566),
            .I(N__15557));
    InMux I__2351 (
            .O(N__15565),
            .I(N__15557));
    LocalMux I__2350 (
            .O(N__15562),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    LocalMux I__2349 (
            .O(N__15557),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    InMux I__2348 (
            .O(N__15552),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__2347 (
            .O(N__15549),
            .I(N__15544));
    InMux I__2346 (
            .O(N__15548),
            .I(N__15539));
    InMux I__2345 (
            .O(N__15547),
            .I(N__15539));
    LocalMux I__2344 (
            .O(N__15544),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    LocalMux I__2343 (
            .O(N__15539),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    InMux I__2342 (
            .O(N__15534),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__2341 (
            .O(N__15531),
            .I(bfn_15_10_0_));
    InMux I__2340 (
            .O(N__15528),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    InMux I__2339 (
            .O(N__15525),
            .I(N__15521));
    InMux I__2338 (
            .O(N__15524),
            .I(N__15518));
    LocalMux I__2337 (
            .O(N__15521),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__2336 (
            .O(N__15518),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    CEMux I__2335 (
            .O(N__15513),
            .I(N__15510));
    LocalMux I__2334 (
            .O(N__15510),
            .I(N__15506));
    CEMux I__2333 (
            .O(N__15509),
            .I(N__15501));
    Span4Mux_v I__2332 (
            .O(N__15506),
            .I(N__15498));
    CEMux I__2331 (
            .O(N__15505),
            .I(N__15495));
    CEMux I__2330 (
            .O(N__15504),
            .I(N__15492));
    LocalMux I__2329 (
            .O(N__15501),
            .I(N__15483));
    Span4Mux_v I__2328 (
            .O(N__15498),
            .I(N__15483));
    LocalMux I__2327 (
            .O(N__15495),
            .I(N__15483));
    LocalMux I__2326 (
            .O(N__15492),
            .I(N__15483));
    Odrv4 I__2325 (
            .O(N__15483),
            .I(\this_vga_signals.N_852_0 ));
    InMux I__2324 (
            .O(N__15480),
            .I(N__15477));
    LocalMux I__2323 (
            .O(N__15477),
            .I(N__15469));
    SRMux I__2322 (
            .O(N__15476),
            .I(N__15456));
    SRMux I__2321 (
            .O(N__15475),
            .I(N__15456));
    SRMux I__2320 (
            .O(N__15474),
            .I(N__15456));
    SRMux I__2319 (
            .O(N__15473),
            .I(N__15456));
    SRMux I__2318 (
            .O(N__15472),
            .I(N__15456));
    Glb2LocalMux I__2317 (
            .O(N__15469),
            .I(N__15456));
    GlobalMux I__2316 (
            .O(N__15456),
            .I(N__15453));
    gio2CtrlBuf I__2315 (
            .O(N__15453),
            .I(\this_vga_signals.N_1098_g ));
    InMux I__2314 (
            .O(N__15450),
            .I(N__15447));
    LocalMux I__2313 (
            .O(N__15447),
            .I(N__15444));
    Span12Mux_v I__2312 (
            .O(N__15444),
            .I(N__15441));
    Span12Mux_h I__2311 (
            .O(N__15441),
            .I(N__15438));
    Odrv12 I__2310 (
            .O(N__15438),
            .I(port_clk_c));
    InMux I__2309 (
            .O(N__15435),
            .I(N__15432));
    LocalMux I__2308 (
            .O(N__15432),
            .I(N__15429));
    Odrv4 I__2307 (
            .O(N__15429),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    InMux I__2306 (
            .O(N__15426),
            .I(N__15423));
    LocalMux I__2305 (
            .O(N__15423),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    InMux I__2304 (
            .O(N__15420),
            .I(N__15417));
    LocalMux I__2303 (
            .O(N__15417),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    InMux I__2302 (
            .O(N__15414),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__2301 (
            .O(N__15411),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__2300 (
            .O(N__15408),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__2299 (
            .O(N__15405),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1 ));
    InMux I__2298 (
            .O(N__15402),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1 ));
    InMux I__2297 (
            .O(N__15399),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1 ));
    InMux I__2296 (
            .O(N__15396),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1 ));
    InMux I__2295 (
            .O(N__15393),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1 ));
    InMux I__2294 (
            .O(N__15390),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1 ));
    InMux I__2293 (
            .O(N__15387),
            .I(\this_ppu.un1_M_count_q_1_cry_6_s1 ));
    InMux I__2292 (
            .O(N__15384),
            .I(N__15381));
    LocalMux I__2291 (
            .O(N__15381),
            .I(N__15378));
    Odrv4 I__2290 (
            .O(N__15378),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    CascadeMux I__2289 (
            .O(N__15375),
            .I(N__15372));
    InMux I__2288 (
            .O(N__15372),
            .I(N__15367));
    CascadeMux I__2287 (
            .O(N__15371),
            .I(N__15361));
    CascadeMux I__2286 (
            .O(N__15370),
            .I(N__15358));
    LocalMux I__2285 (
            .O(N__15367),
            .I(N__15355));
    InMux I__2284 (
            .O(N__15366),
            .I(N__15350));
    InMux I__2283 (
            .O(N__15365),
            .I(N__15350));
    InMux I__2282 (
            .O(N__15364),
            .I(N__15343));
    InMux I__2281 (
            .O(N__15361),
            .I(N__15343));
    InMux I__2280 (
            .O(N__15358),
            .I(N__15343));
    Odrv4 I__2279 (
            .O(N__15355),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__2278 (
            .O(N__15350),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__2277 (
            .O(N__15343),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    CascadeMux I__2276 (
            .O(N__15336),
            .I(\this_vga_signals.un6_vvisibilitylto8_0_cascade_ ));
    CascadeMux I__2275 (
            .O(N__15333),
            .I(\this_vga_signals.un6_vvisibilitylt9_0_cascade_ ));
    CascadeMux I__2274 (
            .O(N__15330),
            .I(this_vga_signals_vvisibility_1_cascade_));
    InMux I__2273 (
            .O(N__15327),
            .I(N__15322));
    InMux I__2272 (
            .O(N__15326),
            .I(N__15319));
    CascadeMux I__2271 (
            .O(N__15325),
            .I(N__15316));
    LocalMux I__2270 (
            .O(N__15322),
            .I(N__15313));
    LocalMux I__2269 (
            .O(N__15319),
            .I(N__15310));
    InMux I__2268 (
            .O(N__15316),
            .I(N__15307));
    Sp12to4 I__2267 (
            .O(N__15313),
            .I(N__15304));
    Span4Mux_v I__2266 (
            .O(N__15310),
            .I(N__15299));
    LocalMux I__2265 (
            .O(N__15307),
            .I(N__15299));
    Span12Mux_s9_v I__2264 (
            .O(N__15304),
            .I(N__15296));
    Span4Mux_h I__2263 (
            .O(N__15299),
            .I(N__15293));
    Span12Mux_v I__2262 (
            .O(N__15296),
            .I(N__15290));
    Span4Mux_h I__2261 (
            .O(N__15293),
            .I(N__15287));
    Odrv12 I__2260 (
            .O(N__15290),
            .I(\this_vga_signals.vvisibility ));
    Odrv4 I__2259 (
            .O(N__15287),
            .I(\this_vga_signals.vvisibility ));
    InMux I__2258 (
            .O(N__15282),
            .I(N__15279));
    LocalMux I__2257 (
            .O(N__15279),
            .I(\this_vga_signals.vaddress_ac0_9_0_a0_0 ));
    CascadeMux I__2256 (
            .O(N__15276),
            .I(\this_ppu.N_1195_0_1_cascade_ ));
    CascadeMux I__2255 (
            .O(N__15273),
            .I(N__15269));
    InMux I__2254 (
            .O(N__15272),
            .I(N__15264));
    InMux I__2253 (
            .O(N__15269),
            .I(N__15264));
    LocalMux I__2252 (
            .O(N__15264),
            .I(N__15260));
    InMux I__2251 (
            .O(N__15263),
            .I(N__15257));
    Odrv4 I__2250 (
            .O(N__15260),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    LocalMux I__2249 (
            .O(N__15257),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    InMux I__2248 (
            .O(N__15252),
            .I(N__15249));
    LocalMux I__2247 (
            .O(N__15249),
            .I(N__15246));
    Span4Mux_h I__2246 (
            .O(N__15246),
            .I(N__15242));
    InMux I__2245 (
            .O(N__15245),
            .I(N__15239));
    Odrv4 I__2244 (
            .O(N__15242),
            .I(\this_vga_signals.vaddress_c3_0 ));
    LocalMux I__2243 (
            .O(N__15239),
            .I(\this_vga_signals.vaddress_c3_0 ));
    InMux I__2242 (
            .O(N__15234),
            .I(N__15229));
    InMux I__2241 (
            .O(N__15233),
            .I(N__15224));
    InMux I__2240 (
            .O(N__15232),
            .I(N__15224));
    LocalMux I__2239 (
            .O(N__15229),
            .I(N__15220));
    LocalMux I__2238 (
            .O(N__15224),
            .I(N__15217));
    InMux I__2237 (
            .O(N__15223),
            .I(N__15213));
    Span4Mux_h I__2236 (
            .O(N__15220),
            .I(N__15209));
    Span4Mux_h I__2235 (
            .O(N__15217),
            .I(N__15206));
    InMux I__2234 (
            .O(N__15216),
            .I(N__15203));
    LocalMux I__2233 (
            .O(N__15213),
            .I(N__15200));
    InMux I__2232 (
            .O(N__15212),
            .I(N__15197));
    Odrv4 I__2231 (
            .O(N__15209),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__2230 (
            .O(N__15206),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__2229 (
            .O(N__15203),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__2228 (
            .O(N__15200),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__2227 (
            .O(N__15197),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    CascadeMux I__2226 (
            .O(N__15186),
            .I(N__15183));
    InMux I__2225 (
            .O(N__15183),
            .I(N__15179));
    InMux I__2224 (
            .O(N__15182),
            .I(N__15174));
    LocalMux I__2223 (
            .O(N__15179),
            .I(N__15171));
    InMux I__2222 (
            .O(N__15178),
            .I(N__15166));
    InMux I__2221 (
            .O(N__15177),
            .I(N__15166));
    LocalMux I__2220 (
            .O(N__15174),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv4 I__2219 (
            .O(N__15171),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__2218 (
            .O(N__15166),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    InMux I__2217 (
            .O(N__15159),
            .I(N__15156));
    LocalMux I__2216 (
            .O(N__15156),
            .I(N__15153));
    Span4Mux_h I__2215 (
            .O(N__15153),
            .I(N__15150));
    Odrv4 I__2214 (
            .O(N__15150),
            .I(\this_vga_signals.if_m8_0_a3_1_1_1 ));
    CascadeMux I__2213 (
            .O(N__15147),
            .I(N__15143));
    CascadeMux I__2212 (
            .O(N__15146),
            .I(N__15138));
    InMux I__2211 (
            .O(N__15143),
            .I(N__15135));
    InMux I__2210 (
            .O(N__15142),
            .I(N__15132));
    InMux I__2209 (
            .O(N__15141),
            .I(N__15127));
    InMux I__2208 (
            .O(N__15138),
            .I(N__15127));
    LocalMux I__2207 (
            .O(N__15135),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__2206 (
            .O(N__15132),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__2205 (
            .O(N__15127),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    InMux I__2204 (
            .O(N__15120),
            .I(N__15117));
    LocalMux I__2203 (
            .O(N__15117),
            .I(\this_vga_signals.g2 ));
    InMux I__2202 (
            .O(N__15114),
            .I(N__15111));
    LocalMux I__2201 (
            .O(N__15111),
            .I(N__15107));
    CascadeMux I__2200 (
            .O(N__15110),
            .I(N__15101));
    Span4Mux_h I__2199 (
            .O(N__15107),
            .I(N__15096));
    InMux I__2198 (
            .O(N__15106),
            .I(N__15093));
    InMux I__2197 (
            .O(N__15105),
            .I(N__15088));
    InMux I__2196 (
            .O(N__15104),
            .I(N__15088));
    InMux I__2195 (
            .O(N__15101),
            .I(N__15085));
    InMux I__2194 (
            .O(N__15100),
            .I(N__15080));
    InMux I__2193 (
            .O(N__15099),
            .I(N__15080));
    Odrv4 I__2192 (
            .O(N__15096),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2191 (
            .O(N__15093),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2190 (
            .O(N__15088),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2189 (
            .O(N__15085),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2188 (
            .O(N__15080),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    CascadeMux I__2187 (
            .O(N__15069),
            .I(N__15066));
    InMux I__2186 (
            .O(N__15066),
            .I(N__15063));
    LocalMux I__2185 (
            .O(N__15063),
            .I(\this_vga_signals.g1_3 ));
    CascadeMux I__2184 (
            .O(N__15060),
            .I(N__15057));
    InMux I__2183 (
            .O(N__15057),
            .I(N__15054));
    LocalMux I__2182 (
            .O(N__15054),
            .I(N__15051));
    Span4Mux_h I__2181 (
            .O(N__15051),
            .I(N__15044));
    InMux I__2180 (
            .O(N__15050),
            .I(N__15041));
    InMux I__2179 (
            .O(N__15049),
            .I(N__15038));
    InMux I__2178 (
            .O(N__15048),
            .I(N__15033));
    InMux I__2177 (
            .O(N__15047),
            .I(N__15033));
    Odrv4 I__2176 (
            .O(N__15044),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__2175 (
            .O(N__15041),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__2174 (
            .O(N__15038),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__2173 (
            .O(N__15033),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__2172 (
            .O(N__15024),
            .I(N__15020));
    CascadeMux I__2171 (
            .O(N__15023),
            .I(N__15013));
    LocalMux I__2170 (
            .O(N__15020),
            .I(N__15010));
    InMux I__2169 (
            .O(N__15019),
            .I(N__15005));
    InMux I__2168 (
            .O(N__15018),
            .I(N__15000));
    InMux I__2167 (
            .O(N__15017),
            .I(N__15000));
    InMux I__2166 (
            .O(N__15016),
            .I(N__14997));
    InMux I__2165 (
            .O(N__15013),
            .I(N__14994));
    Span4Mux_h I__2164 (
            .O(N__15010),
            .I(N__14991));
    InMux I__2163 (
            .O(N__15009),
            .I(N__14988));
    InMux I__2162 (
            .O(N__15008),
            .I(N__14985));
    LocalMux I__2161 (
            .O(N__15005),
            .I(N__14980));
    LocalMux I__2160 (
            .O(N__15000),
            .I(N__14980));
    LocalMux I__2159 (
            .O(N__14997),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2158 (
            .O(N__14994),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__2157 (
            .O(N__14991),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2156 (
            .O(N__14988),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2155 (
            .O(N__14985),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__2154 (
            .O(N__14980),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    CascadeMux I__2153 (
            .O(N__14967),
            .I(N__14962));
    InMux I__2152 (
            .O(N__14966),
            .I(N__14953));
    InMux I__2151 (
            .O(N__14965),
            .I(N__14946));
    InMux I__2150 (
            .O(N__14962),
            .I(N__14946));
    InMux I__2149 (
            .O(N__14961),
            .I(N__14946));
    InMux I__2148 (
            .O(N__14960),
            .I(N__14943));
    InMux I__2147 (
            .O(N__14959),
            .I(N__14940));
    InMux I__2146 (
            .O(N__14958),
            .I(N__14937));
    InMux I__2145 (
            .O(N__14957),
            .I(N__14934));
    InMux I__2144 (
            .O(N__14956),
            .I(N__14931));
    LocalMux I__2143 (
            .O(N__14953),
            .I(N__14926));
    LocalMux I__2142 (
            .O(N__14946),
            .I(N__14921));
    LocalMux I__2141 (
            .O(N__14943),
            .I(N__14921));
    LocalMux I__2140 (
            .O(N__14940),
            .I(N__14916));
    LocalMux I__2139 (
            .O(N__14937),
            .I(N__14909));
    LocalMux I__2138 (
            .O(N__14934),
            .I(N__14909));
    LocalMux I__2137 (
            .O(N__14931),
            .I(N__14909));
    InMux I__2136 (
            .O(N__14930),
            .I(N__14906));
    InMux I__2135 (
            .O(N__14929),
            .I(N__14902));
    Span4Mux_h I__2134 (
            .O(N__14926),
            .I(N__14897));
    Span4Mux_h I__2133 (
            .O(N__14921),
            .I(N__14897));
    InMux I__2132 (
            .O(N__14920),
            .I(N__14894));
    InMux I__2131 (
            .O(N__14919),
            .I(N__14891));
    Span4Mux_v I__2130 (
            .O(N__14916),
            .I(N__14886));
    Span4Mux_v I__2129 (
            .O(N__14909),
            .I(N__14886));
    LocalMux I__2128 (
            .O(N__14906),
            .I(N__14883));
    InMux I__2127 (
            .O(N__14905),
            .I(N__14880));
    LocalMux I__2126 (
            .O(N__14902),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__2125 (
            .O(N__14897),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2124 (
            .O(N__14894),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2123 (
            .O(N__14891),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__2122 (
            .O(N__14886),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__2121 (
            .O(N__14883),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2120 (
            .O(N__14880),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__2119 (
            .O(N__14865),
            .I(N__14862));
    LocalMux I__2118 (
            .O(N__14862),
            .I(N__14859));
    Span4Mux_h I__2117 (
            .O(N__14859),
            .I(N__14856));
    Odrv4 I__2116 (
            .O(N__14856),
            .I(\this_vga_signals.if_m2 ));
    SRMux I__2115 (
            .O(N__14853),
            .I(N__14850));
    LocalMux I__2114 (
            .O(N__14850),
            .I(N__14845));
    SRMux I__2113 (
            .O(N__14849),
            .I(N__14842));
    SRMux I__2112 (
            .O(N__14848),
            .I(N__14839));
    Span4Mux_h I__2111 (
            .O(N__14845),
            .I(N__14835));
    LocalMux I__2110 (
            .O(N__14842),
            .I(N__14832));
    LocalMux I__2109 (
            .O(N__14839),
            .I(N__14829));
    InMux I__2108 (
            .O(N__14838),
            .I(N__14826));
    Odrv4 I__2107 (
            .O(N__14835),
            .I(\this_vga_signals.N_1098_1 ));
    Odrv4 I__2106 (
            .O(N__14832),
            .I(\this_vga_signals.N_1098_1 ));
    Odrv4 I__2105 (
            .O(N__14829),
            .I(\this_vga_signals.N_1098_1 ));
    LocalMux I__2104 (
            .O(N__14826),
            .I(\this_vga_signals.N_1098_1 ));
    InMux I__2103 (
            .O(N__14817),
            .I(N__14814));
    LocalMux I__2102 (
            .O(N__14814),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    CascadeMux I__2101 (
            .O(N__14811),
            .I(N__14808));
    InMux I__2100 (
            .O(N__14808),
            .I(N__14802));
    InMux I__2099 (
            .O(N__14807),
            .I(N__14795));
    InMux I__2098 (
            .O(N__14806),
            .I(N__14795));
    InMux I__2097 (
            .O(N__14805),
            .I(N__14795));
    LocalMux I__2096 (
            .O(N__14802),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__2095 (
            .O(N__14795),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    InMux I__2094 (
            .O(N__14790),
            .I(N__14787));
    LocalMux I__2093 (
            .O(N__14787),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_0_N_2L1 ));
    InMux I__2092 (
            .O(N__14784),
            .I(N__14779));
    InMux I__2091 (
            .O(N__14783),
            .I(N__14774));
    InMux I__2090 (
            .O(N__14782),
            .I(N__14774));
    LocalMux I__2089 (
            .O(N__14779),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__2088 (
            .O(N__14774),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    CascadeMux I__2087 (
            .O(N__14769),
            .I(\this_vga_signals.SUM_2_i_1_2_3_cascade_ ));
    InMux I__2086 (
            .O(N__14766),
            .I(N__14762));
    InMux I__2085 (
            .O(N__14765),
            .I(N__14759));
    LocalMux I__2084 (
            .O(N__14762),
            .I(\this_vga_signals.SUM_2_i_1_1_3 ));
    LocalMux I__2083 (
            .O(N__14759),
            .I(\this_vga_signals.SUM_2_i_1_1_3 ));
    CascadeMux I__2082 (
            .O(N__14754),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_x0_cascade_ ));
    CascadeMux I__2081 (
            .O(N__14751),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ));
    InMux I__2080 (
            .O(N__14748),
            .I(N__14741));
    InMux I__2079 (
            .O(N__14747),
            .I(N__14736));
    InMux I__2078 (
            .O(N__14746),
            .I(N__14736));
    CascadeMux I__2077 (
            .O(N__14745),
            .I(N__14733));
    InMux I__2076 (
            .O(N__14744),
            .I(N__14729));
    LocalMux I__2075 (
            .O(N__14741),
            .I(N__14724));
    LocalMux I__2074 (
            .O(N__14736),
            .I(N__14724));
    InMux I__2073 (
            .O(N__14733),
            .I(N__14721));
    InMux I__2072 (
            .O(N__14732),
            .I(N__14718));
    LocalMux I__2071 (
            .O(N__14729),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__2070 (
            .O(N__14724),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__2069 (
            .O(N__14721),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__2068 (
            .O(N__14718),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    CascadeMux I__2067 (
            .O(N__14709),
            .I(N__14704));
    CascadeMux I__2066 (
            .O(N__14708),
            .I(N__14700));
    InMux I__2065 (
            .O(N__14707),
            .I(N__14697));
    InMux I__2064 (
            .O(N__14704),
            .I(N__14694));
    InMux I__2063 (
            .O(N__14703),
            .I(N__14689));
    InMux I__2062 (
            .O(N__14700),
            .I(N__14689));
    LocalMux I__2061 (
            .O(N__14697),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__2060 (
            .O(N__14694),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__2059 (
            .O(N__14689),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    CascadeMux I__2058 (
            .O(N__14682),
            .I(N__14679));
    InMux I__2057 (
            .O(N__14679),
            .I(N__14673));
    InMux I__2056 (
            .O(N__14678),
            .I(N__14673));
    LocalMux I__2055 (
            .O(N__14673),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_N_2L1 ));
    InMux I__2054 (
            .O(N__14670),
            .I(N__14667));
    LocalMux I__2053 (
            .O(N__14667),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_x1 ));
    InMux I__2052 (
            .O(N__14664),
            .I(N__14655));
    InMux I__2051 (
            .O(N__14663),
            .I(N__14650));
    InMux I__2050 (
            .O(N__14662),
            .I(N__14650));
    InMux I__2049 (
            .O(N__14661),
            .I(N__14647));
    InMux I__2048 (
            .O(N__14660),
            .I(N__14640));
    InMux I__2047 (
            .O(N__14659),
            .I(N__14640));
    InMux I__2046 (
            .O(N__14658),
            .I(N__14640));
    LocalMux I__2045 (
            .O(N__14655),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__2044 (
            .O(N__14650),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__2043 (
            .O(N__14647),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__2042 (
            .O(N__14640),
            .I(\this_vga_signals.vaddress_5 ));
    InMux I__2041 (
            .O(N__14631),
            .I(N__14628));
    LocalMux I__2040 (
            .O(N__14628),
            .I(N__14625));
    Odrv4 I__2039 (
            .O(N__14625),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_0 ));
    InMux I__2038 (
            .O(N__14622),
            .I(N__14614));
    InMux I__2037 (
            .O(N__14621),
            .I(N__14611));
    InMux I__2036 (
            .O(N__14620),
            .I(N__14607));
    InMux I__2035 (
            .O(N__14619),
            .I(N__14604));
    InMux I__2034 (
            .O(N__14618),
            .I(N__14599));
    InMux I__2033 (
            .O(N__14617),
            .I(N__14599));
    LocalMux I__2032 (
            .O(N__14614),
            .I(N__14594));
    LocalMux I__2031 (
            .O(N__14611),
            .I(N__14594));
    InMux I__2030 (
            .O(N__14610),
            .I(N__14591));
    LocalMux I__2029 (
            .O(N__14607),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__2028 (
            .O(N__14604),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__2027 (
            .O(N__14599),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    Odrv4 I__2026 (
            .O(N__14594),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__2025 (
            .O(N__14591),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    InMux I__2024 (
            .O(N__14580),
            .I(N__14573));
    InMux I__2023 (
            .O(N__14579),
            .I(N__14573));
    InMux I__2022 (
            .O(N__14578),
            .I(N__14565));
    LocalMux I__2021 (
            .O(N__14573),
            .I(N__14562));
    InMux I__2020 (
            .O(N__14572),
            .I(N__14555));
    InMux I__2019 (
            .O(N__14571),
            .I(N__14555));
    InMux I__2018 (
            .O(N__14570),
            .I(N__14555));
    InMux I__2017 (
            .O(N__14569),
            .I(N__14550));
    InMux I__2016 (
            .O(N__14568),
            .I(N__14550));
    LocalMux I__2015 (
            .O(N__14565),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__2014 (
            .O(N__14562),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__2013 (
            .O(N__14555),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__2012 (
            .O(N__14550),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    CascadeMux I__2011 (
            .O(N__14541),
            .I(\this_vga_signals.g2_0_a2_5Z0Z_1_cascade_ ));
    InMux I__2010 (
            .O(N__14538),
            .I(N__14535));
    LocalMux I__2009 (
            .O(N__14535),
            .I(\this_vga_signals.g2_0_a2_2 ));
    InMux I__2008 (
            .O(N__14532),
            .I(N__14529));
    LocalMux I__2007 (
            .O(N__14529),
            .I(N__14526));
    Span4Mux_h I__2006 (
            .O(N__14526),
            .I(N__14523));
    Odrv4 I__2005 (
            .O(N__14523),
            .I(\this_vga_signals.g2_0_a2_5 ));
    CEMux I__2004 (
            .O(N__14520),
            .I(N__14517));
    LocalMux I__2003 (
            .O(N__14517),
            .I(N__14514));
    Odrv4 I__2002 (
            .O(N__14514),
            .I(\this_vga_signals.N_852_1 ));
    InMux I__2001 (
            .O(N__14511),
            .I(N__14508));
    LocalMux I__2000 (
            .O(N__14508),
            .I(N__14502));
    InMux I__1999 (
            .O(N__14507),
            .I(N__14495));
    InMux I__1998 (
            .O(N__14506),
            .I(N__14495));
    InMux I__1997 (
            .O(N__14505),
            .I(N__14492));
    Span12Mux_s11_h I__1996 (
            .O(N__14502),
            .I(N__14489));
    InMux I__1995 (
            .O(N__14501),
            .I(N__14484));
    InMux I__1994 (
            .O(N__14500),
            .I(N__14484));
    LocalMux I__1993 (
            .O(N__14495),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1992 (
            .O(N__14492),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv12 I__1991 (
            .O(N__14489),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1990 (
            .O(N__14484),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    InMux I__1989 (
            .O(N__14475),
            .I(N__14472));
    LocalMux I__1988 (
            .O(N__14472),
            .I(\this_vga_signals.un2_hsynclt6_0 ));
    InMux I__1987 (
            .O(N__14469),
            .I(N__14466));
    LocalMux I__1986 (
            .O(N__14466),
            .I(N__14456));
    InMux I__1985 (
            .O(N__14465),
            .I(N__14451));
    InMux I__1984 (
            .O(N__14464),
            .I(N__14451));
    CascadeMux I__1983 (
            .O(N__14463),
            .I(N__14445));
    InMux I__1982 (
            .O(N__14462),
            .I(N__14442));
    InMux I__1981 (
            .O(N__14461),
            .I(N__14439));
    CascadeMux I__1980 (
            .O(N__14460),
            .I(N__14435));
    InMux I__1979 (
            .O(N__14459),
            .I(N__14432));
    Span4Mux_v I__1978 (
            .O(N__14456),
            .I(N__14426));
    LocalMux I__1977 (
            .O(N__14451),
            .I(N__14426));
    InMux I__1976 (
            .O(N__14450),
            .I(N__14423));
    InMux I__1975 (
            .O(N__14449),
            .I(N__14416));
    InMux I__1974 (
            .O(N__14448),
            .I(N__14416));
    InMux I__1973 (
            .O(N__14445),
            .I(N__14416));
    LocalMux I__1972 (
            .O(N__14442),
            .I(N__14413));
    LocalMux I__1971 (
            .O(N__14439),
            .I(N__14396));
    InMux I__1970 (
            .O(N__14438),
            .I(N__14393));
    InMux I__1969 (
            .O(N__14435),
            .I(N__14390));
    LocalMux I__1968 (
            .O(N__14432),
            .I(N__14387));
    InMux I__1967 (
            .O(N__14431),
            .I(N__14384));
    Span4Mux_v I__1966 (
            .O(N__14426),
            .I(N__14379));
    LocalMux I__1965 (
            .O(N__14423),
            .I(N__14379));
    LocalMux I__1964 (
            .O(N__14416),
            .I(N__14374));
    Span4Mux_h I__1963 (
            .O(N__14413),
            .I(N__14374));
    InMux I__1962 (
            .O(N__14412),
            .I(N__14367));
    InMux I__1961 (
            .O(N__14411),
            .I(N__14367));
    InMux I__1960 (
            .O(N__14410),
            .I(N__14367));
    InMux I__1959 (
            .O(N__14409),
            .I(N__14356));
    InMux I__1958 (
            .O(N__14408),
            .I(N__14356));
    InMux I__1957 (
            .O(N__14407),
            .I(N__14356));
    InMux I__1956 (
            .O(N__14406),
            .I(N__14356));
    InMux I__1955 (
            .O(N__14405),
            .I(N__14356));
    InMux I__1954 (
            .O(N__14404),
            .I(N__14343));
    InMux I__1953 (
            .O(N__14403),
            .I(N__14343));
    InMux I__1952 (
            .O(N__14402),
            .I(N__14343));
    InMux I__1951 (
            .O(N__14401),
            .I(N__14343));
    InMux I__1950 (
            .O(N__14400),
            .I(N__14343));
    InMux I__1949 (
            .O(N__14399),
            .I(N__14343));
    Odrv4 I__1948 (
            .O(N__14396),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1947 (
            .O(N__14393),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1946 (
            .O(N__14390),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1945 (
            .O(N__14387),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1944 (
            .O(N__14384),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1943 (
            .O(N__14379),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1942 (
            .O(N__14374),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1941 (
            .O(N__14367),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1940 (
            .O(N__14356),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1939 (
            .O(N__14343),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    InMux I__1938 (
            .O(N__14322),
            .I(N__14319));
    LocalMux I__1937 (
            .O(N__14319),
            .I(N__14316));
    Span4Mux_h I__1936 (
            .O(N__14316),
            .I(N__14313));
    Odrv4 I__1935 (
            .O(N__14313),
            .I(\this_vga_signals.un2_hsynclt7 ));
    InMux I__1934 (
            .O(N__14310),
            .I(N__14306));
    InMux I__1933 (
            .O(N__14309),
            .I(N__14303));
    LocalMux I__1932 (
            .O(N__14306),
            .I(\this_vga_signals.un2_hsynclto3_0 ));
    LocalMux I__1931 (
            .O(N__14303),
            .I(\this_vga_signals.un2_hsynclto3_0 ));
    CascadeMux I__1930 (
            .O(N__14298),
            .I(N__14290));
    CascadeMux I__1929 (
            .O(N__14297),
            .I(N__14285));
    CascadeMux I__1928 (
            .O(N__14296),
            .I(N__14282));
    CascadeMux I__1927 (
            .O(N__14295),
            .I(N__14279));
    InMux I__1926 (
            .O(N__14294),
            .I(N__14271));
    InMux I__1925 (
            .O(N__14293),
            .I(N__14271));
    InMux I__1924 (
            .O(N__14290),
            .I(N__14271));
    CascadeMux I__1923 (
            .O(N__14289),
            .I(N__14267));
    CascadeMux I__1922 (
            .O(N__14288),
            .I(N__14263));
    InMux I__1921 (
            .O(N__14285),
            .I(N__14258));
    InMux I__1920 (
            .O(N__14282),
            .I(N__14255));
    InMux I__1919 (
            .O(N__14279),
            .I(N__14249));
    InMux I__1918 (
            .O(N__14278),
            .I(N__14249));
    LocalMux I__1917 (
            .O(N__14271),
            .I(N__14245));
    InMux I__1916 (
            .O(N__14270),
            .I(N__14242));
    InMux I__1915 (
            .O(N__14267),
            .I(N__14239));
    CascadeMux I__1914 (
            .O(N__14266),
            .I(N__14234));
    InMux I__1913 (
            .O(N__14263),
            .I(N__14229));
    InMux I__1912 (
            .O(N__14262),
            .I(N__14229));
    InMux I__1911 (
            .O(N__14261),
            .I(N__14226));
    LocalMux I__1910 (
            .O(N__14258),
            .I(N__14221));
    LocalMux I__1909 (
            .O(N__14255),
            .I(N__14221));
    CascadeMux I__1908 (
            .O(N__14254),
            .I(N__14212));
    LocalMux I__1907 (
            .O(N__14249),
            .I(N__14206));
    InMux I__1906 (
            .O(N__14248),
            .I(N__14203));
    Span4Mux_v I__1905 (
            .O(N__14245),
            .I(N__14196));
    LocalMux I__1904 (
            .O(N__14242),
            .I(N__14196));
    LocalMux I__1903 (
            .O(N__14239),
            .I(N__14196));
    InMux I__1902 (
            .O(N__14238),
            .I(N__14189));
    InMux I__1901 (
            .O(N__14237),
            .I(N__14189));
    InMux I__1900 (
            .O(N__14234),
            .I(N__14189));
    LocalMux I__1899 (
            .O(N__14229),
            .I(N__14186));
    LocalMux I__1898 (
            .O(N__14226),
            .I(N__14181));
    Span4Mux_h I__1897 (
            .O(N__14221),
            .I(N__14181));
    InMux I__1896 (
            .O(N__14220),
            .I(N__14170));
    InMux I__1895 (
            .O(N__14219),
            .I(N__14170));
    InMux I__1894 (
            .O(N__14218),
            .I(N__14170));
    InMux I__1893 (
            .O(N__14217),
            .I(N__14170));
    InMux I__1892 (
            .O(N__14216),
            .I(N__14170));
    InMux I__1891 (
            .O(N__14215),
            .I(N__14161));
    InMux I__1890 (
            .O(N__14212),
            .I(N__14161));
    InMux I__1889 (
            .O(N__14211),
            .I(N__14161));
    InMux I__1888 (
            .O(N__14210),
            .I(N__14161));
    InMux I__1887 (
            .O(N__14209),
            .I(N__14158));
    Odrv4 I__1886 (
            .O(N__14206),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1885 (
            .O(N__14203),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__1884 (
            .O(N__14196),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1883 (
            .O(N__14189),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__1882 (
            .O(N__14186),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__1881 (
            .O(N__14181),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1880 (
            .O(N__14170),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1879 (
            .O(N__14161),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1878 (
            .O(N__14158),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    CascadeMux I__1877 (
            .O(N__14139),
            .I(N__14134));
    CascadeMux I__1876 (
            .O(N__14138),
            .I(N__14129));
    InMux I__1875 (
            .O(N__14137),
            .I(N__14118));
    InMux I__1874 (
            .O(N__14134),
            .I(N__14118));
    InMux I__1873 (
            .O(N__14133),
            .I(N__14115));
    InMux I__1872 (
            .O(N__14132),
            .I(N__14108));
    InMux I__1871 (
            .O(N__14129),
            .I(N__14108));
    InMux I__1870 (
            .O(N__14128),
            .I(N__14108));
    InMux I__1869 (
            .O(N__14127),
            .I(N__14105));
    InMux I__1868 (
            .O(N__14126),
            .I(N__14100));
    InMux I__1867 (
            .O(N__14125),
            .I(N__14100));
    InMux I__1866 (
            .O(N__14124),
            .I(N__14095));
    InMux I__1865 (
            .O(N__14123),
            .I(N__14095));
    LocalMux I__1864 (
            .O(N__14118),
            .I(N__14091));
    LocalMux I__1863 (
            .O(N__14115),
            .I(N__14083));
    LocalMux I__1862 (
            .O(N__14108),
            .I(N__14080));
    LocalMux I__1861 (
            .O(N__14105),
            .I(N__14073));
    LocalMux I__1860 (
            .O(N__14100),
            .I(N__14073));
    LocalMux I__1859 (
            .O(N__14095),
            .I(N__14073));
    InMux I__1858 (
            .O(N__14094),
            .I(N__14070));
    Span4Mux_v I__1857 (
            .O(N__14091),
            .I(N__14067));
    InMux I__1856 (
            .O(N__14090),
            .I(N__14060));
    InMux I__1855 (
            .O(N__14089),
            .I(N__14060));
    InMux I__1854 (
            .O(N__14088),
            .I(N__14060));
    InMux I__1853 (
            .O(N__14087),
            .I(N__14050));
    InMux I__1852 (
            .O(N__14086),
            .I(N__14047));
    Span4Mux_h I__1851 (
            .O(N__14083),
            .I(N__14042));
    Span4Mux_h I__1850 (
            .O(N__14080),
            .I(N__14042));
    Span4Mux_v I__1849 (
            .O(N__14073),
            .I(N__14039));
    LocalMux I__1848 (
            .O(N__14070),
            .I(N__14036));
    Sp12to4 I__1847 (
            .O(N__14067),
            .I(N__14031));
    LocalMux I__1846 (
            .O(N__14060),
            .I(N__14031));
    InMux I__1845 (
            .O(N__14059),
            .I(N__14026));
    InMux I__1844 (
            .O(N__14058),
            .I(N__14026));
    InMux I__1843 (
            .O(N__14057),
            .I(N__14019));
    InMux I__1842 (
            .O(N__14056),
            .I(N__14019));
    InMux I__1841 (
            .O(N__14055),
            .I(N__14019));
    InMux I__1840 (
            .O(N__14054),
            .I(N__14016));
    InMux I__1839 (
            .O(N__14053),
            .I(N__14013));
    LocalMux I__1838 (
            .O(N__14050),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1837 (
            .O(N__14047),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1836 (
            .O(N__14042),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1835 (
            .O(N__14039),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1834 (
            .O(N__14036),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv12 I__1833 (
            .O(N__14031),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1832 (
            .O(N__14026),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1831 (
            .O(N__14019),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1830 (
            .O(N__14016),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1829 (
            .O(N__14013),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__1828 (
            .O(N__13992),
            .I(N__13989));
    LocalMux I__1827 (
            .O(N__13989),
            .I(\this_vga_signals.un4_hsynclto7_0 ));
    InMux I__1826 (
            .O(N__13986),
            .I(N__13983));
    LocalMux I__1825 (
            .O(N__13983),
            .I(N__13980));
    Span4Mux_h I__1824 (
            .O(N__13980),
            .I(N__13977));
    Odrv4 I__1823 (
            .O(N__13977),
            .I(M_this_map_ram_write_data_1));
    InMux I__1822 (
            .O(N__13974),
            .I(N__13971));
    LocalMux I__1821 (
            .O(N__13971),
            .I(\this_vga_signals.SUM_2_i_1_1_1_3 ));
    CascadeMux I__1820 (
            .O(N__13968),
            .I(\this_vga_signals.N_1_3_1_cascade_ ));
    CascadeMux I__1819 (
            .O(N__13965),
            .I(N__13962));
    InMux I__1818 (
            .O(N__13962),
            .I(N__13959));
    LocalMux I__1817 (
            .O(N__13959),
            .I(\this_vga_signals.SUM_2_i_1_2_3 ));
    IoInMux I__1816 (
            .O(N__13956),
            .I(N__13953));
    LocalMux I__1815 (
            .O(N__13953),
            .I(N__13950));
    Span4Mux_s3_v I__1814 (
            .O(N__13950),
            .I(N__13947));
    Span4Mux_h I__1813 (
            .O(N__13947),
            .I(N__13944));
    Span4Mux_v I__1812 (
            .O(N__13944),
            .I(N__13941));
    Sp12to4 I__1811 (
            .O(N__13941),
            .I(N__13938));
    Span12Mux_v I__1810 (
            .O(N__13938),
            .I(N__13935));
    Odrv12 I__1809 (
            .O(N__13935),
            .I(this_vga_signals_vsync_1_i));
    InMux I__1808 (
            .O(N__13932),
            .I(N__13929));
    LocalMux I__1807 (
            .O(N__13929),
            .I(\this_vga_signals.un2_vsynclt8 ));
    InMux I__1806 (
            .O(N__13926),
            .I(N__13923));
    LocalMux I__1805 (
            .O(N__13923),
            .I(N__13917));
    InMux I__1804 (
            .O(N__13922),
            .I(N__13914));
    InMux I__1803 (
            .O(N__13921),
            .I(N__13909));
    InMux I__1802 (
            .O(N__13920),
            .I(N__13909));
    Odrv4 I__1801 (
            .O(N__13917),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d ));
    LocalMux I__1800 (
            .O(N__13914),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d ));
    LocalMux I__1799 (
            .O(N__13909),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d ));
    InMux I__1798 (
            .O(N__13902),
            .I(N__13898));
    InMux I__1797 (
            .O(N__13901),
            .I(N__13895));
    LocalMux I__1796 (
            .O(N__13898),
            .I(\this_vga_signals.mult1_un54_sum_0_3 ));
    LocalMux I__1795 (
            .O(N__13895),
            .I(\this_vga_signals.mult1_un54_sum_0_3 ));
    InMux I__1794 (
            .O(N__13890),
            .I(N__13887));
    LocalMux I__1793 (
            .O(N__13887),
            .I(N__13881));
    InMux I__1792 (
            .O(N__13886),
            .I(N__13877));
    CascadeMux I__1791 (
            .O(N__13885),
            .I(N__13874));
    CascadeMux I__1790 (
            .O(N__13884),
            .I(N__13871));
    Span4Mux_h I__1789 (
            .O(N__13881),
            .I(N__13864));
    InMux I__1788 (
            .O(N__13880),
            .I(N__13861));
    LocalMux I__1787 (
            .O(N__13877),
            .I(N__13858));
    InMux I__1786 (
            .O(N__13874),
            .I(N__13855));
    InMux I__1785 (
            .O(N__13871),
            .I(N__13848));
    InMux I__1784 (
            .O(N__13870),
            .I(N__13848));
    InMux I__1783 (
            .O(N__13869),
            .I(N__13848));
    InMux I__1782 (
            .O(N__13868),
            .I(N__13840));
    InMux I__1781 (
            .O(N__13867),
            .I(N__13837));
    Span4Mux_v I__1780 (
            .O(N__13864),
            .I(N__13832));
    LocalMux I__1779 (
            .O(N__13861),
            .I(N__13832));
    Span4Mux_v I__1778 (
            .O(N__13858),
            .I(N__13825));
    LocalMux I__1777 (
            .O(N__13855),
            .I(N__13825));
    LocalMux I__1776 (
            .O(N__13848),
            .I(N__13825));
    InMux I__1775 (
            .O(N__13847),
            .I(N__13816));
    InMux I__1774 (
            .O(N__13846),
            .I(N__13816));
    InMux I__1773 (
            .O(N__13845),
            .I(N__13816));
    InMux I__1772 (
            .O(N__13844),
            .I(N__13816));
    InMux I__1771 (
            .O(N__13843),
            .I(N__13813));
    LocalMux I__1770 (
            .O(N__13840),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1769 (
            .O(N__13837),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__1768 (
            .O(N__13832),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__1767 (
            .O(N__13825),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1766 (
            .O(N__13816),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1765 (
            .O(N__13813),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    CascadeMux I__1764 (
            .O(N__13800),
            .I(N__13788));
    InMux I__1763 (
            .O(N__13799),
            .I(N__13778));
    InMux I__1762 (
            .O(N__13798),
            .I(N__13778));
    InMux I__1761 (
            .O(N__13797),
            .I(N__13769));
    InMux I__1760 (
            .O(N__13796),
            .I(N__13769));
    InMux I__1759 (
            .O(N__13795),
            .I(N__13769));
    InMux I__1758 (
            .O(N__13794),
            .I(N__13769));
    InMux I__1757 (
            .O(N__13793),
            .I(N__13758));
    InMux I__1756 (
            .O(N__13792),
            .I(N__13758));
    InMux I__1755 (
            .O(N__13791),
            .I(N__13758));
    InMux I__1754 (
            .O(N__13788),
            .I(N__13758));
    InMux I__1753 (
            .O(N__13787),
            .I(N__13753));
    InMux I__1752 (
            .O(N__13786),
            .I(N__13753));
    CascadeMux I__1751 (
            .O(N__13785),
            .I(N__13749));
    CascadeMux I__1750 (
            .O(N__13784),
            .I(N__13744));
    InMux I__1749 (
            .O(N__13783),
            .I(N__13741));
    LocalMux I__1748 (
            .O(N__13778),
            .I(N__13736));
    LocalMux I__1747 (
            .O(N__13769),
            .I(N__13736));
    InMux I__1746 (
            .O(N__13768),
            .I(N__13731));
    InMux I__1745 (
            .O(N__13767),
            .I(N__13731));
    LocalMux I__1744 (
            .O(N__13758),
            .I(N__13728));
    LocalMux I__1743 (
            .O(N__13753),
            .I(N__13725));
    InMux I__1742 (
            .O(N__13752),
            .I(N__13721));
    InMux I__1741 (
            .O(N__13749),
            .I(N__13718));
    InMux I__1740 (
            .O(N__13748),
            .I(N__13715));
    InMux I__1739 (
            .O(N__13747),
            .I(N__13710));
    InMux I__1738 (
            .O(N__13744),
            .I(N__13710));
    LocalMux I__1737 (
            .O(N__13741),
            .I(N__13705));
    Span4Mux_v I__1736 (
            .O(N__13736),
            .I(N__13705));
    LocalMux I__1735 (
            .O(N__13731),
            .I(N__13702));
    Span4Mux_v I__1734 (
            .O(N__13728),
            .I(N__13697));
    Span4Mux_h I__1733 (
            .O(N__13725),
            .I(N__13697));
    InMux I__1732 (
            .O(N__13724),
            .I(N__13694));
    LocalMux I__1731 (
            .O(N__13721),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1730 (
            .O(N__13718),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1729 (
            .O(N__13715),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1728 (
            .O(N__13710),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1727 (
            .O(N__13705),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1726 (
            .O(N__13702),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1725 (
            .O(N__13697),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1724 (
            .O(N__13694),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    CascadeMux I__1723 (
            .O(N__13677),
            .I(\this_vga_signals.un2_hsynclto3_0_cascade_ ));
    InMux I__1722 (
            .O(N__13674),
            .I(N__13671));
    LocalMux I__1721 (
            .O(N__13671),
            .I(\this_vga_signals.M_hcounter_d7lto7_1 ));
    InMux I__1720 (
            .O(N__13668),
            .I(N__13661));
    InMux I__1719 (
            .O(N__13667),
            .I(N__13661));
    InMux I__1718 (
            .O(N__13666),
            .I(N__13656));
    LocalMux I__1717 (
            .O(N__13661),
            .I(N__13652));
    InMux I__1716 (
            .O(N__13660),
            .I(N__13649));
    InMux I__1715 (
            .O(N__13659),
            .I(N__13646));
    LocalMux I__1714 (
            .O(N__13656),
            .I(N__13640));
    InMux I__1713 (
            .O(N__13655),
            .I(N__13637));
    Span4Mux_v I__1712 (
            .O(N__13652),
            .I(N__13632));
    LocalMux I__1711 (
            .O(N__13649),
            .I(N__13632));
    LocalMux I__1710 (
            .O(N__13646),
            .I(N__13624));
    InMux I__1709 (
            .O(N__13645),
            .I(N__13621));
    InMux I__1708 (
            .O(N__13644),
            .I(N__13616));
    InMux I__1707 (
            .O(N__13643),
            .I(N__13616));
    Span4Mux_v I__1706 (
            .O(N__13640),
            .I(N__13609));
    LocalMux I__1705 (
            .O(N__13637),
            .I(N__13609));
    Span4Mux_v I__1704 (
            .O(N__13632),
            .I(N__13609));
    InMux I__1703 (
            .O(N__13631),
            .I(N__13606));
    InMux I__1702 (
            .O(N__13630),
            .I(N__13597));
    InMux I__1701 (
            .O(N__13629),
            .I(N__13597));
    InMux I__1700 (
            .O(N__13628),
            .I(N__13597));
    InMux I__1699 (
            .O(N__13627),
            .I(N__13597));
    Odrv4 I__1698 (
            .O(N__13624),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1697 (
            .O(N__13621),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1696 (
            .O(N__13616),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__1695 (
            .O(N__13609),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1694 (
            .O(N__13606),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1693 (
            .O(N__13597),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    CascadeMux I__1692 (
            .O(N__13584),
            .I(\this_vga_signals.M_hcounter_d7lt7_0_cascade_ ));
    InMux I__1691 (
            .O(N__13581),
            .I(N__13574));
    InMux I__1690 (
            .O(N__13580),
            .I(N__13574));
    InMux I__1689 (
            .O(N__13579),
            .I(N__13571));
    LocalMux I__1688 (
            .O(N__13574),
            .I(N__13565));
    LocalMux I__1687 (
            .O(N__13571),
            .I(N__13556));
    InMux I__1686 (
            .O(N__13570),
            .I(N__13549));
    InMux I__1685 (
            .O(N__13569),
            .I(N__13549));
    InMux I__1684 (
            .O(N__13568),
            .I(N__13549));
    Span4Mux_h I__1683 (
            .O(N__13565),
            .I(N__13546));
    InMux I__1682 (
            .O(N__13564),
            .I(N__13543));
    CascadeMux I__1681 (
            .O(N__13563),
            .I(N__13539));
    CascadeMux I__1680 (
            .O(N__13562),
            .I(N__13536));
    CascadeMux I__1679 (
            .O(N__13561),
            .I(N__13533));
    InMux I__1678 (
            .O(N__13560),
            .I(N__13529));
    InMux I__1677 (
            .O(N__13559),
            .I(N__13526));
    Span4Mux_v I__1676 (
            .O(N__13556),
            .I(N__13521));
    LocalMux I__1675 (
            .O(N__13549),
            .I(N__13521));
    Span4Mux_v I__1674 (
            .O(N__13546),
            .I(N__13516));
    LocalMux I__1673 (
            .O(N__13543),
            .I(N__13516));
    InMux I__1672 (
            .O(N__13542),
            .I(N__13513));
    InMux I__1671 (
            .O(N__13539),
            .I(N__13504));
    InMux I__1670 (
            .O(N__13536),
            .I(N__13504));
    InMux I__1669 (
            .O(N__13533),
            .I(N__13504));
    InMux I__1668 (
            .O(N__13532),
            .I(N__13504));
    LocalMux I__1667 (
            .O(N__13529),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1666 (
            .O(N__13526),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__1665 (
            .O(N__13521),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__1664 (
            .O(N__13516),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1663 (
            .O(N__13513),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1662 (
            .O(N__13504),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    CascadeMux I__1661 (
            .O(N__13491),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_cascade_ ));
    InMux I__1660 (
            .O(N__13488),
            .I(N__13484));
    InMux I__1659 (
            .O(N__13487),
            .I(N__13481));
    LocalMux I__1658 (
            .O(N__13484),
            .I(N__13478));
    LocalMux I__1657 (
            .O(N__13481),
            .I(\this_vga_signals.g0_0_0_a2_0 ));
    Odrv4 I__1656 (
            .O(N__13478),
            .I(\this_vga_signals.g0_0_0_a2_0 ));
    InMux I__1655 (
            .O(N__13473),
            .I(N__13467));
    InMux I__1654 (
            .O(N__13472),
            .I(N__13462));
    InMux I__1653 (
            .O(N__13471),
            .I(N__13462));
    InMux I__1652 (
            .O(N__13470),
            .I(N__13459));
    LocalMux I__1651 (
            .O(N__13467),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1650 (
            .O(N__13462),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1649 (
            .O(N__13459),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    InMux I__1648 (
            .O(N__13452),
            .I(N__13446));
    CascadeMux I__1647 (
            .O(N__13451),
            .I(N__13438));
    CascadeMux I__1646 (
            .O(N__13450),
            .I(N__13432));
    InMux I__1645 (
            .O(N__13449),
            .I(N__13429));
    LocalMux I__1644 (
            .O(N__13446),
            .I(N__13426));
    InMux I__1643 (
            .O(N__13445),
            .I(N__13423));
    InMux I__1642 (
            .O(N__13444),
            .I(N__13420));
    InMux I__1641 (
            .O(N__13443),
            .I(N__13417));
    InMux I__1640 (
            .O(N__13442),
            .I(N__13408));
    InMux I__1639 (
            .O(N__13441),
            .I(N__13408));
    InMux I__1638 (
            .O(N__13438),
            .I(N__13408));
    InMux I__1637 (
            .O(N__13437),
            .I(N__13408));
    InMux I__1636 (
            .O(N__13436),
            .I(N__13401));
    InMux I__1635 (
            .O(N__13435),
            .I(N__13401));
    InMux I__1634 (
            .O(N__13432),
            .I(N__13401));
    LocalMux I__1633 (
            .O(N__13429),
            .I(N__13398));
    Odrv4 I__1632 (
            .O(N__13426),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1631 (
            .O(N__13423),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1630 (
            .O(N__13420),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1629 (
            .O(N__13417),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1628 (
            .O(N__13408),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1627 (
            .O(N__13401),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    Odrv4 I__1626 (
            .O(N__13398),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    CascadeMux I__1625 (
            .O(N__13383),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_0_cascade_ ));
    InMux I__1624 (
            .O(N__13380),
            .I(N__13371));
    InMux I__1623 (
            .O(N__13379),
            .I(N__13368));
    CascadeMux I__1622 (
            .O(N__13378),
            .I(N__13360));
    CascadeMux I__1621 (
            .O(N__13377),
            .I(N__13356));
    CascadeMux I__1620 (
            .O(N__13376),
            .I(N__13353));
    InMux I__1619 (
            .O(N__13375),
            .I(N__13350));
    InMux I__1618 (
            .O(N__13374),
            .I(N__13347));
    LocalMux I__1617 (
            .O(N__13371),
            .I(N__13342));
    LocalMux I__1616 (
            .O(N__13368),
            .I(N__13342));
    InMux I__1615 (
            .O(N__13367),
            .I(N__13335));
    InMux I__1614 (
            .O(N__13366),
            .I(N__13335));
    InMux I__1613 (
            .O(N__13365),
            .I(N__13335));
    InMux I__1612 (
            .O(N__13364),
            .I(N__13332));
    InMux I__1611 (
            .O(N__13363),
            .I(N__13329));
    InMux I__1610 (
            .O(N__13360),
            .I(N__13322));
    InMux I__1609 (
            .O(N__13359),
            .I(N__13322));
    InMux I__1608 (
            .O(N__13356),
            .I(N__13322));
    InMux I__1607 (
            .O(N__13353),
            .I(N__13319));
    LocalMux I__1606 (
            .O(N__13350),
            .I(\this_vga_signals.mult1_un68_sum_axb1_661 ));
    LocalMux I__1605 (
            .O(N__13347),
            .I(\this_vga_signals.mult1_un68_sum_axb1_661 ));
    Odrv4 I__1604 (
            .O(N__13342),
            .I(\this_vga_signals.mult1_un68_sum_axb1_661 ));
    LocalMux I__1603 (
            .O(N__13335),
            .I(\this_vga_signals.mult1_un68_sum_axb1_661 ));
    LocalMux I__1602 (
            .O(N__13332),
            .I(\this_vga_signals.mult1_un68_sum_axb1_661 ));
    LocalMux I__1601 (
            .O(N__13329),
            .I(\this_vga_signals.mult1_un68_sum_axb1_661 ));
    LocalMux I__1600 (
            .O(N__13322),
            .I(\this_vga_signals.mult1_un68_sum_axb1_661 ));
    LocalMux I__1599 (
            .O(N__13319),
            .I(\this_vga_signals.mult1_un68_sum_axb1_661 ));
    InMux I__1598 (
            .O(N__13302),
            .I(N__13299));
    LocalMux I__1597 (
            .O(N__13299),
            .I(\this_vga_signals.g0_i_x4_0_a3_2 ));
    CascadeMux I__1596 (
            .O(N__13296),
            .I(N__13293));
    InMux I__1595 (
            .O(N__13293),
            .I(N__13290));
    LocalMux I__1594 (
            .O(N__13290),
            .I(N__13287));
    Odrv4 I__1593 (
            .O(N__13287),
            .I(\this_vga_signals.vaddress_0_6 ));
    InMux I__1592 (
            .O(N__13284),
            .I(N__13281));
    LocalMux I__1591 (
            .O(N__13281),
            .I(\this_vga_signals.g0_i_x4_0_a3_0 ));
    InMux I__1590 (
            .O(N__13278),
            .I(N__13275));
    LocalMux I__1589 (
            .O(N__13275),
            .I(\this_vga_signals.vsync_1_3 ));
    CascadeMux I__1588 (
            .O(N__13272),
            .I(\this_vga_signals.vsync_1_2_cascade_ ));
    CascadeMux I__1587 (
            .O(N__13269),
            .I(\this_vga_signals.mult1_un68_sum_axb1_661_cascade_ ));
    InMux I__1586 (
            .O(N__13266),
            .I(N__13263));
    LocalMux I__1585 (
            .O(N__13263),
            .I(\this_vga_signals.g0_2_0_a2_1 ));
    CascadeMux I__1584 (
            .O(N__13260),
            .I(\this_vga_signals.if_N_5_cascade_ ));
    CascadeMux I__1583 (
            .O(N__13257),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ));
    CascadeMux I__1582 (
            .O(N__13254),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_1_cascade_ ));
    CascadeMux I__1581 (
            .O(N__13251),
            .I(\this_vga_signals.mult1_un61_sum_c3_cascade_ ));
    InMux I__1580 (
            .O(N__13248),
            .I(N__13242));
    InMux I__1579 (
            .O(N__13247),
            .I(N__13242));
    LocalMux I__1578 (
            .O(N__13242),
            .I(N__13239));
    Odrv4 I__1577 (
            .O(N__13239),
            .I(\this_vga_signals.N_4_0_1_0 ));
    CascadeMux I__1576 (
            .O(N__13236),
            .I(\this_vga_signals.mult1_un47_sum_c3_cascade_ ));
    InMux I__1575 (
            .O(N__13233),
            .I(N__13230));
    LocalMux I__1574 (
            .O(N__13230),
            .I(\this_vga_signals.g1_2 ));
    CascadeMux I__1573 (
            .O(N__13227),
            .I(\this_vga_signals.SUM_3_0_cascade_ ));
    CascadeMux I__1572 (
            .O(N__13224),
            .I(N__13221));
    InMux I__1571 (
            .O(N__13221),
            .I(N__13218));
    LocalMux I__1570 (
            .O(N__13218),
            .I(\this_vga_signals.mult1_un61_sum_axb1_0 ));
    InMux I__1569 (
            .O(N__13215),
            .I(N__13212));
    LocalMux I__1568 (
            .O(N__13212),
            .I(N__13209));
    Span4Mux_v I__1567 (
            .O(N__13209),
            .I(N__13206));
    Odrv4 I__1566 (
            .O(N__13206),
            .I(M_this_map_ram_write_data_4));
    InMux I__1565 (
            .O(N__13203),
            .I(N__13200));
    LocalMux I__1564 (
            .O(N__13200),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i_0 ));
    CascadeMux I__1563 (
            .O(N__13197),
            .I(\this_vga_signals.N_18_cascade_ ));
    InMux I__1562 (
            .O(N__13194),
            .I(N__13191));
    LocalMux I__1561 (
            .O(N__13191),
            .I(\this_vga_signals.g1_0_0_1 ));
    InMux I__1560 (
            .O(N__13188),
            .I(N__13185));
    LocalMux I__1559 (
            .O(N__13185),
            .I(\this_vga_signals.vaddress_1_6 ));
    CascadeMux I__1558 (
            .O(N__13182),
            .I(\this_vga_signals.N_6_cascade_ ));
    InMux I__1557 (
            .O(N__13179),
            .I(N__13173));
    InMux I__1556 (
            .O(N__13178),
            .I(N__13173));
    LocalMux I__1555 (
            .O(N__13173),
            .I(\this_vga_signals.g1_1_1 ));
    InMux I__1554 (
            .O(N__13170),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__1553 (
            .O(N__13167),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__1552 (
            .O(N__13164),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__1551 (
            .O(N__13161),
            .I(bfn_11_14_0_));
    InMux I__1550 (
            .O(N__13158),
            .I(N__13155));
    LocalMux I__1549 (
            .O(N__13155),
            .I(\this_vga_signals.un4_hsynclt9 ));
    InMux I__1548 (
            .O(N__13152),
            .I(N__13147));
    InMux I__1547 (
            .O(N__13151),
            .I(N__13144));
    InMux I__1546 (
            .O(N__13150),
            .I(N__13141));
    LocalMux I__1545 (
            .O(N__13147),
            .I(N__13138));
    LocalMux I__1544 (
            .O(N__13144),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__1543 (
            .O(N__13141),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    Odrv4 I__1542 (
            .O(N__13138),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    CascadeMux I__1541 (
            .O(N__13131),
            .I(N__13127));
    CascadeMux I__1540 (
            .O(N__13130),
            .I(N__13123));
    InMux I__1539 (
            .O(N__13127),
            .I(N__13120));
    InMux I__1538 (
            .O(N__13126),
            .I(N__13115));
    InMux I__1537 (
            .O(N__13123),
            .I(N__13115));
    LocalMux I__1536 (
            .O(N__13120),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    LocalMux I__1535 (
            .O(N__13115),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    CascadeMux I__1534 (
            .O(N__13110),
            .I(\this_vga_signals.M_pcounter_q_3_1_cascade_ ));
    InMux I__1533 (
            .O(N__13107),
            .I(N__13101));
    InMux I__1532 (
            .O(N__13106),
            .I(N__13101));
    LocalMux I__1531 (
            .O(N__13101),
            .I(N__13098));
    Odrv4 I__1530 (
            .O(N__13098),
            .I(N_3_0));
    CascadeMux I__1529 (
            .O(N__13095),
            .I(N_3_0_cascade_));
    InMux I__1528 (
            .O(N__13092),
            .I(N__13089));
    LocalMux I__1527 (
            .O(N__13089),
            .I(N__13083));
    InMux I__1526 (
            .O(N__13088),
            .I(N__13078));
    InMux I__1525 (
            .O(N__13087),
            .I(N__13078));
    InMux I__1524 (
            .O(N__13086),
            .I(N__13075));
    Span4Mux_h I__1523 (
            .O(N__13083),
            .I(N__13072));
    LocalMux I__1522 (
            .O(N__13078),
            .I(\this_vga_signals.M_pcounter_q_i_3_1 ));
    LocalMux I__1521 (
            .O(N__13075),
            .I(\this_vga_signals.M_pcounter_q_i_3_1 ));
    Odrv4 I__1520 (
            .O(N__13072),
            .I(\this_vga_signals.M_pcounter_q_i_3_1 ));
    InMux I__1519 (
            .O(N__13065),
            .I(N__13062));
    LocalMux I__1518 (
            .O(N__13062),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_1 ));
    InMux I__1517 (
            .O(N__13059),
            .I(N__13056));
    LocalMux I__1516 (
            .O(N__13056),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_a0_0 ));
    InMux I__1515 (
            .O(N__13053),
            .I(N__13046));
    InMux I__1514 (
            .O(N__13052),
            .I(N__13042));
    CascadeMux I__1513 (
            .O(N__13051),
            .I(N__13038));
    CascadeMux I__1512 (
            .O(N__13050),
            .I(N__13033));
    InMux I__1511 (
            .O(N__13049),
            .I(N__13027));
    LocalMux I__1510 (
            .O(N__13046),
            .I(N__13024));
    InMux I__1509 (
            .O(N__13045),
            .I(N__13021));
    LocalMux I__1508 (
            .O(N__13042),
            .I(N__13018));
    InMux I__1507 (
            .O(N__13041),
            .I(N__13015));
    InMux I__1506 (
            .O(N__13038),
            .I(N__13008));
    InMux I__1505 (
            .O(N__13037),
            .I(N__13008));
    InMux I__1504 (
            .O(N__13036),
            .I(N__13008));
    InMux I__1503 (
            .O(N__13033),
            .I(N__12999));
    InMux I__1502 (
            .O(N__13032),
            .I(N__12999));
    InMux I__1501 (
            .O(N__13031),
            .I(N__12999));
    InMux I__1500 (
            .O(N__13030),
            .I(N__12999));
    LocalMux I__1499 (
            .O(N__13027),
            .I(\this_vga_signals.SUM_3 ));
    Odrv4 I__1498 (
            .O(N__13024),
            .I(\this_vga_signals.SUM_3 ));
    LocalMux I__1497 (
            .O(N__13021),
            .I(\this_vga_signals.SUM_3 ));
    Odrv4 I__1496 (
            .O(N__13018),
            .I(\this_vga_signals.SUM_3 ));
    LocalMux I__1495 (
            .O(N__13015),
            .I(\this_vga_signals.SUM_3 ));
    LocalMux I__1494 (
            .O(N__13008),
            .I(\this_vga_signals.SUM_3 ));
    LocalMux I__1493 (
            .O(N__12999),
            .I(\this_vga_signals.SUM_3 ));
    CascadeMux I__1492 (
            .O(N__12984),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz_cascade_ ));
    InMux I__1491 (
            .O(N__12981),
            .I(N__12976));
    InMux I__1490 (
            .O(N__12980),
            .I(N__12970));
    InMux I__1489 (
            .O(N__12979),
            .I(N__12962));
    LocalMux I__1488 (
            .O(N__12976),
            .I(N__12959));
    InMux I__1487 (
            .O(N__12975),
            .I(N__12956));
    InMux I__1486 (
            .O(N__12974),
            .I(N__12951));
    InMux I__1485 (
            .O(N__12973),
            .I(N__12951));
    LocalMux I__1484 (
            .O(N__12970),
            .I(N__12948));
    InMux I__1483 (
            .O(N__12969),
            .I(N__12945));
    InMux I__1482 (
            .O(N__12968),
            .I(N__12936));
    InMux I__1481 (
            .O(N__12967),
            .I(N__12936));
    InMux I__1480 (
            .O(N__12966),
            .I(N__12936));
    InMux I__1479 (
            .O(N__12965),
            .I(N__12936));
    LocalMux I__1478 (
            .O(N__12962),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9 ));
    Odrv4 I__1477 (
            .O(N__12959),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9 ));
    LocalMux I__1476 (
            .O(N__12956),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9 ));
    LocalMux I__1475 (
            .O(N__12951),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9 ));
    Odrv4 I__1474 (
            .O(N__12948),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9 ));
    LocalMux I__1473 (
            .O(N__12945),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9 ));
    LocalMux I__1472 (
            .O(N__12936),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9 ));
    InMux I__1471 (
            .O(N__12921),
            .I(N__12918));
    LocalMux I__1470 (
            .O(N__12918),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ));
    InMux I__1469 (
            .O(N__12915),
            .I(N__12912));
    LocalMux I__1468 (
            .O(N__12912),
            .I(\this_vga_signals.if_N_6_0 ));
    InMux I__1467 (
            .O(N__12909),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__1466 (
            .O(N__12906),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__1465 (
            .O(N__12903),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__1464 (
            .O(N__12900),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__1463 (
            .O(N__12897),
            .I(N__12894));
    LocalMux I__1462 (
            .O(N__12894),
            .I(\this_vga_signals.g1_0 ));
    CascadeMux I__1461 (
            .O(N__12891),
            .I(\this_vga_signals.g0_i_x4_2_0_0_1_cascade_ ));
    CascadeMux I__1460 (
            .O(N__12888),
            .I(N__12885));
    InMux I__1459 (
            .O(N__12885),
            .I(N__12882));
    LocalMux I__1458 (
            .O(N__12882),
            .I(\this_vga_signals.g0_i_x4_0_0 ));
    CascadeMux I__1457 (
            .O(N__12879),
            .I(\this_vga_signals.N_3_cascade_ ));
    InMux I__1456 (
            .O(N__12876),
            .I(N__12873));
    LocalMux I__1455 (
            .O(N__12873),
            .I(\this_vga_signals.N_4_0_0 ));
    CascadeMux I__1454 (
            .O(N__12870),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0_0_cascade_ ));
    InMux I__1453 (
            .O(N__12867),
            .I(N__12864));
    LocalMux I__1452 (
            .O(N__12864),
            .I(N__12861));
    Odrv4 I__1451 (
            .O(N__12861),
            .I(\this_vga_signals.mult1_un75_sum_c2_0_0_0 ));
    CascadeMux I__1450 (
            .O(N__12858),
            .I(N__12855));
    InMux I__1449 (
            .O(N__12855),
            .I(N__12852));
    LocalMux I__1448 (
            .O(N__12852),
            .I(\this_vga_signals.g0_2_1 ));
    CascadeMux I__1447 (
            .O(N__12849),
            .I(N__12844));
    InMux I__1446 (
            .O(N__12848),
            .I(N__12841));
    InMux I__1445 (
            .O(N__12847),
            .I(N__12836));
    InMux I__1444 (
            .O(N__12844),
            .I(N__12836));
    LocalMux I__1443 (
            .O(N__12841),
            .I(\this_vga_signals.N_5_0_0 ));
    LocalMux I__1442 (
            .O(N__12836),
            .I(\this_vga_signals.N_5_0_0 ));
    InMux I__1441 (
            .O(N__12831),
            .I(N__12828));
    LocalMux I__1440 (
            .O(N__12828),
            .I(N__12825));
    Span4Mux_v I__1439 (
            .O(N__12825),
            .I(N__12822));
    Span4Mux_v I__1438 (
            .O(N__12822),
            .I(N__12818));
    InMux I__1437 (
            .O(N__12821),
            .I(N__12815));
    Odrv4 I__1436 (
            .O(N__12818),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1435 (
            .O(N__12815),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    InMux I__1434 (
            .O(N__12810),
            .I(N__12807));
    LocalMux I__1433 (
            .O(N__12807),
            .I(\this_vga_signals.mult1_un68_sum_ac0_2 ));
    CascadeMux I__1432 (
            .O(N__12804),
            .I(\this_vga_signals.mult1_un68_sum_ac0_2_cascade_ ));
    InMux I__1431 (
            .O(N__12801),
            .I(N__12798));
    LocalMux I__1430 (
            .O(N__12798),
            .I(\this_vga_signals.g1_0_3 ));
    InMux I__1429 (
            .O(N__12795),
            .I(N__12792));
    LocalMux I__1428 (
            .O(N__12792),
            .I(\this_vga_signals.g0_2_0_a2 ));
    CascadeMux I__1427 (
            .O(N__12789),
            .I(N__12786));
    InMux I__1426 (
            .O(N__12786),
            .I(N__12780));
    InMux I__1425 (
            .O(N__12785),
            .I(N__12780));
    LocalMux I__1424 (
            .O(N__12780),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    CascadeMux I__1423 (
            .O(N__12777),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ));
    InMux I__1422 (
            .O(N__12774),
            .I(N__12771));
    LocalMux I__1421 (
            .O(N__12771),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    InMux I__1420 (
            .O(N__12768),
            .I(N__12765));
    LocalMux I__1419 (
            .O(N__12765),
            .I(\this_vga_signals.g0_1_2 ));
    InMux I__1418 (
            .O(N__12762),
            .I(N__12759));
    LocalMux I__1417 (
            .O(N__12759),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_x1 ));
    CascadeMux I__1416 (
            .O(N__12756),
            .I(\this_vga_signals.g3_0_cascade_ ));
    InMux I__1415 (
            .O(N__12753),
            .I(N__12750));
    LocalMux I__1414 (
            .O(N__12750),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0_2 ));
    CascadeMux I__1413 (
            .O(N__12747),
            .I(\this_vga_signals.g0_0_a2_0_0_cascade_ ));
    InMux I__1412 (
            .O(N__12744),
            .I(N__12741));
    LocalMux I__1411 (
            .O(N__12741),
            .I(\this_vga_signals.g1_0_a2_1 ));
    CascadeMux I__1410 (
            .O(N__12738),
            .I(N__12735));
    InMux I__1409 (
            .O(N__12735),
            .I(N__12732));
    LocalMux I__1408 (
            .O(N__12732),
            .I(\this_vga_signals.vaddress_1_5 ));
    CascadeMux I__1407 (
            .O(N__12729),
            .I(N__12726));
    InMux I__1406 (
            .O(N__12726),
            .I(N__12723));
    LocalMux I__1405 (
            .O(N__12723),
            .I(N__12720));
    Span4Mux_h I__1404 (
            .O(N__12720),
            .I(N__12717));
    Odrv4 I__1403 (
            .O(N__12717),
            .I(\this_vga_signals.mult1_un47_sum_c3_0_0 ));
    CascadeMux I__1402 (
            .O(N__12714),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_x0_cascade_ ));
    InMux I__1401 (
            .O(N__12711),
            .I(N__12708));
    LocalMux I__1400 (
            .O(N__12708),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_ns ));
    CascadeMux I__1399 (
            .O(N__12705),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_ns_cascade_ ));
    InMux I__1398 (
            .O(N__12702),
            .I(N__12699));
    LocalMux I__1397 (
            .O(N__12699),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_0 ));
    InMux I__1396 (
            .O(N__12696),
            .I(N__12693));
    LocalMux I__1395 (
            .O(N__12693),
            .I(\this_vga_signals.g0_i_x4_1 ));
    InMux I__1394 (
            .O(N__12690),
            .I(N__12687));
    LocalMux I__1393 (
            .O(N__12687),
            .I(\this_vga_signals.g0_i_x4_0_1 ));
    InMux I__1392 (
            .O(N__12684),
            .I(N__12681));
    LocalMux I__1391 (
            .O(N__12681),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0 ));
    InMux I__1390 (
            .O(N__12678),
            .I(N__12674));
    InMux I__1389 (
            .O(N__12677),
            .I(N__12670));
    LocalMux I__1388 (
            .O(N__12674),
            .I(N__12666));
    InMux I__1387 (
            .O(N__12673),
            .I(N__12663));
    LocalMux I__1386 (
            .O(N__12670),
            .I(N__12660));
    InMux I__1385 (
            .O(N__12669),
            .I(N__12657));
    Span4Mux_v I__1384 (
            .O(N__12666),
            .I(N__12641));
    LocalMux I__1383 (
            .O(N__12663),
            .I(N__12641));
    Span4Mux_v I__1382 (
            .O(N__12660),
            .I(N__12636));
    LocalMux I__1381 (
            .O(N__12657),
            .I(N__12636));
    InMux I__1380 (
            .O(N__12656),
            .I(N__12631));
    InMux I__1379 (
            .O(N__12655),
            .I(N__12631));
    InMux I__1378 (
            .O(N__12654),
            .I(N__12624));
    InMux I__1377 (
            .O(N__12653),
            .I(N__12624));
    InMux I__1376 (
            .O(N__12652),
            .I(N__12624));
    InMux I__1375 (
            .O(N__12651),
            .I(N__12619));
    InMux I__1374 (
            .O(N__12650),
            .I(N__12619));
    InMux I__1373 (
            .O(N__12649),
            .I(N__12616));
    InMux I__1372 (
            .O(N__12648),
            .I(N__12609));
    InMux I__1371 (
            .O(N__12647),
            .I(N__12609));
    InMux I__1370 (
            .O(N__12646),
            .I(N__12609));
    Odrv4 I__1369 (
            .O(N__12641),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    Odrv4 I__1368 (
            .O(N__12636),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1367 (
            .O(N__12631),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1366 (
            .O(N__12624),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1365 (
            .O(N__12619),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1364 (
            .O(N__12616),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1363 (
            .O(N__12609),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    InMux I__1362 (
            .O(N__12594),
            .I(N__12591));
    LocalMux I__1361 (
            .O(N__12591),
            .I(N__12588));
    Odrv4 I__1360 (
            .O(N__12588),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0 ));
    InMux I__1359 (
            .O(N__12585),
            .I(N__12581));
    InMux I__1358 (
            .O(N__12584),
            .I(N__12578));
    LocalMux I__1357 (
            .O(N__12581),
            .I(N__12573));
    LocalMux I__1356 (
            .O(N__12578),
            .I(N__12573));
    Odrv4 I__1355 (
            .O(N__12573),
            .I(\this_vga_signals.SUM_3_0_0 ));
    InMux I__1354 (
            .O(N__12570),
            .I(N__12566));
    InMux I__1353 (
            .O(N__12569),
            .I(N__12563));
    LocalMux I__1352 (
            .O(N__12566),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    LocalMux I__1351 (
            .O(N__12563),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    IoInMux I__1350 (
            .O(N__12558),
            .I(N__12555));
    LocalMux I__1349 (
            .O(N__12555),
            .I(N__12552));
    IoSpan4Mux I__1348 (
            .O(N__12552),
            .I(N__12549));
    Span4Mux_s3_v I__1347 (
            .O(N__12549),
            .I(N__12546));
    Sp12to4 I__1346 (
            .O(N__12546),
            .I(N__12543));
    Span12Mux_v I__1345 (
            .O(N__12543),
            .I(N__12540));
    Odrv12 I__1344 (
            .O(N__12540),
            .I(this_vga_signals_hsync_1_i));
    IoInMux I__1343 (
            .O(N__12537),
            .I(N__12534));
    LocalMux I__1342 (
            .O(N__12534),
            .I(N__12531));
    Span4Mux_s3_v I__1341 (
            .O(N__12531),
            .I(N__12528));
    Sp12to4 I__1340 (
            .O(N__12528),
            .I(N__12525));
    Span12Mux_s11_h I__1339 (
            .O(N__12525),
            .I(N__12522));
    Span12Mux_v I__1338 (
            .O(N__12522),
            .I(N__12519));
    Odrv12 I__1337 (
            .O(N__12519),
            .I(this_vga_signals_hvisibility_i));
    CascadeMux I__1336 (
            .O(N__12516),
            .I(\this_vga_signals.g3_0_1_cascade_ ));
    InMux I__1335 (
            .O(N__12513),
            .I(N__12510));
    LocalMux I__1334 (
            .O(N__12510),
            .I(\this_vga_signals.g3_0 ));
    CascadeMux I__1333 (
            .O(N__12507),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_ ));
    InMux I__1332 (
            .O(N__12504),
            .I(N__12497));
    InMux I__1331 (
            .O(N__12503),
            .I(N__12490));
    InMux I__1330 (
            .O(N__12502),
            .I(N__12490));
    InMux I__1329 (
            .O(N__12501),
            .I(N__12490));
    InMux I__1328 (
            .O(N__12500),
            .I(N__12487));
    LocalMux I__1327 (
            .O(N__12497),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_1 ));
    LocalMux I__1326 (
            .O(N__12490),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_1 ));
    LocalMux I__1325 (
            .O(N__12487),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_1 ));
    InMux I__1324 (
            .O(N__12480),
            .I(N__12477));
    LocalMux I__1323 (
            .O(N__12477),
            .I(\this_vga_signals.N_6_1_0 ));
    InMux I__1322 (
            .O(N__12474),
            .I(N__12471));
    LocalMux I__1321 (
            .O(N__12471),
            .I(N__12468));
    Span4Mux_v I__1320 (
            .O(N__12468),
            .I(N__12464));
    InMux I__1319 (
            .O(N__12467),
            .I(N__12461));
    Odrv4 I__1318 (
            .O(N__12464),
            .I(\this_vga_signals.N_234 ));
    LocalMux I__1317 (
            .O(N__12461),
            .I(\this_vga_signals.N_234 ));
    CascadeMux I__1316 (
            .O(N__12456),
            .I(\this_vga_signals.SUM_3_cascade_ ));
    CascadeMux I__1315 (
            .O(N__12453),
            .I(N__12450));
    InMux I__1314 (
            .O(N__12450),
            .I(N__12447));
    LocalMux I__1313 (
            .O(N__12447),
            .I(\this_vga_signals.g0_6_1 ));
    CascadeMux I__1312 (
            .O(N__12444),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9_cascade_ ));
    InMux I__1311 (
            .O(N__12441),
            .I(N__12438));
    LocalMux I__1310 (
            .O(N__12438),
            .I(\this_vga_signals.mult1_un61_sum_axb1_1 ));
    InMux I__1309 (
            .O(N__12435),
            .I(N__12432));
    LocalMux I__1308 (
            .O(N__12432),
            .I(N__12429));
    Span4Mux_h I__1307 (
            .O(N__12429),
            .I(N__12426));
    Odrv4 I__1306 (
            .O(N__12426),
            .I(\this_vga_signals.g1_2_0_0 ));
    InMux I__1305 (
            .O(N__12423),
            .I(N__12420));
    LocalMux I__1304 (
            .O(N__12420),
            .I(N__12415));
    InMux I__1303 (
            .O(N__12419),
            .I(N__12410));
    InMux I__1302 (
            .O(N__12418),
            .I(N__12410));
    Span4Mux_h I__1301 (
            .O(N__12415),
            .I(N__12405));
    LocalMux I__1300 (
            .O(N__12410),
            .I(N__12405));
    Odrv4 I__1299 (
            .O(N__12405),
            .I(\this_vga_signals.mult1_un68_sum_axb1 ));
    InMux I__1298 (
            .O(N__12402),
            .I(N__12399));
    LocalMux I__1297 (
            .O(N__12399),
            .I(\this_vga_signals.g1_7 ));
    InMux I__1296 (
            .O(N__12396),
            .I(N__12393));
    LocalMux I__1295 (
            .O(N__12393),
            .I(\this_vga_signals.g0_i_x4_3_0 ));
    CascadeMux I__1294 (
            .O(N__12390),
            .I(\this_vga_signals.mult1_un61_sum_axb1_3_0_cascade_ ));
    InMux I__1293 (
            .O(N__12387),
            .I(N__12384));
    LocalMux I__1292 (
            .O(N__12384),
            .I(\this_vga_signals.g1_1_0 ));
    InMux I__1291 (
            .O(N__12381),
            .I(N__12378));
    LocalMux I__1290 (
            .O(N__12378),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_1 ));
    CascadeMux I__1289 (
            .O(N__12375),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_1_cascade_ ));
    InMux I__1288 (
            .O(N__12372),
            .I(N__12369));
    LocalMux I__1287 (
            .O(N__12369),
            .I(\this_vga_signals.g1_0_1_0 ));
    CascadeMux I__1286 (
            .O(N__12366),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_ ));
    CascadeMux I__1285 (
            .O(N__12363),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_3_cascade_ ));
    CascadeMux I__1284 (
            .O(N__12360),
            .I(N__12357));
    InMux I__1283 (
            .O(N__12357),
            .I(N__12354));
    LocalMux I__1282 (
            .O(N__12354),
            .I(N__12348));
    InMux I__1281 (
            .O(N__12353),
            .I(N__12343));
    InMux I__1280 (
            .O(N__12352),
            .I(N__12343));
    InMux I__1279 (
            .O(N__12351),
            .I(N__12340));
    Odrv12 I__1278 (
            .O(N__12348),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0));
    LocalMux I__1277 (
            .O(N__12343),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0));
    LocalMux I__1276 (
            .O(N__12340),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0));
    CascadeMux I__1275 (
            .O(N__12333),
            .I(N__12329));
    InMux I__1274 (
            .O(N__12332),
            .I(N__12325));
    InMux I__1273 (
            .O(N__12329),
            .I(N__12320));
    InMux I__1272 (
            .O(N__12328),
            .I(N__12320));
    LocalMux I__1271 (
            .O(N__12325),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0));
    LocalMux I__1270 (
            .O(N__12320),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0));
    InMux I__1269 (
            .O(N__12315),
            .I(N__12312));
    LocalMux I__1268 (
            .O(N__12312),
            .I(N__12309));
    Span4Mux_h I__1267 (
            .O(N__12309),
            .I(N__12306));
    Odrv4 I__1266 (
            .O(N__12306),
            .I(\this_vga_signals.d_N_3_1_i ));
    InMux I__1265 (
            .O(N__12303),
            .I(N__12300));
    LocalMux I__1264 (
            .O(N__12300),
            .I(\this_vga_signals.M_hcounter_q_RNIO08E8Z0Z_3 ));
    CascadeMux I__1263 (
            .O(N__12297),
            .I(N__12289));
    CascadeMux I__1262 (
            .O(N__12296),
            .I(N__12286));
    InMux I__1261 (
            .O(N__12295),
            .I(N__12282));
    InMux I__1260 (
            .O(N__12294),
            .I(N__12277));
    InMux I__1259 (
            .O(N__12293),
            .I(N__12277));
    InMux I__1258 (
            .O(N__12292),
            .I(N__12268));
    InMux I__1257 (
            .O(N__12289),
            .I(N__12268));
    InMux I__1256 (
            .O(N__12286),
            .I(N__12268));
    InMux I__1255 (
            .O(N__12285),
            .I(N__12268));
    LocalMux I__1254 (
            .O(N__12282),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3));
    LocalMux I__1253 (
            .O(N__12277),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3));
    LocalMux I__1252 (
            .O(N__12268),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3));
    CascadeMux I__1251 (
            .O(N__12261),
            .I(\this_vga_signals.g1_0_1_cascade_ ));
    CascadeMux I__1250 (
            .O(N__12258),
            .I(\this_vga_signals.g1_2_0_cascade_ ));
    CascadeMux I__1249 (
            .O(N__12255),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_0_0_cascade_ ));
    InMux I__1248 (
            .O(N__12252),
            .I(N__12249));
    LocalMux I__1247 (
            .O(N__12249),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1_0_0_1 ));
    InMux I__1246 (
            .O(N__12246),
            .I(N__12243));
    LocalMux I__1245 (
            .O(N__12243),
            .I(\this_vga_signals.mult1_un89_sum_c3_1_0_0_1 ));
    InMux I__1244 (
            .O(N__12240),
            .I(N__12230));
    InMux I__1243 (
            .O(N__12239),
            .I(N__12221));
    InMux I__1242 (
            .O(N__12238),
            .I(N__12221));
    InMux I__1241 (
            .O(N__12237),
            .I(N__12221));
    InMux I__1240 (
            .O(N__12236),
            .I(N__12221));
    InMux I__1239 (
            .O(N__12235),
            .I(N__12218));
    InMux I__1238 (
            .O(N__12234),
            .I(N__12213));
    InMux I__1237 (
            .O(N__12233),
            .I(N__12213));
    LocalMux I__1236 (
            .O(N__12230),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0));
    LocalMux I__1235 (
            .O(N__12221),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0));
    LocalMux I__1234 (
            .O(N__12218),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0));
    LocalMux I__1233 (
            .O(N__12213),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0));
    InMux I__1232 (
            .O(N__12204),
            .I(N__12201));
    LocalMux I__1231 (
            .O(N__12201),
            .I(\this_vga_signals.N_4_2 ));
    CascadeMux I__1230 (
            .O(N__12198),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_0_cascade_ ));
    CascadeMux I__1229 (
            .O(N__12195),
            .I(N__12192));
    InMux I__1228 (
            .O(N__12192),
            .I(N__12189));
    LocalMux I__1227 (
            .O(N__12189),
            .I(N__12186));
    Span4Mux_h I__1226 (
            .O(N__12186),
            .I(N__12183));
    Odrv4 I__1225 (
            .O(N__12183),
            .I(M_this_vga_signals_address_7));
    InMux I__1224 (
            .O(N__12180),
            .I(N__12177));
    LocalMux I__1223 (
            .O(N__12177),
            .I(\this_vga_signals.g1 ));
    InMux I__1222 (
            .O(N__12174),
            .I(N__12168));
    InMux I__1221 (
            .O(N__12173),
            .I(N__12168));
    LocalMux I__1220 (
            .O(N__12168),
            .I(N__12165));
    Odrv4 I__1219 (
            .O(N__12165),
            .I(\this_vga_signals.if_m2_0 ));
    InMux I__1218 (
            .O(N__12162),
            .I(N__12159));
    LocalMux I__1217 (
            .O(N__12159),
            .I(\this_vga_signals.if_m2_1 ));
    CascadeMux I__1216 (
            .O(N__12156),
            .I(\this_vga_signals.if_m2_1_cascade_ ));
    CascadeMux I__1215 (
            .O(N__12153),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ));
    InMux I__1214 (
            .O(N__12150),
            .I(N__12142));
    InMux I__1213 (
            .O(N__12149),
            .I(N__12137));
    InMux I__1212 (
            .O(N__12148),
            .I(N__12137));
    InMux I__1211 (
            .O(N__12147),
            .I(N__12134));
    InMux I__1210 (
            .O(N__12146),
            .I(N__12131));
    InMux I__1209 (
            .O(N__12145),
            .I(N__12128));
    LocalMux I__1208 (
            .O(N__12142),
            .I(N__12122));
    LocalMux I__1207 (
            .O(N__12137),
            .I(N__12119));
    LocalMux I__1206 (
            .O(N__12134),
            .I(N__12116));
    LocalMux I__1205 (
            .O(N__12131),
            .I(N__12113));
    LocalMux I__1204 (
            .O(N__12128),
            .I(N__12110));
    InMux I__1203 (
            .O(N__12127),
            .I(N__12107));
    InMux I__1202 (
            .O(N__12126),
            .I(N__12104));
    InMux I__1201 (
            .O(N__12125),
            .I(N__12101));
    Odrv12 I__1200 (
            .O(N__12122),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__1199 (
            .O(N__12119),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__1198 (
            .O(N__12116),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__1197 (
            .O(N__12113),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__1196 (
            .O(N__12110),
            .I(M_this_vga_ramdac_en_0));
    LocalMux I__1195 (
            .O(N__12107),
            .I(M_this_vga_ramdac_en_0));
    LocalMux I__1194 (
            .O(N__12104),
            .I(M_this_vga_ramdac_en_0));
    LocalMux I__1193 (
            .O(N__12101),
            .I(M_this_vga_ramdac_en_0));
    CascadeMux I__1192 (
            .O(N__12084),
            .I(N__12081));
    InMux I__1191 (
            .O(N__12081),
            .I(N__12078));
    LocalMux I__1190 (
            .O(N__12078),
            .I(N__12075));
    Span4Mux_h I__1189 (
            .O(N__12075),
            .I(N__12072));
    Span4Mux_v I__1188 (
            .O(N__12072),
            .I(N__12069));
    Odrv4 I__1187 (
            .O(N__12069),
            .I(M_this_vga_signals_address_2));
    InMux I__1186 (
            .O(N__12066),
            .I(N__12063));
    LocalMux I__1185 (
            .O(N__12063),
            .I(\this_vga_signals.g0_i_x4_0_4 ));
    InMux I__1184 (
            .O(N__12060),
            .I(N__12057));
    LocalMux I__1183 (
            .O(N__12057),
            .I(N__12054));
    Odrv12 I__1182 (
            .O(N__12054),
            .I(\this_vga_ramdac.m6 ));
    CascadeMux I__1181 (
            .O(N__12051),
            .I(G_463_cascade_));
    InMux I__1180 (
            .O(N__12048),
            .I(N__12045));
    LocalMux I__1179 (
            .O(N__12045),
            .I(N__12042));
    Span4Mux_v I__1178 (
            .O(N__12042),
            .I(N__12038));
    InMux I__1177 (
            .O(N__12041),
            .I(N__12035));
    Odrv4 I__1176 (
            .O(N__12038),
            .I(\this_vga_ramdac.N_2807_reto ));
    LocalMux I__1175 (
            .O(N__12035),
            .I(\this_vga_ramdac.N_2807_reto ));
    InMux I__1174 (
            .O(N__12030),
            .I(N__12024));
    InMux I__1173 (
            .O(N__12029),
            .I(N__12024));
    LocalMux I__1172 (
            .O(N__12024),
            .I(N_2_0));
    InMux I__1171 (
            .O(N__12021),
            .I(N__12018));
    LocalMux I__1170 (
            .O(N__12018),
            .I(M_this_vga_signals_pixel_clk_0_0));
    InMux I__1169 (
            .O(N__12015),
            .I(N__12005));
    InMux I__1168 (
            .O(N__12014),
            .I(N__12005));
    InMux I__1167 (
            .O(N__12013),
            .I(N__11996));
    InMux I__1166 (
            .O(N__12012),
            .I(N__11996));
    InMux I__1165 (
            .O(N__12011),
            .I(N__11996));
    InMux I__1164 (
            .O(N__12010),
            .I(N__11996));
    LocalMux I__1163 (
            .O(N__12005),
            .I(G_463));
    LocalMux I__1162 (
            .O(N__11996),
            .I(G_463));
    InMux I__1161 (
            .O(N__11991),
            .I(N__11988));
    LocalMux I__1160 (
            .O(N__11988),
            .I(N__11985));
    Odrv12 I__1159 (
            .O(N__11985),
            .I(\this_vga_ramdac.m19 ));
    InMux I__1158 (
            .O(N__11982),
            .I(N__11979));
    LocalMux I__1157 (
            .O(N__11979),
            .I(N__11976));
    Span4Mux_v I__1156 (
            .O(N__11976),
            .I(N__11972));
    CascadeMux I__1155 (
            .O(N__11975),
            .I(N__11969));
    Span4Mux_h I__1154 (
            .O(N__11972),
            .I(N__11966));
    InMux I__1153 (
            .O(N__11969),
            .I(N__11963));
    Odrv4 I__1152 (
            .O(N__11966),
            .I(\this_vga_ramdac.N_2810_reto ));
    LocalMux I__1151 (
            .O(N__11963),
            .I(\this_vga_ramdac.N_2810_reto ));
    InMux I__1150 (
            .O(N__11958),
            .I(N__11955));
    LocalMux I__1149 (
            .O(N__11955),
            .I(M_this_map_ram_write_data_0));
    InMux I__1148 (
            .O(N__11952),
            .I(N__11949));
    LocalMux I__1147 (
            .O(N__11949),
            .I(N__11946));
    Span4Mux_h I__1146 (
            .O(N__11946),
            .I(N__11943));
    Odrv4 I__1145 (
            .O(N__11943),
            .I(M_this_map_ram_write_data_5));
    InMux I__1144 (
            .O(N__11940),
            .I(N__11937));
    LocalMux I__1143 (
            .O(N__11937),
            .I(M_this_map_ram_write_data_6));
    CascadeMux I__1142 (
            .O(N__11934),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_ ));
    InMux I__1141 (
            .O(N__11931),
            .I(N__11927));
    InMux I__1140 (
            .O(N__11930),
            .I(N__11924));
    LocalMux I__1139 (
            .O(N__11927),
            .I(\this_vga_signals.mult1_un61_sum_axb1_2 ));
    LocalMux I__1138 (
            .O(N__11924),
            .I(\this_vga_signals.mult1_un61_sum_axb1_2 ));
    InMux I__1137 (
            .O(N__11919),
            .I(N__11916));
    LocalMux I__1136 (
            .O(N__11916),
            .I(N__11913));
    Odrv12 I__1135 (
            .O(N__11913),
            .I(\this_vga_ramdac.N_24_mux ));
    InMux I__1134 (
            .O(N__11910),
            .I(N__11906));
    CascadeMux I__1133 (
            .O(N__11909),
            .I(N__11903));
    LocalMux I__1132 (
            .O(N__11906),
            .I(N__11900));
    InMux I__1131 (
            .O(N__11903),
            .I(N__11897));
    Odrv12 I__1130 (
            .O(N__11900),
            .I(\this_vga_ramdac.N_2806_reto ));
    LocalMux I__1129 (
            .O(N__11897),
            .I(\this_vga_ramdac.N_2806_reto ));
    InMux I__1128 (
            .O(N__11892),
            .I(N__11886));
    InMux I__1127 (
            .O(N__11891),
            .I(N__11883));
    InMux I__1126 (
            .O(N__11890),
            .I(N__11878));
    InMux I__1125 (
            .O(N__11889),
            .I(N__11875));
    LocalMux I__1124 (
            .O(N__11886),
            .I(N__11870));
    LocalMux I__1123 (
            .O(N__11883),
            .I(N__11870));
    InMux I__1122 (
            .O(N__11882),
            .I(N__11867));
    InMux I__1121 (
            .O(N__11881),
            .I(N__11864));
    LocalMux I__1120 (
            .O(N__11878),
            .I(N__11858));
    LocalMux I__1119 (
            .O(N__11875),
            .I(N__11858));
    Span4Mux_v I__1118 (
            .O(N__11870),
            .I(N__11853));
    LocalMux I__1117 (
            .O(N__11867),
            .I(N__11853));
    LocalMux I__1116 (
            .O(N__11864),
            .I(N__11850));
    CascadeMux I__1115 (
            .O(N__11863),
            .I(N__11847));
    Span4Mux_v I__1114 (
            .O(N__11858),
            .I(N__11844));
    Span4Mux_h I__1113 (
            .O(N__11853),
            .I(N__11839));
    Span4Mux_v I__1112 (
            .O(N__11850),
            .I(N__11839));
    InMux I__1111 (
            .O(N__11847),
            .I(N__11836));
    Odrv4 I__1110 (
            .O(N__11844),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    Odrv4 I__1109 (
            .O(N__11839),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    LocalMux I__1108 (
            .O(N__11836),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    CascadeMux I__1107 (
            .O(N__11829),
            .I(\this_vga_signals.M_pcounter_q_3_0_cascade_ ));
    CascadeMux I__1106 (
            .O(N__11826),
            .I(N_2_0_cascade_));
    InMux I__1105 (
            .O(N__11823),
            .I(N__11820));
    LocalMux I__1104 (
            .O(N__11820),
            .I(N__11817));
    Span12Mux_v I__1103 (
            .O(N__11817),
            .I(N__11814));
    Odrv12 I__1102 (
            .O(N__11814),
            .I(\this_vga_ramdac.i2_mux_0 ));
    InMux I__1101 (
            .O(N__11811),
            .I(N__11808));
    LocalMux I__1100 (
            .O(N__11808),
            .I(N__11804));
    CascadeMux I__1099 (
            .O(N__11807),
            .I(N__11801));
    Span4Mux_v I__1098 (
            .O(N__11804),
            .I(N__11798));
    InMux I__1097 (
            .O(N__11801),
            .I(N__11795));
    Odrv4 I__1096 (
            .O(N__11798),
            .I(\this_vga_ramdac.N_2811_reto ));
    LocalMux I__1095 (
            .O(N__11795),
            .I(\this_vga_ramdac.N_2811_reto ));
    InMux I__1094 (
            .O(N__11790),
            .I(N__11787));
    LocalMux I__1093 (
            .O(N__11787),
            .I(N__11784));
    Span12Mux_v I__1092 (
            .O(N__11784),
            .I(N__11781));
    Odrv12 I__1091 (
            .O(N__11781),
            .I(\this_vga_ramdac.m16 ));
    InMux I__1090 (
            .O(N__11778),
            .I(N__11774));
    CascadeMux I__1089 (
            .O(N__11777),
            .I(N__11771));
    LocalMux I__1088 (
            .O(N__11774),
            .I(N__11768));
    InMux I__1087 (
            .O(N__11771),
            .I(N__11765));
    Odrv12 I__1086 (
            .O(N__11768),
            .I(\this_vga_ramdac.N_2809_reto ));
    LocalMux I__1085 (
            .O(N__11765),
            .I(\this_vga_ramdac.N_2809_reto ));
    InMux I__1084 (
            .O(N__11760),
            .I(N__11757));
    LocalMux I__1083 (
            .O(N__11757),
            .I(N__11754));
    Span4Mux_v I__1082 (
            .O(N__11754),
            .I(N__11751));
    Odrv4 I__1081 (
            .O(N__11751),
            .I(\this_vga_ramdac.i2_mux ));
    InMux I__1080 (
            .O(N__11748),
            .I(N__11745));
    LocalMux I__1079 (
            .O(N__11745),
            .I(N__11741));
    CascadeMux I__1078 (
            .O(N__11744),
            .I(N__11738));
    Span4Mux_h I__1077 (
            .O(N__11741),
            .I(N__11735));
    InMux I__1076 (
            .O(N__11738),
            .I(N__11732));
    Odrv4 I__1075 (
            .O(N__11735),
            .I(\this_vga_ramdac.N_2808_reto ));
    LocalMux I__1074 (
            .O(N__11732),
            .I(\this_vga_ramdac.N_2808_reto ));
    CascadeMux I__1073 (
            .O(N__11727),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_ ));
    InMux I__1072 (
            .O(N__11724),
            .I(N__11721));
    LocalMux I__1071 (
            .O(N__11721),
            .I(N__11718));
    Odrv4 I__1070 (
            .O(N__11718),
            .I(\this_vga_signals.g1_0_0 ));
    InMux I__1069 (
            .O(N__11715),
            .I(N__11712));
    LocalMux I__1068 (
            .O(N__11712),
            .I(\this_vga_signals.N_3_2_0_1 ));
    CascadeMux I__1067 (
            .O(N__11709),
            .I(\this_vga_signals.mult1_un61_sum_axb1_3_cascade_ ));
    InMux I__1066 (
            .O(N__11706),
            .I(N__11703));
    LocalMux I__1065 (
            .O(N__11703),
            .I(\this_vga_signals.g1_1 ));
    InMux I__1064 (
            .O(N__11700),
            .I(N__11697));
    LocalMux I__1063 (
            .O(N__11697),
            .I(\this_vga_signals.g0_0 ));
    CascadeMux I__1062 (
            .O(N__11694),
            .I(\this_vga_signals.g0_5_1_cascade_ ));
    InMux I__1061 (
            .O(N__11691),
            .I(N__11688));
    LocalMux I__1060 (
            .O(N__11688),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0_0_0_0 ));
    CascadeMux I__1059 (
            .O(N__11685),
            .I(N__11682));
    InMux I__1058 (
            .O(N__11682),
            .I(N__11679));
    LocalMux I__1057 (
            .O(N__11679),
            .I(N__11676));
    Odrv4 I__1056 (
            .O(N__11676),
            .I(\this_vga_signals.g1_0_0_0 ));
    CascadeMux I__1055 (
            .O(N__11673),
            .I(N__11670));
    InMux I__1054 (
            .O(N__11670),
            .I(N__11667));
    LocalMux I__1053 (
            .O(N__11667),
            .I(\this_vga_signals.g1_2_1 ));
    CascadeMux I__1052 (
            .O(N__11664),
            .I(\this_vga_signals.if_i4_mux_cascade_ ));
    CascadeMux I__1051 (
            .O(N__11661),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ));
    InMux I__1050 (
            .O(N__11658),
            .I(N__11655));
    LocalMux I__1049 (
            .O(N__11655),
            .I(\this_vga_signals.g1_0_2 ));
    InMux I__1048 (
            .O(N__11652),
            .I(N__11649));
    LocalMux I__1047 (
            .O(N__11649),
            .I(\this_vga_signals.g0_1 ));
    InMux I__1046 (
            .O(N__11646),
            .I(N__11643));
    LocalMux I__1045 (
            .O(N__11643),
            .I(\this_vga_signals.g1_4_0 ));
    CascadeMux I__1044 (
            .O(N__11640),
            .I(N__11637));
    InMux I__1043 (
            .O(N__11637),
            .I(N__11634));
    LocalMux I__1042 (
            .O(N__11634),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    CascadeMux I__1041 (
            .O(N__11631),
            .I(\this_vga_signals.g1_7_cascade_ ));
    CascadeMux I__1040 (
            .O(N__11628),
            .I(\this_vga_signals.N_6_0_cascade_ ));
    CascadeMux I__1039 (
            .O(N__11625),
            .I(N__11620));
    InMux I__1038 (
            .O(N__11624),
            .I(N__11616));
    InMux I__1037 (
            .O(N__11623),
            .I(N__11609));
    InMux I__1036 (
            .O(N__11620),
            .I(N__11609));
    InMux I__1035 (
            .O(N__11619),
            .I(N__11609));
    LocalMux I__1034 (
            .O(N__11616),
            .I(N__11606));
    LocalMux I__1033 (
            .O(N__11609),
            .I(N__11601));
    Span4Mux_h I__1032 (
            .O(N__11606),
            .I(N__11598));
    InMux I__1031 (
            .O(N__11605),
            .I(N__11593));
    InMux I__1030 (
            .O(N__11604),
            .I(N__11593));
    Span4Mux_h I__1029 (
            .O(N__11601),
            .I(N__11590));
    Odrv4 I__1028 (
            .O(N__11598),
            .I(M_this_vram_read_data_1));
    LocalMux I__1027 (
            .O(N__11593),
            .I(M_this_vram_read_data_1));
    Odrv4 I__1026 (
            .O(N__11590),
            .I(M_this_vram_read_data_1));
    CascadeMux I__1025 (
            .O(N__11583),
            .I(N__11576));
    CascadeMux I__1024 (
            .O(N__11582),
            .I(N__11572));
    InMux I__1023 (
            .O(N__11581),
            .I(N__11569));
    CascadeMux I__1022 (
            .O(N__11580),
            .I(N__11566));
    CascadeMux I__1021 (
            .O(N__11579),
            .I(N__11563));
    InMux I__1020 (
            .O(N__11576),
            .I(N__11556));
    InMux I__1019 (
            .O(N__11575),
            .I(N__11556));
    InMux I__1018 (
            .O(N__11572),
            .I(N__11556));
    LocalMux I__1017 (
            .O(N__11569),
            .I(N__11553));
    InMux I__1016 (
            .O(N__11566),
            .I(N__11548));
    InMux I__1015 (
            .O(N__11563),
            .I(N__11548));
    LocalMux I__1014 (
            .O(N__11556),
            .I(N__11545));
    Span4Mux_h I__1013 (
            .O(N__11553),
            .I(N__11542));
    LocalMux I__1012 (
            .O(N__11548),
            .I(M_this_vram_read_data_3));
    Odrv4 I__1011 (
            .O(N__11545),
            .I(M_this_vram_read_data_3));
    Odrv4 I__1010 (
            .O(N__11542),
            .I(M_this_vram_read_data_3));
    CascadeMux I__1009 (
            .O(N__11535),
            .I(\this_vga_signals.g1_1_0_0_0_cascade_ ));
    CascadeMux I__1008 (
            .O(N__11532),
            .I(\this_vga_signals.g1_0_1_0_0_cascade_ ));
    CascadeMux I__1007 (
            .O(N__11529),
            .I(N__11526));
    InMux I__1006 (
            .O(N__11526),
            .I(N__11523));
    LocalMux I__1005 (
            .O(N__11523),
            .I(N__11520));
    Span4Mux_v I__1004 (
            .O(N__11520),
            .I(N__11517));
    Odrv4 I__1003 (
            .O(N__11517),
            .I(M_this_vga_signals_address_0));
    InMux I__1002 (
            .O(N__11514),
            .I(N__11511));
    LocalMux I__1001 (
            .O(N__11511),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1_0 ));
    InMux I__1000 (
            .O(N__11508),
            .I(N__11505));
    LocalMux I__999 (
            .O(N__11505),
            .I(N__11502));
    Odrv12 I__998 (
            .O(N__11502),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1 ));
    CascadeMux I__997 (
            .O(N__11499),
            .I(N__11496));
    InMux I__996 (
            .O(N__11496),
            .I(N__11493));
    LocalMux I__995 (
            .O(N__11493),
            .I(N__11490));
    Span4Mux_v I__994 (
            .O(N__11490),
            .I(N__11487));
    Odrv4 I__993 (
            .O(N__11487),
            .I(M_this_vga_signals_address_3));
    CascadeMux I__992 (
            .O(N__11484),
            .I(\this_vga_signals.mult1_un61_sum_axb1_cascade_ ));
    CascadeMux I__991 (
            .O(N__11481),
            .I(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_cascade_));
    InMux I__990 (
            .O(N__11478),
            .I(N__11475));
    LocalMux I__989 (
            .O(N__11475),
            .I(N__11472));
    Odrv4 I__988 (
            .O(N__11472),
            .I(\this_vga_signals.if_i4_mux ));
    CascadeMux I__987 (
            .O(N__11469),
            .I(N__11466));
    InMux I__986 (
            .O(N__11466),
            .I(N__11463));
    LocalMux I__985 (
            .O(N__11463),
            .I(N__11460));
    Odrv4 I__984 (
            .O(N__11460),
            .I(M_this_vga_signals_address_1));
    CascadeMux I__983 (
            .O(N__11457),
            .I(N__11454));
    InMux I__982 (
            .O(N__11454),
            .I(N__11451));
    LocalMux I__981 (
            .O(N__11451),
            .I(N__11448));
    Span4Mux_v I__980 (
            .O(N__11448),
            .I(N__11445));
    Odrv4 I__979 (
            .O(N__11445),
            .I(M_this_vga_signals_address_6));
    InMux I__978 (
            .O(N__11442),
            .I(N__11439));
    LocalMux I__977 (
            .O(N__11439),
            .I(\this_vga_signals.mult1_un82_sum_c3 ));
    CascadeMux I__976 (
            .O(N__11436),
            .I(N__11433));
    InMux I__975 (
            .O(N__11433),
            .I(N__11430));
    LocalMux I__974 (
            .O(N__11430),
            .I(\this_vga_signals.N_219 ));
    InMux I__973 (
            .O(N__11427),
            .I(N__11418));
    InMux I__972 (
            .O(N__11426),
            .I(N__11418));
    InMux I__971 (
            .O(N__11425),
            .I(N__11418));
    LocalMux I__970 (
            .O(N__11418),
            .I(N__11415));
    Span4Mux_v I__969 (
            .O(N__11415),
            .I(N__11410));
    InMux I__968 (
            .O(N__11414),
            .I(N__11405));
    InMux I__967 (
            .O(N__11413),
            .I(N__11405));
    Odrv4 I__966 (
            .O(N__11410),
            .I(M_this_vram_read_data_2));
    LocalMux I__965 (
            .O(N__11405),
            .I(M_this_vram_read_data_2));
    InMux I__964 (
            .O(N__11400),
            .I(N__11392));
    InMux I__963 (
            .O(N__11399),
            .I(N__11385));
    InMux I__962 (
            .O(N__11398),
            .I(N__11385));
    InMux I__961 (
            .O(N__11397),
            .I(N__11385));
    InMux I__960 (
            .O(N__11396),
            .I(N__11380));
    InMux I__959 (
            .O(N__11395),
            .I(N__11380));
    LocalMux I__958 (
            .O(N__11392),
            .I(N__11375));
    LocalMux I__957 (
            .O(N__11385),
            .I(N__11375));
    LocalMux I__956 (
            .O(N__11380),
            .I(M_this_vram_read_data_0));
    Odrv4 I__955 (
            .O(N__11375),
            .I(M_this_vram_read_data_0));
    CascadeMux I__954 (
            .O(N__11370),
            .I(N__11367));
    CascadeBuf I__953 (
            .O(N__11367),
            .I(N__11364));
    CascadeMux I__952 (
            .O(N__11364),
            .I(N__11361));
    InMux I__951 (
            .O(N__11361),
            .I(N__11358));
    LocalMux I__950 (
            .O(N__11358),
            .I(N__11354));
    InMux I__949 (
            .O(N__11357),
            .I(N__11351));
    Span4Mux_v I__948 (
            .O(N__11354),
            .I(N__11348));
    LocalMux I__947 (
            .O(N__11351),
            .I(M_this_map_address_qZ0Z_4));
    Odrv4 I__946 (
            .O(N__11348),
            .I(M_this_map_address_qZ0Z_4));
    InMux I__945 (
            .O(N__11343),
            .I(un1_M_this_map_address_q_cry_3));
    CascadeMux I__944 (
            .O(N__11340),
            .I(N__11337));
    CascadeBuf I__943 (
            .O(N__11337),
            .I(N__11334));
    CascadeMux I__942 (
            .O(N__11334),
            .I(N__11331));
    InMux I__941 (
            .O(N__11331),
            .I(N__11328));
    LocalMux I__940 (
            .O(N__11328),
            .I(N__11324));
    InMux I__939 (
            .O(N__11327),
            .I(N__11321));
    Span4Mux_v I__938 (
            .O(N__11324),
            .I(N__11318));
    LocalMux I__937 (
            .O(N__11321),
            .I(M_this_map_address_qZ0Z_5));
    Odrv4 I__936 (
            .O(N__11318),
            .I(M_this_map_address_qZ0Z_5));
    InMux I__935 (
            .O(N__11313),
            .I(un1_M_this_map_address_q_cry_4));
    CascadeMux I__934 (
            .O(N__11310),
            .I(N__11307));
    CascadeBuf I__933 (
            .O(N__11307),
            .I(N__11304));
    CascadeMux I__932 (
            .O(N__11304),
            .I(N__11301));
    InMux I__931 (
            .O(N__11301),
            .I(N__11298));
    LocalMux I__930 (
            .O(N__11298),
            .I(N__11294));
    InMux I__929 (
            .O(N__11297),
            .I(N__11291));
    Span4Mux_v I__928 (
            .O(N__11294),
            .I(N__11288));
    LocalMux I__927 (
            .O(N__11291),
            .I(M_this_map_address_qZ0Z_6));
    Odrv4 I__926 (
            .O(N__11288),
            .I(M_this_map_address_qZ0Z_6));
    InMux I__925 (
            .O(N__11283),
            .I(un1_M_this_map_address_q_cry_5));
    CascadeMux I__924 (
            .O(N__11280),
            .I(N__11277));
    CascadeBuf I__923 (
            .O(N__11277),
            .I(N__11274));
    CascadeMux I__922 (
            .O(N__11274),
            .I(N__11271));
    InMux I__921 (
            .O(N__11271),
            .I(N__11268));
    LocalMux I__920 (
            .O(N__11268),
            .I(N__11264));
    InMux I__919 (
            .O(N__11267),
            .I(N__11261));
    Span4Mux_v I__918 (
            .O(N__11264),
            .I(N__11258));
    LocalMux I__917 (
            .O(N__11261),
            .I(M_this_map_address_qZ0Z_7));
    Odrv4 I__916 (
            .O(N__11258),
            .I(M_this_map_address_qZ0Z_7));
    InMux I__915 (
            .O(N__11253),
            .I(un1_M_this_map_address_q_cry_6));
    CascadeMux I__914 (
            .O(N__11250),
            .I(N__11247));
    CascadeBuf I__913 (
            .O(N__11247),
            .I(N__11244));
    CascadeMux I__912 (
            .O(N__11244),
            .I(N__11241));
    InMux I__911 (
            .O(N__11241),
            .I(N__11238));
    LocalMux I__910 (
            .O(N__11238),
            .I(N__11234));
    InMux I__909 (
            .O(N__11237),
            .I(N__11231));
    Span4Mux_v I__908 (
            .O(N__11234),
            .I(N__11228));
    LocalMux I__907 (
            .O(N__11231),
            .I(M_this_map_address_qZ0Z_8));
    Odrv4 I__906 (
            .O(N__11228),
            .I(M_this_map_address_qZ0Z_8));
    InMux I__905 (
            .O(N__11223),
            .I(bfn_7_25_0_));
    InMux I__904 (
            .O(N__11220),
            .I(un1_M_this_map_address_q_cry_8));
    CascadeMux I__903 (
            .O(N__11217),
            .I(N__11214));
    CascadeBuf I__902 (
            .O(N__11214),
            .I(N__11211));
    CascadeMux I__901 (
            .O(N__11211),
            .I(N__11208));
    InMux I__900 (
            .O(N__11208),
            .I(N__11205));
    LocalMux I__899 (
            .O(N__11205),
            .I(N__11201));
    InMux I__898 (
            .O(N__11204),
            .I(N__11198));
    Span4Mux_v I__897 (
            .O(N__11201),
            .I(N__11195));
    LocalMux I__896 (
            .O(N__11198),
            .I(M_this_map_address_qZ0Z_9));
    Odrv4 I__895 (
            .O(N__11195),
            .I(M_this_map_address_qZ0Z_9));
    CascadeMux I__894 (
            .O(N__11190),
            .I(N__11187));
    InMux I__893 (
            .O(N__11187),
            .I(N__11184));
    LocalMux I__892 (
            .O(N__11184),
            .I(M_this_vga_signals_address_5));
    CascadeMux I__891 (
            .O(N__11181),
            .I(N__11178));
    InMux I__890 (
            .O(N__11178),
            .I(N__11175));
    LocalMux I__889 (
            .O(N__11175),
            .I(M_this_vga_signals_address_4));
    IoInMux I__888 (
            .O(N__11172),
            .I(N__11169));
    LocalMux I__887 (
            .O(N__11169),
            .I(N__11166));
    Span4Mux_s2_h I__886 (
            .O(N__11166),
            .I(N__11163));
    Sp12to4 I__885 (
            .O(N__11163),
            .I(N__11160));
    Span12Mux_v I__884 (
            .O(N__11160),
            .I(N__11157));
    Odrv12 I__883 (
            .O(N__11157),
            .I(rgb_c_3));
    IoInMux I__882 (
            .O(N__11154),
            .I(N__11151));
    LocalMux I__881 (
            .O(N__11151),
            .I(N__11148));
    Odrv12 I__880 (
            .O(N__11148),
            .I(this_vga_signals_vvisibility_i));
    IoInMux I__879 (
            .O(N__11145),
            .I(N__11142));
    LocalMux I__878 (
            .O(N__11142),
            .I(N__11139));
    IoSpan4Mux I__877 (
            .O(N__11139),
            .I(N__11136));
    Span4Mux_s3_h I__876 (
            .O(N__11136),
            .I(N__11133));
    Sp12to4 I__875 (
            .O(N__11133),
            .I(N__11130));
    Span12Mux_v I__874 (
            .O(N__11130),
            .I(N__11127));
    Odrv12 I__873 (
            .O(N__11127),
            .I(rgb_c_5));
    IoInMux I__872 (
            .O(N__11124),
            .I(N__11121));
    LocalMux I__871 (
            .O(N__11121),
            .I(N__11118));
    IoSpan4Mux I__870 (
            .O(N__11118),
            .I(N__11115));
    Span4Mux_s3_h I__869 (
            .O(N__11115),
            .I(N__11112));
    Odrv4 I__868 (
            .O(N__11112),
            .I(rgb_c_1));
    CascadeMux I__867 (
            .O(N__11109),
            .I(N__11106));
    CascadeBuf I__866 (
            .O(N__11106),
            .I(N__11103));
    CascadeMux I__865 (
            .O(N__11103),
            .I(N__11100));
    InMux I__864 (
            .O(N__11100),
            .I(N__11097));
    LocalMux I__863 (
            .O(N__11097),
            .I(N__11093));
    InMux I__862 (
            .O(N__11096),
            .I(N__11090));
    Span4Mux_v I__861 (
            .O(N__11093),
            .I(N__11087));
    LocalMux I__860 (
            .O(N__11090),
            .I(M_this_map_address_qZ0Z_0));
    Odrv4 I__859 (
            .O(N__11087),
            .I(M_this_map_address_qZ0Z_0));
    CascadeMux I__858 (
            .O(N__11082),
            .I(N__11079));
    CascadeBuf I__857 (
            .O(N__11079),
            .I(N__11076));
    CascadeMux I__856 (
            .O(N__11076),
            .I(N__11073));
    InMux I__855 (
            .O(N__11073),
            .I(N__11070));
    LocalMux I__854 (
            .O(N__11070),
            .I(N__11066));
    InMux I__853 (
            .O(N__11069),
            .I(N__11063));
    Span4Mux_v I__852 (
            .O(N__11066),
            .I(N__11060));
    LocalMux I__851 (
            .O(N__11063),
            .I(M_this_map_address_qZ0Z_1));
    Odrv4 I__850 (
            .O(N__11060),
            .I(M_this_map_address_qZ0Z_1));
    InMux I__849 (
            .O(N__11055),
            .I(un1_M_this_map_address_q_cry_0));
    CascadeMux I__848 (
            .O(N__11052),
            .I(N__11049));
    CascadeBuf I__847 (
            .O(N__11049),
            .I(N__11046));
    CascadeMux I__846 (
            .O(N__11046),
            .I(N__11043));
    InMux I__845 (
            .O(N__11043),
            .I(N__11040));
    LocalMux I__844 (
            .O(N__11040),
            .I(N__11036));
    InMux I__843 (
            .O(N__11039),
            .I(N__11033));
    Span4Mux_v I__842 (
            .O(N__11036),
            .I(N__11030));
    LocalMux I__841 (
            .O(N__11033),
            .I(M_this_map_address_qZ0Z_2));
    Odrv4 I__840 (
            .O(N__11030),
            .I(M_this_map_address_qZ0Z_2));
    InMux I__839 (
            .O(N__11025),
            .I(un1_M_this_map_address_q_cry_1));
    CascadeMux I__838 (
            .O(N__11022),
            .I(N__11019));
    CascadeBuf I__837 (
            .O(N__11019),
            .I(N__11016));
    CascadeMux I__836 (
            .O(N__11016),
            .I(N__11013));
    InMux I__835 (
            .O(N__11013),
            .I(N__11010));
    LocalMux I__834 (
            .O(N__11010),
            .I(N__11006));
    InMux I__833 (
            .O(N__11009),
            .I(N__11003));
    Span4Mux_v I__832 (
            .O(N__11006),
            .I(N__11000));
    LocalMux I__831 (
            .O(N__11003),
            .I(M_this_map_address_qZ0Z_3));
    Odrv4 I__830 (
            .O(N__11000),
            .I(M_this_map_address_qZ0Z_3));
    InMux I__829 (
            .O(N__10995),
            .I(un1_M_this_map_address_q_cry_2));
    IoInMux I__828 (
            .O(N__10992),
            .I(N__10989));
    LocalMux I__827 (
            .O(N__10989),
            .I(N__10986));
    Span4Mux_s0_h I__826 (
            .O(N__10986),
            .I(N__10983));
    Sp12to4 I__825 (
            .O(N__10983),
            .I(N__10980));
    Odrv12 I__824 (
            .O(N__10980),
            .I(port_data_rw_0_i));
    IoInMux I__823 (
            .O(N__10977),
            .I(N__10974));
    LocalMux I__822 (
            .O(N__10974),
            .I(N__10971));
    Span4Mux_s3_h I__821 (
            .O(N__10971),
            .I(N__10968));
    Sp12to4 I__820 (
            .O(N__10968),
            .I(N__10965));
    Odrv12 I__819 (
            .O(N__10965),
            .I(rgb_c_0));
    IoInMux I__818 (
            .O(N__10962),
            .I(N__10959));
    LocalMux I__817 (
            .O(N__10959),
            .I(N__10956));
    Span4Mux_s3_h I__816 (
            .O(N__10956),
            .I(N__10953));
    Odrv4 I__815 (
            .O(N__10953),
            .I(rgb_c_2));
    IoInMux I__814 (
            .O(N__10950),
            .I(N__10947));
    LocalMux I__813 (
            .O(N__10947),
            .I(N__10944));
    Span4Mux_s3_h I__812 (
            .O(N__10944),
            .I(N__10941));
    Span4Mux_v I__811 (
            .O(N__10941),
            .I(N__10938));
    Sp12to4 I__810 (
            .O(N__10938),
            .I(N__10935));
    Odrv12 I__809 (
            .O(N__10935),
            .I(rgb_c_4));
    IoInMux I__808 (
            .O(N__10932),
            .I(N__10929));
    LocalMux I__807 (
            .O(N__10929),
            .I(N__10926));
    Odrv12 I__806 (
            .O(N__10926),
            .I(port_nmib_0_i));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_20_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_19_0_));
    defparam IN_MUX_bfv_20_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_20_0_ (
            .carryinitin(\this_ppu.un1_M_vaddress_q_cry_7 ),
            .carryinitout(bfn_20_20_0_));
    defparam IN_MUX_bfv_19_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_19_0_));
    defparam IN_MUX_bfv_19_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_20_0_ (
            .carryinitin(\this_ppu.un1_M_haddress_q_cry_7 ),
            .carryinitout(bfn_19_20_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(M_this_data_count_q_cry_7),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_24_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_16_0_));
    defparam IN_MUX_bfv_24_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_19_0_));
    defparam IN_MUX_bfv_19_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_17_0_));
    defparam IN_MUX_bfv_19_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_18_0_ (
            .carryinitin(\this_ppu.un1_M_vaddress_q_3_cry_7 ),
            .carryinitout(bfn_19_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\this_ppu.un1_M_haddress_q_2_cry_7 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_28_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_28_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_28_21_0_));
    defparam IN_MUX_bfv_28_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_28_22_0_ (
            .carryinitin(un1_M_this_external_address_q_cry_7),
            .carryinitout(bfn_28_22_0_));
    defparam IN_MUX_bfv_21_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_13_0_));
    defparam IN_MUX_bfv_21_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_14_0_ (
            .carryinitin(un1_M_this_sprites_address_q_cry_7),
            .carryinitout(bfn_21_14_0_));
    defparam IN_MUX_bfv_7_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_24_0_));
    defparam IN_MUX_bfv_7_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_25_0_ (
            .carryinitin(un1_M_this_map_address_q_cry_7),
            .carryinitout(bfn_7_25_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNI67JU6_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__17160),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_1098_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_9  (
            .USERSIGNALTOGLOBALBUFFER(N__34657),
            .GLOBALBUFFEROUTPUT(M_this_reset_cond_out_g_0));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__17316),
            .GLOBALBUFFEROUTPUT(N_515_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_ppu.port_data_rw_0_i_LC_1_20_3 .C_ON=1'b0;
    defparam \this_ppu.port_data_rw_0_i_LC_1_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.port_data_rw_0_i_LC_1_20_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \this_ppu.port_data_rw_0_i_LC_1_20_3  (
            .in0(N__21404),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26567),
            .lcout(port_data_rw_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_4_14_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_4_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(N__11910),
            .in2(_gnd_net_),
            .in3(N__11882),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_15_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_15_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_15_1  (
            .in0(N__11891),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11748),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_16_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_16_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_16_3  (
            .in0(N__11892),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11982),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI497S8_9_LC_5_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI497S8_9_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI497S8_9_LC_5_11_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI497S8_9_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__21408),
            .in2(_gnd_net_),
            .in3(N__15326),
            .lcout(port_nmib_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_5_15_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_5_15_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_5_15_6  (
            .in0(N__11778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11889),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_27_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_27_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_27_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM8094_0_9_LC_5_29_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM8094_0_9_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM8094_0_9_LC_5_29_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIM8094_0_9_LC_5_29_3  (
            .in0(N__15327),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_vvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_6_16_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_6_16_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_6_16_6  (
            .in0(N__11811),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11890),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_16_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__11881),
            .in2(_gnd_net_),
            .in3(N__12048),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_0_LC_7_24_0.C_ON=1'b1;
    defparam M_this_map_address_q_0_LC_7_24_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_0_LC_7_24_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_0_LC_7_24_0 (
            .in0(N__17574),
            .in1(N__11096),
            .in2(N__17433),
            .in3(N__17436),
            .lcout(M_this_map_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_7_24_0_),
            .carryout(un1_M_this_map_address_q_cry_0),
            .clk(N__34632),
            .ce(),
            .sr(N__28662));
    defparam M_this_map_address_q_1_LC_7_24_1.C_ON=1'b1;
    defparam M_this_map_address_q_1_LC_7_24_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_1_LC_7_24_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_1_LC_7_24_1 (
            .in0(N__17578),
            .in1(N__11069),
            .in2(_gnd_net_),
            .in3(N__11055),
            .lcout(M_this_map_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_0),
            .carryout(un1_M_this_map_address_q_cry_1),
            .clk(N__34632),
            .ce(),
            .sr(N__28662));
    defparam M_this_map_address_q_2_LC_7_24_2.C_ON=1'b1;
    defparam M_this_map_address_q_2_LC_7_24_2.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_2_LC_7_24_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_2_LC_7_24_2 (
            .in0(N__17575),
            .in1(N__11039),
            .in2(_gnd_net_),
            .in3(N__11025),
            .lcout(M_this_map_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_1),
            .carryout(un1_M_this_map_address_q_cry_2),
            .clk(N__34632),
            .ce(),
            .sr(N__28662));
    defparam M_this_map_address_q_3_LC_7_24_3.C_ON=1'b1;
    defparam M_this_map_address_q_3_LC_7_24_3.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_3_LC_7_24_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_3_LC_7_24_3 (
            .in0(N__17579),
            .in1(N__11009),
            .in2(_gnd_net_),
            .in3(N__10995),
            .lcout(M_this_map_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_2),
            .carryout(un1_M_this_map_address_q_cry_3),
            .clk(N__34632),
            .ce(),
            .sr(N__28662));
    defparam M_this_map_address_q_4_LC_7_24_4.C_ON=1'b1;
    defparam M_this_map_address_q_4_LC_7_24_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_4_LC_7_24_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_4_LC_7_24_4 (
            .in0(N__17576),
            .in1(N__11357),
            .in2(_gnd_net_),
            .in3(N__11343),
            .lcout(M_this_map_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_3),
            .carryout(un1_M_this_map_address_q_cry_4),
            .clk(N__34632),
            .ce(),
            .sr(N__28662));
    defparam M_this_map_address_q_5_LC_7_24_5.C_ON=1'b1;
    defparam M_this_map_address_q_5_LC_7_24_5.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_5_LC_7_24_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_5_LC_7_24_5 (
            .in0(N__17580),
            .in1(N__11327),
            .in2(_gnd_net_),
            .in3(N__11313),
            .lcout(M_this_map_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_4),
            .carryout(un1_M_this_map_address_q_cry_5),
            .clk(N__34632),
            .ce(),
            .sr(N__28662));
    defparam M_this_map_address_q_6_LC_7_24_6.C_ON=1'b1;
    defparam M_this_map_address_q_6_LC_7_24_6.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_6_LC_7_24_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_6_LC_7_24_6 (
            .in0(N__17577),
            .in1(N__11297),
            .in2(_gnd_net_),
            .in3(N__11283),
            .lcout(M_this_map_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_5),
            .carryout(un1_M_this_map_address_q_cry_6),
            .clk(N__34632),
            .ce(),
            .sr(N__28662));
    defparam M_this_map_address_q_7_LC_7_24_7.C_ON=1'b1;
    defparam M_this_map_address_q_7_LC_7_24_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_7_LC_7_24_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_7_LC_7_24_7 (
            .in0(N__17581),
            .in1(N__11267),
            .in2(_gnd_net_),
            .in3(N__11253),
            .lcout(M_this_map_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_6),
            .carryout(un1_M_this_map_address_q_cry_7),
            .clk(N__34632),
            .ce(),
            .sr(N__28662));
    defparam M_this_map_address_q_8_LC_7_25_0.C_ON=1'b1;
    defparam M_this_map_address_q_8_LC_7_25_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_8_LC_7_25_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_8_LC_7_25_0 (
            .in0(N__17582),
            .in1(N__11237),
            .in2(_gnd_net_),
            .in3(N__11223),
            .lcout(M_this_map_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_7_25_0_),
            .carryout(un1_M_this_map_address_q_cry_8),
            .clk(N__34639),
            .ce(),
            .sr(N__28659));
    defparam M_this_map_address_q_9_LC_7_25_1.C_ON=1'b0;
    defparam M_this_map_address_q_9_LC_7_25_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_9_LC_7_25_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_map_address_q_9_LC_7_25_1 (
            .in0(N__11204),
            .in1(N__17583),
            .in2(_gnd_net_),
            .in3(N__11220),
            .lcout(M_this_map_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34639),
            .ce(),
            .sr(N__28659));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3J5O7_9_LC_9_6_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3J5O7_9_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3J5O7_9_LC_9_6_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3J5O7_9_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__12148),
            .in2(_gnd_net_),
            .in3(N__12831),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI7VUTC_9_LC_9_6_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI7VUTC_9_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI7VUTC_9_LC_9_6_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI7VUTC_9_LC_9_6_7  (
            .in0(N__12149),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12677),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_7_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_7_1 .LUT_INIT=16'b0110001101001101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_7_1  (
            .in0(N__11605),
            .in1(N__11414),
            .in2(N__11580),
            .in3(N__11396),
            .lcout(\this_vga_ramdac.m19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_7_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_7_3 .LUT_INIT=16'b0100010110010111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_7_3  (
            .in0(N__11604),
            .in1(N__11413),
            .in2(N__11579),
            .in3(N__11395),
            .lcout(\this_vga_ramdac.m16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIEDCEO4_9_LC_9_7_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIEDCEO4_9_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIEDCEO4_9_LC_9_7_4 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIEDCEO4_9_LC_9_7_4  (
            .in0(N__12146),
            .in1(N__11508),
            .in2(_gnd_net_),
            .in3(N__11442),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_8_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_8_1 .LUT_INIT=16'b0101010100100010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_8_1  (
            .in0(N__11581),
            .in1(N__11624),
            .in2(_gnd_net_),
            .in3(N__11400),
            .lcout(\this_vga_ramdac.N_24_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIF2OJ6_6_LC_9_8_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIF2OJ6_6_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIF2OJ6_6_LC_9_8_5 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIF2OJ6_6_LC_9_8_5  (
            .in0(N__12126),
            .in1(N__14469),
            .in2(N__11436),
            .in3(N__12474),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_9_8_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_9_8_6 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_9_8_6  (
            .in0(N__11478),
            .in1(N__12315),
            .in2(N__12360),
            .in3(N__12423),
            .lcout(\this_vga_signals.mult1_un82_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_9_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_9_0 .LUT_INIT=16'b0011001000111111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_9_0  (
            .in0(N__11399),
            .in1(N__11427),
            .in2(N__11583),
            .in3(N__11623),
            .lcout(\this_vga_ramdac.m6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_9_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_9_9_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_9_9_1  (
            .in0(N__13668),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13581),
            .lcout(\this_vga_signals.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIKHT15_9_LC_9_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIKHT15_9_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIKHT15_9_LC_9_9_3 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIKHT15_9_LC_9_9_3  (
            .in0(N__13667),
            .in1(N__13580),
            .in2(N__15325),
            .in3(N__13890),
            .lcout(M_this_vga_ramdac_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_9_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_9_4 .LUT_INIT=16'b0010001101001011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_9_4  (
            .in0(N__11397),
            .in1(N__11426),
            .in2(N__11582),
            .in3(N__11619),
            .lcout(\this_vga_ramdac.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_9_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_9_5 .LUT_INIT=16'b0000011101110101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_9_5  (
            .in0(N__11425),
            .in1(N__11398),
            .in2(N__11625),
            .in3(N__11575),
            .lcout(\this_vga_ramdac.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_18_LC_9_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_18_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_18_LC_9_10_0 .LUT_INIT=16'b1011100010001011;
    LogicCell40 \this_vga_signals.un4_haddress_g0_18_LC_9_10_0  (
            .in0(N__14961),
            .in1(N__12162),
            .in2(N__11685),
            .in3(N__12678),
            .lcout(),
            .ltout(\this_vga_signals.g1_1_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNITO6PD6_2_LC_9_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNITO6PD6_2_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNITO6PD6_2_LC_9_10_1 .LUT_INIT=16'b1110101110000010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNITO6PD6_2_LC_9_10_1  (
            .in0(N__14958),
            .in1(N__12396),
            .in2(N__11535),
            .in3(N__12246),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIAQLVLB_2_LC_9_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIAQLVLB_2_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIAQLVLB_2_LC_9_10_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIAQLVLB_2_LC_9_10_2  (
            .in0(N__12125),
            .in1(N__11514),
            .in2(N__11532),
            .in3(N__11658),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_16_LC_9_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_16_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_16_LC_9_10_3 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \this_vga_signals.un4_haddress_g0_16_LC_9_10_3  (
            .in0(N__12174),
            .in1(N__14965),
            .in2(N__12333),
            .in3(N__12353),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_9_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_9_10_6 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_9_10_6  (
            .in0(N__12352),
            .in1(N__12328),
            .in2(N__14967),
            .in3(N__12173),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG45VS_9_LC_9_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG45VS_9_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG45VS_9_LC_9_10_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIG45VS_9_LC_9_10_7  (
            .in0(N__12145),
            .in1(N__12295),
            .in2(_gnd_net_),
            .in3(N__12240),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_9_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_9_11_0 .LUT_INIT=16'b1100000110000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_9_11_0  (
            .in0(N__13052),
            .in1(N__12980),
            .in2(N__14296),
            .in3(N__14462),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_9_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_9_11_1 .LUT_INIT=16'b1100011111000001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_9_11_1  (
            .in0(N__13794),
            .in1(N__14123),
            .in2(N__11484),
            .in3(N__12652),
            .lcout(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0),
            .ltout(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m4_LC_9_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m4_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m4_LC_9_11_2 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \this_vga_signals.un4_haddress_if_m4_LC_9_11_2  (
            .in0(N__14865),
            .in1(N__13797),
            .in2(N__11481),
            .in3(N__12293),
            .lcout(\this_vga_signals.if_i4_mux ),
            .ltout(\this_vga_signals.if_i4_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_1_LC_9_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_1_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_1_LC_9_11_3 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \this_vga_signals.un4_haddress_g0_1_LC_9_11_3  (
            .in0(N__12294),
            .in1(N__11706),
            .in2(N__11664),
            .in3(N__11652),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIQSM9K2_2_LC_9_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIQSM9K2_2_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIQSM9K2_2_LC_9_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIQSM9K2_2_LC_9_11_4  (
            .in0(N__11724),
            .in1(N__12594),
            .in2(N__11661),
            .in3(N__11646),
            .lcout(\this_vga_signals.g1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIAJMMB_2_LC_9_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIAJMMB_2_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIAJMMB_2_LC_9_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIAJMMB_2_LC_9_11_5  (
            .in0(N__13796),
            .in1(N__14957),
            .in2(_gnd_net_),
            .in3(N__12235),
            .lcout(\this_vga_signals.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI2BF2A_2_LC_9_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI2BF2A_2_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI2BF2A_2_LC_9_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI2BF2A_2_LC_9_11_6  (
            .in0(N__12654),
            .in1(N__12435),
            .in2(_gnd_net_),
            .in3(N__12585),
            .lcout(\this_vga_signals.g1_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_11_7 .LUT_INIT=16'b1000011111100001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_11_7  (
            .in0(N__13795),
            .in1(N__14124),
            .in2(N__11640),
            .in3(N__12653),
            .lcout(this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_7_LC_9_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_7_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_7_LC_9_12_0 .LUT_INIT=16'b0101111100000101;
    LogicCell40 \this_vga_signals.un4_haddress_g1_7_LC_9_12_0  (
            .in0(N__13786),
            .in1(_gnd_net_),
            .in2(N__14138),
            .in3(N__12646),
            .lcout(\this_vga_signals.g1_7 ),
            .ltout(\this_vga_signals.g1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_7_LC_9_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_7_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_7_LC_9_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_haddress_g0_7_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__14956),
            .in2(N__11631),
            .in3(N__11930),
            .lcout(),
            .ltout(\this_vga_signals.N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_m2_LC_9_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_m2_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_m2_LC_9_12_2 .LUT_INIT=16'b1011111100000100;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_m2_LC_9_12_2  (
            .in0(N__11715),
            .in1(N__12372),
            .in2(N__11628),
            .in3(N__11691),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_4_LC_9_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_4_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_4_LC_9_12_3 .LUT_INIT=16'b0100101011011010;
    LogicCell40 \this_vga_signals.un4_haddress_g0_4_LC_9_12_3  (
            .in0(N__14465),
            .in1(N__12584),
            .in2(N__11673),
            .in3(N__14293),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_10_LC_9_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_10_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_10_LC_9_12_4 .LUT_INIT=16'b1111101001011111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_10_LC_9_12_4  (
            .in0(N__14294),
            .in1(_gnd_net_),
            .in2(N__11727),
            .in3(N__14133),
            .lcout(\this_vga_signals.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_20_LC_9_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_20_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_20_LC_9_12_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_haddress_g0_20_LC_9_12_5  (
            .in0(N__12647),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14128),
            .lcout(\this_vga_signals.N_3_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_2_LC_9_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_2_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_2_LC_9_12_6 .LUT_INIT=16'b1100000110000011;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_2_LC_9_12_6  (
            .in0(N__13049),
            .in1(N__12979),
            .in2(N__14298),
            .in3(N__14464),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axb1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_0_LC_9_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_0_LC_9_12_7 .LUT_INIT=16'b1011010000101101;
    LogicCell40 \this_vga_signals.un4_haddress_g1_0_LC_9_12_7  (
            .in0(N__12648),
            .in1(N__14132),
            .in2(N__11709),
            .in3(N__13787),
            .lcout(\this_vga_signals.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_6_LC_9_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_6_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_6_LC_9_13_0 .LUT_INIT=16'b1111011111101111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_6_LC_9_13_0  (
            .in0(N__14088),
            .in1(N__14270),
            .in2(N__12453),
            .in3(N__12973),
            .lcout(\this_vga_signals.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_5_1_LC_9_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_5_1_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_5_1_LC_9_13_2 .LUT_INIT=16'b0010001001000100;
    LogicCell40 \this_vga_signals.un4_haddress_g0_5_1_LC_9_13_2  (
            .in0(N__14089),
            .in1(N__13767),
            .in2(_gnd_net_),
            .in3(N__12649),
            .lcout(),
            .ltout(\this_vga_signals.g0_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_5_LC_9_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_5_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_5_LC_9_13_3 .LUT_INIT=16'b0011100111000110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_5_LC_9_13_3  (
            .in0(N__11931),
            .in1(N__11700),
            .in2(N__11694),
            .in3(N__12504),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_0_0_LC_9_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_0_0_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_0_0_LC_9_13_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_haddress_g1_0_0_LC_9_13_4  (
            .in0(N__14090),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13768),
            .lcout(\this_vga_signals.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_1_9_LC_9_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_1_9_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_1_9_LC_9_13_5 .LUT_INIT=16'b1101110110111011;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_1_9_LC_9_13_5  (
            .in0(N__13660),
            .in1(N__13564),
            .in2(_gnd_net_),
            .in3(N__13880),
            .lcout(\this_vga_signals.g1_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_1_LC_9_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_1_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_1_LC_9_13_6 .LUT_INIT=16'b1100000110000011;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_1_LC_9_13_6  (
            .in0(N__13045),
            .in1(N__12974),
            .in2(N__14289),
            .in3(N__14450),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_14_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_14_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_14_1  (
            .in0(N__11919),
            .in1(N__34733),
            .in2(N__11909),
            .in3(N__12014),
            .lcout(\this_vga_ramdac.N_2806_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34594),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_14_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_14_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_ret_LC_9_14_2  (
            .in0(N__12015),
            .in1(N__34734),
            .in2(N__11863),
            .in3(N__12150),
            .lcout(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34594),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_9_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_9_14_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_9_14_5  (
            .in0(N__13092),
            .in1(N__12569),
            .in2(_gnd_net_),
            .in3(N__17071),
            .lcout(),
            .ltout(\this_vga_signals.M_pcounter_q_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_9_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_9_14_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__13150),
            .in2(N__11829),
            .in3(N__17310),
            .lcout(N_2_0),
            .ltout(N_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_9_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_9_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11826),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_pcounter_q_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34594),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_15_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_15_0 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_15_0  (
            .in0(N__34726),
            .in1(N__11823),
            .in2(N__11807),
            .in3(N__12013),
            .lcout(\this_vga_ramdac.N_2811_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34601),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_15_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_15_1 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_15_1  (
            .in0(N__12011),
            .in1(N__11790),
            .in2(N__11777),
            .in3(N__34724),
            .lcout(\this_vga_ramdac.N_2809_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34601),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_15_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_15_2 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_15_2  (
            .in0(N__34723),
            .in1(N__11760),
            .in2(N__11744),
            .in3(N__12010),
            .lcout(\this_vga_ramdac.N_2808_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34601),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.G_463_LC_9_15_4 .C_ON=1'b0;
    defparam \this_ppu.G_463_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.G_463_LC_9_15_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.G_463_LC_9_15_4  (
            .in0(N__12021),
            .in1(N__13106),
            .in2(_gnd_net_),
            .in3(N__12029),
            .lcout(G_463),
            .ltout(G_463_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_9_15_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_9_15_5 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_9_15_5  (
            .in0(N__12041),
            .in1(N__12060),
            .in2(N__12051),
            .in3(N__34722),
            .lcout(\this_vga_ramdac.N_2807_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34601),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_9_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_9_15_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__13107),
            .in2(_gnd_net_),
            .in3(N__12030),
            .lcout(M_this_vga_signals_pixel_clk_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34601),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_15_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_15_7 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_15_7  (
            .in0(N__12012),
            .in1(N__11991),
            .in2(N__11975),
            .in3(N__34725),
            .lcout(\this_vga_ramdac.N_2810_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34601),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_LC_9_25_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_LC_9_25_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_LC_9_25_3  (
            .in0(N__34158),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17427),
            .lcout(M_this_map_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_5_LC_9_25_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_5_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_5_LC_9_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_5_LC_9_25_5  (
            .in0(N__33459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17428),
            .lcout(M_this_map_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_6_LC_9_27_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_6_LC_9_27_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_6_LC_9_27_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_6_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(N__35439),
            .in2(_gnd_net_),
            .in3(N__17397),
            .lcout(M_this_map_ram_write_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_LC_10_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_LC_10_9_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_LC_10_9_0  (
            .in0(N__12795),
            .in1(N__12684),
            .in2(N__16092),
            .in3(N__12702),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_10_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_10_9_1 .LUT_INIT=16'b0111110101000001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_10_9_1  (
            .in0(N__16170),
            .in1(N__12066),
            .in2(N__11934),
            .in3(N__12180),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI8AIVHV_9_LC_10_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI8AIVHV_9_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI8AIVHV_9_LC_10_9_2 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI8AIVHV_9_LC_10_9_2  (
            .in0(N__12867),
            .in1(N__12127),
            .in2(N__12198),
            .in3(N__12744),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_10_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_10_9_3 .LUT_INIT=16'b1011001011101000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_10_9_3  (
            .in0(N__16116),
            .in1(N__12696),
            .in2(N__16175),
            .in3(N__12801),
            .lcout(\this_vga_signals.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__16776),
            .in2(_gnd_net_),
            .in3(N__16542),
            .lcout(\this_vga_signals.vaddress_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_0_LC_10_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_0_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_0_LC_10_9_5 .LUT_INIT=16'b0010011000101010;
    LogicCell40 \this_vga_signals.M_lcounter_q_0_LC_10_9_5  (
            .in0(N__16861),
            .in1(N__17309),
            .in2(N__17022),
            .in3(N__17116),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34545),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_10_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_10_10_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_m2_0_LC_10_10_0  (
            .in0(N__12239),
            .in1(N__13791),
            .in2(N__12297),
            .in3(N__12419),
            .lcout(\this_vga_signals.if_m2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m2_1_LC_10_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m2_1_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m2_1_LC_10_10_1 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \this_vga_signals.un4_haddress_if_m2_1_LC_10_10_1  (
            .in0(N__12418),
            .in1(N__12285),
            .in2(N__13800),
            .in3(N__12236),
            .lcout(\this_vga_signals.if_m2_1 ),
            .ltout(\this_vga_signals.if_m2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_10_2 .LUT_INIT=16'b0101110010100011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_10_2  (
            .in0(N__14966),
            .in1(N__12303),
            .in2(N__12156),
            .in3(N__12332),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI43G6H2_9_LC_10_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI43G6H2_9_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI43G6H2_9_LC_10_10_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI43G6H2_9_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12153),
            .in3(N__12147),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_4_LC_10_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_4_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_4_LC_10_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_4_LC_10_10_4  (
            .in0(N__12690),
            .in1(N__12774),
            .in2(N__12729),
            .in3(N__13452),
            .lcout(\this_vga_signals.g0_i_x4_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam d_m1_2_LC_10_10_5.C_ON=1'b0;
    defparam d_m1_2_LC_10_10_5.SEQ_MODE=4'b0000;
    defparam d_m1_2_LC_10_10_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 d_m1_2_LC_10_10_5 (
            .in0(N__12351),
            .in1(N__12292),
            .in2(_gnd_net_),
            .in3(N__12238),
            .lcout(this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIV3EFO_2_LC_10_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIV3EFO_2_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIV3EFO_2_LC_10_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIV3EFO_2_LC_10_10_6  (
            .in0(N__12237),
            .in1(N__13793),
            .in2(N__12296),
            .in3(N__14960),
            .lcout(\this_vga_signals.d_N_3_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIO08E8_3_LC_10_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIO08E8_3_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIO08E8_3_LC_10_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIO08E8_3_LC_10_10_7  (
            .in0(N__13792),
            .in1(N__14127),
            .in2(_gnd_net_),
            .in3(N__12669),
            .lcout(\this_vga_signals.M_hcounter_q_RNIO08E8Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_10_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_10_11_0 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_10_11_0  (
            .in0(N__14125),
            .in1(N__12821),
            .in2(N__14297),
            .in3(N__12501),
            .lcout(this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_0_1_LC_10_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_0_1_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_0_1_LC_10_11_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_haddress_g1_0_1_LC_10_11_1  (
            .in0(N__14930),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13798),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_2_LC_10_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_2_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_2_LC_10_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g1_2_LC_10_11_2  (
            .in0(N__12234),
            .in1(N__12847),
            .in2(N__12261),
            .in3(N__12503),
            .lcout(),
            .ltout(\this_vga_signals.g1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_2_LC_10_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_2_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_2_LC_10_11_3 .LUT_INIT=16'b0000111110001011;
    LogicCell40 \this_vga_signals.un4_haddress_g0_2_LC_10_11_3  (
            .in0(N__12387),
            .in1(N__12915),
            .in2(N__12258),
            .in3(N__12204),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_o2_0_LC_10_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_o2_0_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_o2_0_LC_10_11_4 .LUT_INIT=16'b0001011101110001;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_o2_0_LC_10_11_4  (
            .in0(N__15024),
            .in1(N__14511),
            .in2(N__12255),
            .in3(N__12252),
            .lcout(\this_vga_signals.mult1_un89_sum_c3_1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_3_LC_10_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_3_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_3_LC_10_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_haddress_g1_3_LC_10_11_5  (
            .in0(N__12502),
            .in1(N__13799),
            .in2(N__12849),
            .in3(N__12233),
            .lcout(\this_vga_signals.N_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_11_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_11_6  (
            .in0(N__14126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12655),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIMID621_5_LC_10_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIMID621_5_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIMID621_5_LC_10_11_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIMID621_5_LC_10_11_7  (
            .in0(N__12656),
            .in1(N__12381),
            .in2(N__12888),
            .in3(N__12402),
            .lcout(\this_vga_signals.g0_i_x4_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_4_LC_10_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_4_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_4_LC_10_12_0 .LUT_INIT=16'b1100100000010011;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_4_LC_10_12_0  (
            .in0(N__14412),
            .in1(N__14220),
            .in2(N__13051),
            .in3(N__12975),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axb1_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_17_LC_10_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_17_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_17_LC_10_12_1 .LUT_INIT=16'b1000011111100001;
    LogicCell40 \this_vga_signals.un4_haddress_g0_17_LC_10_12_1  (
            .in0(N__12651),
            .in1(N__13747),
            .in2(N__12390),
            .in3(N__14057),
            .lcout(\this_vga_signals.g1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_8_LC_10_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_8_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_8_LC_10_12_2 .LUT_INIT=16'b1001101110001001;
    LogicCell40 \this_vga_signals.un4_haddress_g0_8_LC_10_12_2  (
            .in0(N__14056),
            .in1(N__12441),
            .in2(N__13784),
            .in3(N__12650),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_1 ),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_0_LC_10_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_0_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_0_LC_10_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_0_LC_10_12_3  (
            .in0(N__13748),
            .in1(N__12897),
            .in2(N__12375),
            .in3(N__12500),
            .lcout(\this_vga_signals.g1_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_10_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_10_12_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_10_12_4  (
            .in0(N__14055),
            .in1(N__12467),
            .in2(_gnd_net_),
            .in3(N__14216),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_10_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_10_12_5 .LUT_INIT=16'b1111110111110010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_10_12_5  (
            .in0(N__14217),
            .in1(N__13036),
            .in2(N__12366),
            .in3(N__14410),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_12_6 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_12_6  (
            .in0(N__12921),
            .in1(N__12480),
            .in2(N__12363),
            .in3(N__14218),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_10_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_10_12_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_10_12_7  (
            .in0(N__14219),
            .in1(N__13037),
            .in2(N__12507),
            .in3(N__14411),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_10_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_10_13_0 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_10_13_0  (
            .in0(N__13847),
            .in1(N__14401),
            .in2(N__13563),
            .in3(N__13630),
            .lcout(\this_vga_signals.N_6_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_2_9_LC_10_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_2_9_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_2_9_LC_10_13_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_2_9_LC_10_13_1  (
            .in0(N__13629),
            .in1(N__13532),
            .in2(_gnd_net_),
            .in3(N__13846),
            .lcout(\this_vga_signals.N_234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_13_2 .LUT_INIT=16'b1010011100011111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_13_2  (
            .in0(N__13844),
            .in1(N__14400),
            .in2(N__13562),
            .in3(N__13627),
            .lcout(\this_vga_signals.SUM_3 ),
            .ltout(\this_vga_signals.SUM_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_6_1_LC_10_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_6_1_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_6_1_LC_10_13_3 .LUT_INIT=16'b0000010101011111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_6_1_LC_10_13_3  (
            .in0(N__14402),
            .in1(_gnd_net_),
            .in2(N__12456),
            .in3(N__14058),
            .lcout(\this_vga_signals.g0_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_13_4 .LUT_INIT=16'b0011100101100011;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_13_4  (
            .in0(N__13845),
            .in1(N__14399),
            .in2(N__13561),
            .in3(N__13628),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9 ),
            .ltout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIAA7K1_4_LC_10_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIAA7K1_4_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIAA7K1_4_LC_10_13_5 .LUT_INIT=16'b1100000011111100;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIAA7K1_4_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__14059),
            .in2(N__12444),
            .in3(N__14237),
            .lcout(\this_vga_signals.g0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_0_LC_10_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_0_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_0_LC_10_13_6 .LUT_INIT=16'b1100000110000011;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_0_LC_10_13_6  (
            .in0(N__13041),
            .in1(N__12969),
            .in2(N__14266),
            .in3(N__14403),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIC8D41_2_LC_10_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIC8D41_2_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIC8D41_2_LC_10_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIC8D41_2_LC_10_13_7  (
            .in0(N__14404),
            .in1(N__14920),
            .in2(N__13785),
            .in3(N__14238),
            .lcout(\this_vga_signals.g1_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_3_LC_10_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_3_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_3_LC_10_14_0 .LUT_INIT=16'b1100011111000001;
    LogicCell40 \this_vga_signals.un4_haddress_g0_3_LC_10_14_0  (
            .in0(N__13752),
            .in1(N__14086),
            .in2(N__13224),
            .in3(N__12673),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_14_1 .LUT_INIT=16'b1001101100110111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_14_1  (
            .in0(N__13645),
            .in1(N__13542),
            .in2(N__14460),
            .in3(N__13867),
            .lcout(\this_vga_signals.SUM_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_10_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_10_15_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_0_LC_10_15_0  (
            .in0(N__13087),
            .in1(N__12570),
            .in2(_gnd_net_),
            .in3(N__17107),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34588),
            .ce(N__17305),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_10_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_10_15_1 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_1_LC_10_15_1  (
            .in0(N__17108),
            .in1(N__13088),
            .in2(N__13131),
            .in3(N__13151),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34588),
            .ce(N__17305),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_10_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_10_16_1 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_10_16_1  (
            .in0(N__13158),
            .in1(N__14322),
            .in2(N__13885),
            .in3(N__13659),
            .lcout(this_vga_signals_hsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_17_6 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_17_6  (
            .in0(N__13666),
            .in1(N__13579),
            .in2(_gnd_net_),
            .in3(N__13886),
            .lcout(this_vga_signals_hvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_LC_11_8_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_LC_11_8_0 .LUT_INIT=16'b1110011001000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_LC_11_8_0  (
            .in0(N__13248),
            .in1(N__12711),
            .in2(N__15999),
            .in3(N__12513),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI5NOID_3_LC_11_8_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI5NOID_3_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI5NOID_3_LC_11_8_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI5NOID_3_LC_11_8_2  (
            .in0(N__15994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13364),
            .lcout(),
            .ltout(\this_vga_signals.g3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIC44JP1_2_LC_11_8_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIC44JP1_2_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIC44JP1_2_LC_11_8_3 .LUT_INIT=16'b0111110111010111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIC44JP1_2_LC_11_8_3  (
            .in0(N__16089),
            .in1(N__13488),
            .in2(N__12516),
            .in3(N__13449),
            .lcout(\this_vga_signals.g3_0 ),
            .ltout(\this_vga_signals.g3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIGG1CK4_2_LC_11_8_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIGG1CK4_2_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIGG1CK4_2_LC_11_8_4 .LUT_INIT=16'b1010101001011010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIGG1CK4_2_LC_11_8_4  (
            .in0(N__13247),
            .in1(_gnd_net_),
            .in2(N__12756),
            .in3(N__12810),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI90GQ8D_1_LC_11_8_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI90GQ8D_1_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI90GQ8D_1_LC_11_8_5 .LUT_INIT=16'b0110100111110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI90GQ8D_1_LC_11_8_5  (
            .in0(N__14532),
            .in1(N__12753),
            .in2(N__12747),
            .in3(N__13194),
            .lcout(\this_vga_signals.g1_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_11_8_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_11_8_7 .LUT_INIT=16'b1001000110111001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_LC_11_8_7  (
            .in0(N__13203),
            .in1(N__13188),
            .in2(N__12738),
            .in3(N__15114),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x0_LC_11_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x0_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x0_LC_11_9_0 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x0_LC_11_9_0  (
            .in0(N__14619),
            .in1(N__14579),
            .in2(N__13377),
            .in3(N__13926),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_ns_LC_11_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_ns_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_ns_LC_11_9_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_ns_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__13437),
            .in2(N__12714),
            .in3(N__12762),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_ns ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_11_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_11_9_2 .LUT_INIT=16'b1110010111011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_LC_11_9_2  (
            .in0(N__13441),
            .in1(N__15982),
            .in2(N__12705),
            .in3(N__13266),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_11_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_11_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_11_9_3  (
            .in0(N__14580),
            .in1(N__16779),
            .in2(_gnd_net_),
            .in3(N__13178),
            .lcout(\this_vga_signals.g0_i_x4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_1_LC_11_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_1_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_1_LC_11_9_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_1_LC_11_9_4  (
            .in0(N__16541),
            .in1(_gnd_net_),
            .in2(N__13378),
            .in3(N__16084),
            .lcout(\this_vga_signals.g0_i_x4_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_11_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_11_9_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_11_9_5  (
            .in0(N__13375),
            .in1(N__15998),
            .in2(N__12789),
            .in3(N__13442),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_9_6 .LUT_INIT=16'b0001001000100001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_9_6  (
            .in0(N__13359),
            .in1(N__15981),
            .in2(N__13451),
            .in3(N__12785),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_2 ),
            .ltout(\this_vga_signals.mult1_un68_sum_ac0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_11_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_11_9_7 .LUT_INIT=16'b0000110100000111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_LC_11_9_7  (
            .in0(N__16085),
            .in1(N__13179),
            .in2(N__12804),
            .in3(N__12768),
            .lcout(\this_vga_signals.g1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_11_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_11_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_11_10_1  (
            .in0(N__13367),
            .in1(N__15990),
            .in2(N__16778),
            .in3(N__13436),
            .lcout(\this_vga_signals.g0_2_0_a2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_11_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_11_10_2 .LUT_INIT=16'b0011001110011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_11_10_2  (
            .in0(N__14618),
            .in1(N__14571),
            .in2(_gnd_net_),
            .in3(N__13921),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_11_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_11_10_3 .LUT_INIT=16'b0000001100111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__15989),
            .in2(N__12777),
            .in3(N__16762),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_11_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_11_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_2_LC_11_10_4  (
            .in0(N__15987),
            .in1(N__14572),
            .in2(N__13450),
            .in3(N__13365),
            .lcout(\this_vga_signals.g0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_0_a3_LC_11_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_a3_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_a3_LC_11_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_0_a3_LC_11_10_5  (
            .in0(N__13366),
            .in1(N__15988),
            .in2(N__16777),
            .in3(N__13435),
            .lcout(\this_vga_signals.N_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x1_LC_11_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x1_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x1_LC_11_10_6 .LUT_INIT=16'b1100001101101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x1_LC_11_10_6  (
            .in0(N__14617),
            .in1(N__14570),
            .in2(N__13376),
            .in3(N__13920),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_11_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_11_10_7 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_11_10_7  (
            .in0(N__16620),
            .in1(N__16761),
            .in2(_gnd_net_),
            .in3(N__16515),
            .lcout(\this_vga_signals.vaddress_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_11_LC_11_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_11_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_11_LC_11_11_0 .LUT_INIT=16'b1101110110111011;
    LogicCell40 \this_vga_signals.un4_haddress_g0_11_LC_11_11_0  (
            .in0(N__13065),
            .in1(N__14094),
            .in2(_gnd_net_),
            .in3(N__14262),
            .lcout(\this_vga_signals.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIF18M2_5_LC_11_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIF18M2_5_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIF18M2_5_LC_11_11_3 .LUT_INIT=16'b0110010011011001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIF18M2_5_LC_11_11_3  (
            .in0(N__13053),
            .in1(N__12981),
            .in2(N__14288),
            .in3(N__14459),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_x4_2_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI42KN6_5_LC_11_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI42KN6_5_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI42KN6_5_LC_11_11_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI42KN6_5_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12891),
            .in3(N__12848),
            .lcout(\this_vga_signals.g0_i_x4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_0_a2_LC_11_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_0_a2_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_0_a2_LC_11_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_0_a2_LC_11_11_5  (
            .in0(N__13380),
            .in1(N__13902),
            .in2(_gnd_net_),
            .in3(N__13445),
            .lcout(),
            .ltout(\this_vga_signals.N_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_11_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_11_11_6 .LUT_INIT=16'b1101010000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_LC_11_11_6  (
            .in0(N__16078),
            .in1(N__15992),
            .in2(N__12879),
            .in3(N__12876),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_11_7 .LUT_INIT=16'b1011001000101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_11_7  (
            .in0(N__16079),
            .in1(N__16174),
            .in2(N__12870),
            .in3(N__13302),
            .lcout(\this_vga_signals.mult1_un75_sum_c2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIL0C14_6_LC_11_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIL0C14_6_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIL0C14_6_LC_11_12_0 .LUT_INIT=16'b0000111001110000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIL0C14_6_LC_11_12_0  (
            .in0(N__14408),
            .in1(N__13032),
            .in2(N__12858),
            .in3(N__12968),
            .lcout(\this_vga_signals.N_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_a0_0_LC_11_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_a0_0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_a0_0_LC_11_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_a0_0_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__14210),
            .in2(_gnd_net_),
            .in3(N__14406),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_a0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_12_3 .LUT_INIT=16'b1011101010100010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_12_3  (
            .in0(N__12967),
            .in1(N__14215),
            .in2(N__13050),
            .in3(N__14409),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_13_LC_11_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_13_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_13_LC_11_12_4 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \this_vga_signals.un4_haddress_g0_13_LC_11_12_4  (
            .in0(N__14407),
            .in1(N__13031),
            .in2(N__14254),
            .in3(N__12966),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_11_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_11_12_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_11_12_5  (
            .in0(N__14054),
            .in1(N__14211),
            .in2(_gnd_net_),
            .in3(N__14405),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_11_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_11_12_6 .LUT_INIT=16'b1111111101110000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_11_12_6  (
            .in0(N__13059),
            .in1(N__13030),
            .in2(N__12984),
            .in3(N__12965),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_19_LC_11_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_19_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_19_LC_11_12_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un4_haddress_g0_19_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__15009),
            .in2(_gnd_net_),
            .in3(N__14919),
            .lcout(\this_vga_signals.if_N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_13_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__14505),
            .in2(N__15023),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_11_13_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_11_13_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_11_13_1  (
            .in0(N__17268),
            .in1(N__14929),
            .in2(_gnd_net_),
            .in3(N__12909),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__34566),
            .ce(),
            .sr(N__14849));
    defparam \this_vga_signals.M_hcounter_q_3_LC_11_13_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_11_13_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_11_13_2  (
            .in0(N__17306),
            .in1(N__13783),
            .in2(_gnd_net_),
            .in3(N__12906),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__34566),
            .ce(),
            .sr(N__14849));
    defparam \this_vga_signals.M_hcounter_q_4_LC_11_13_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_11_13_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_11_13_3  (
            .in0(N__17269),
            .in1(N__14087),
            .in2(_gnd_net_),
            .in3(N__12903),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__34566),
            .ce(),
            .sr(N__14849));
    defparam \this_vga_signals.M_hcounter_q_5_LC_11_13_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_11_13_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_11_13_4  (
            .in0(N__17307),
            .in1(N__14248),
            .in2(_gnd_net_),
            .in3(N__12900),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__34566),
            .ce(),
            .sr(N__14849));
    defparam \this_vga_signals.M_hcounter_q_6_LC_11_13_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_11_13_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_11_13_5  (
            .in0(N__17270),
            .in1(N__14438),
            .in2(_gnd_net_),
            .in3(N__13170),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__34566),
            .ce(),
            .sr(N__14849));
    defparam \this_vga_signals.M_hcounter_q_7_LC_11_13_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_11_13_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_11_13_6  (
            .in0(N__17308),
            .in1(N__13868),
            .in2(_gnd_net_),
            .in3(N__13167),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__34566),
            .ce(),
            .sr(N__14849));
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_13_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_13_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_11_13_7  (
            .in0(N__17271),
            .in1(N__13560),
            .in2(_gnd_net_),
            .in3(N__13164),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__34566),
            .ce(),
            .sr(N__14849));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_11_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_11_14_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__13655),
            .in2(_gnd_net_),
            .in3(N__13161),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34574),
            .ce(N__14520),
            .sr(N__14853));
    defparam \this_vga_signals.M_hcounter_q_RNISKQ82_7_LC_11_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNISKQ82_7_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNISKQ82_7_LC_11_15_1 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNISKQ82_7_LC_11_15_1  (
            .in0(N__13570),
            .in1(N__13992),
            .in2(N__13884),
            .in3(N__14449),
            .lcout(\this_vga_signals.un4_hsynclt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_11_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_11_15_2 .LUT_INIT=16'b1101110110111011;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_11_15_2  (
            .in0(N__13643),
            .in1(N__13569),
            .in2(_gnd_net_),
            .in3(N__13869),
            .lcout(\this_vga_signals.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_11_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_11_15_3 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_11_15_3  (
            .in0(N__13086),
            .in1(N__13152),
            .in2(N__13130),
            .in3(N__17056),
            .lcout(),
            .ltout(\this_vga_signals.M_pcounter_q_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_11_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_11_15_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__13126),
            .in2(N__13110),
            .in3(N__17301),
            .lcout(N_3_0),
            .ltout(N_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_LC_11_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_11_15_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13095),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_pcounter_q_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34580),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_15_6 .LUT_INIT=16'b1001101100110111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_15_6  (
            .in0(N__13644),
            .in1(N__13568),
            .in2(N__14463),
            .in3(N__13870),
            .lcout(),
            .ltout(\this_vga_signals.SUM_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_LC_11_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_LC_11_15_7 .LUT_INIT=16'b0010011010010001;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_LC_11_15_7  (
            .in0(N__14261),
            .in1(N__13233),
            .in2(N__13227),
            .in3(N__14448),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_4_LC_11_27_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_4_LC_11_27_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_4_LC_11_27_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_4_LC_11_27_5  (
            .in0(_gnd_net_),
            .in1(N__33574),
            .in2(_gnd_net_),
            .in3(N__17432),
            .lcout(M_this_map_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_12_8_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_12_8_1 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_LC_12_8_1  (
            .in0(N__16346),
            .in1(N__15252),
            .in2(N__13965),
            .in3(N__14766),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_a2_0_LC_12_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_a2_0_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_a2_0_LC_12_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_a2_0_LC_12_9_0  (
            .in0(N__15980),
            .in1(N__13444),
            .in2(_gnd_net_),
            .in3(N__13374),
            .lcout(),
            .ltout(\this_vga_signals.N_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQJ81Q1_1_LC_12_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQJ81Q1_1_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQJ81Q1_1_LC_12_9_1 .LUT_INIT=16'b0110000000000110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQJ81Q1_1_LC_12_9_1  (
            .in0(N__16071),
            .in1(N__16155),
            .in2(N__13197),
            .in3(N__13487),
            .lcout(\this_vga_signals.g1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_12_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_12_9_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_12_9_3  (
            .in0(N__16760),
            .in1(N__16628),
            .in2(_gnd_net_),
            .in3(N__16536),
            .lcout(\this_vga_signals.vaddress_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_0_m2_LC_12_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_m2_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_m2_LC_12_9_4 .LUT_INIT=16'b0001100010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_0_m2_LC_12_9_4  (
            .in0(N__16537),
            .in1(N__15106),
            .in2(N__15060),
            .in3(N__14744),
            .lcout(),
            .ltout(\this_vga_signals.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_12_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_12_9_5 .LUT_INIT=16'b0101010101110101;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_LC_12_9_5  (
            .in0(N__14622),
            .in1(N__16780),
            .in2(N__13182),
            .in3(N__14703),
            .lcout(\this_vga_signals.g1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_661_LC_12_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_661_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_661_LC_12_9_6 .LUT_INIT=16'b0001111001111000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_661_LC_12_9_6  (
            .in0(N__14664),
            .in1(N__16759),
            .in2(N__14708),
            .in3(N__13470),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_661 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axb1_661_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__15979),
            .in2(N__13269),
            .in3(N__16781),
            .lcout(\this_vga_signals.g0_2_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_10_0 .LUT_INIT=16'b0001010000010100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_10_0  (
            .in0(N__15159),
            .in1(N__15232),
            .in2(N__15375),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\this_vga_signals.if_N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_12_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_12_10_1 .LUT_INIT=16'b0000110100001110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_LC_12_10_1  (
            .in0(N__15048),
            .in1(N__14659),
            .in2(N__13260),
            .in3(N__15100),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_12_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_12_10_2 .LUT_INIT=16'b0001100010000001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_12_10_2  (
            .in0(N__15983),
            .in1(N__15233),
            .in2(N__13257),
            .in3(N__14568),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_12_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_12_10_3 .LUT_INIT=16'b1010011010101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_12_10_3  (
            .in0(N__16769),
            .in1(N__14660),
            .in2(N__13254),
            .in3(N__13473),
            .lcout(\this_vga_signals.mult1_un61_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a2_0_LC_12_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a2_0_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a2_0_LC_12_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_0_a2_0_LC_12_10_4  (
            .in0(N__15984),
            .in1(N__16770),
            .in2(N__13251),
            .in3(N__13363),
            .lcout(\this_vga_signals.N_4_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_10_5 .LUT_INIT=16'b1000010111100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_10_5  (
            .in0(N__15047),
            .in1(N__14658),
            .in2(N__14745),
            .in3(N__15099),
            .lcout(\this_vga_signals.mult1_un47_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_12_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_12_10_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_LC_12_10_6  (
            .in0(N__16517),
            .in1(N__16768),
            .in2(N__13236),
            .in3(N__14707),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_3_d_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_a2_0_1_LC_12_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_a2_0_1_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_a2_0_1_LC_12_10_7 .LUT_INIT=16'b0101101001010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_a2_0_1_LC_12_10_7  (
            .in0(N__14569),
            .in1(_gnd_net_),
            .in2(N__13491),
            .in3(N__14610),
            .lcout(\this_vga_signals.g0_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIEQV87_2_LC_12_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIEQV87_2_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIEQV87_2_LC_12_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIEQV87_2_LC_12_11_0  (
            .in0(N__13472),
            .in1(N__15986),
            .in2(N__16090),
            .in3(N__16538),
            .lcout(\this_vga_signals.g2_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_12_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_12_11_1 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_12_11_1  (
            .in0(N__15234),
            .in1(N__14663),
            .in2(N__14709),
            .in3(N__13471),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_3_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_12_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_12_11_2 .LUT_INIT=16'b1111111110111101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_12_11_2  (
            .in0(N__14662),
            .in1(N__15050),
            .in2(N__15110),
            .in3(N__14746),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_12_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_12_11_3 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_LC_12_11_3  (
            .in0(N__16771),
            .in1(N__15991),
            .in2(_gnd_net_),
            .in3(N__13901),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_2_LC_12_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_2_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_2_LC_12_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_2_LC_12_11_4  (
            .in0(N__13284),
            .in1(N__13443),
            .in2(N__13383),
            .in3(N__13379),
            .lcout(\this_vga_signals.g0_i_x4_0_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_0_LC_12_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_0_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_0_LC_12_11_6 .LUT_INIT=16'b0110011011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_0_LC_12_11_6  (
            .in0(N__15120),
            .in1(N__16539),
            .in2(N__13296),
            .in3(N__14747),
            .lcout(\this_vga_signals.g0_i_x4_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_11_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_11_7  (
            .in0(N__16540),
            .in1(N__16278),
            .in2(N__16782),
            .in3(N__16425),
            .lcout(\this_vga_signals.vsync_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_12_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_12_0  (
            .in0(N__16083),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16347),
            .lcout(),
            .ltout(\this_vga_signals.vsync_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_12_1 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_12_1  (
            .in0(N__13932),
            .in1(N__13278),
            .in2(N__13272),
            .in3(N__16629),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_12_2 .LUT_INIT=16'b0000000101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_12_2  (
            .in0(N__16775),
            .in1(N__16176),
            .in2(N__16091),
            .in3(N__15993),
            .lcout(\this_vga_signals.un2_vsynclt8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_1_i_o3_LC_12_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_1_i_o3_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_1_i_o3_LC_12_12_7 .LUT_INIT=16'b0000001110101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_1_i_o3_LC_12_12_7  (
            .in0(N__14621),
            .in1(N__14748),
            .in2(N__15069),
            .in3(N__13922),
            .lcout(\this_vga_signals.mult1_un54_sum_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_12_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_12_13_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_12_13_0  (
            .in0(N__15016),
            .in1(N__14507),
            .in2(_gnd_net_),
            .in3(N__17300),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34560),
            .ce(),
            .sr(N__14848));
    defparam \this_vga_signals.M_hcounter_q_0_LC_12_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_12_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__14506),
            .in2(_gnd_net_),
            .in3(N__17299),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34560),
            .ce(),
            .sr(N__14848));
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_14_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_14_0  (
            .in0(N__14209),
            .in1(N__14431),
            .in2(_gnd_net_),
            .in3(N__13843),
            .lcout(\this_vga_signals.M_hcounter_d7lto7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__13724),
            .in2(_gnd_net_),
            .in3(N__14905),
            .lcout(\this_vga_signals.un2_hsynclto3_0 ),
            .ltout(\this_vga_signals.un2_hsynclto3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_14_2 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_14_2  (
            .in0(N__15017),
            .in1(N__14500),
            .in2(N__13677),
            .in3(N__14053),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_d7lt7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_14_3 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_14_3  (
            .in0(N__13674),
            .in1(N__13631),
            .in2(N__13584),
            .in3(N__13559),
            .lcout(\this_vga_signals.M_hcounter_d7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_14_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__14838),
            .in2(_gnd_net_),
            .in3(N__17288),
            .lcout(\this_vga_signals.N_852_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_12_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_12_14_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_12_14_7  (
            .in0(N__14501),
            .in1(N__14309),
            .in2(_gnd_net_),
            .in3(N__15018),
            .lcout(\this_vga_signals.un2_hsynclt6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_4_LC_12_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_4_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_4_LC_12_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIEVMV1_4_LC_12_15_3  (
            .in0(N__14475),
            .in1(N__14137),
            .in2(N__14295),
            .in3(N__14461),
            .lcout(\this_vga_signals.un2_hsynclt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_15_6 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_15_6  (
            .in0(N__14310),
            .in1(N__14278),
            .in2(N__14139),
            .in3(N__15019),
            .lcout(\this_vga_signals.un4_hsynclto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_1_LC_12_25_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_1_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_1_LC_12_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_1_LC_12_25_6  (
            .in0(_gnd_net_),
            .in1(N__33979),
            .in2(_gnd_net_),
            .in3(N__17406),
            .lcout(M_this_map_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIT6RN_8_LC_13_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIT6RN_8_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIT6RN_8_LC_13_9_0 .LUT_INIT=16'b1111001111010011;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIT6RN_8_LC_13_9_0  (
            .in0(N__15142),
            .in1(N__16423),
            .in2(N__15273),
            .in3(N__13974),
            .lcout(\this_vga_signals.SUM_2_i_1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_13_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_13_9_1 .LUT_INIT=16'b0000001100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__14783),
            .in2(N__15371),
            .in3(N__14806),
            .lcout(\this_vga_signals.SUM_2_i_1_1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_13_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_13_9_2 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_13_9_2  (
            .in0(N__14807),
            .in1(N__15364),
            .in2(_gnd_net_),
            .in3(N__14817),
            .lcout(),
            .ltout(\this_vga_signals.N_1_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNITUMI_8_LC_13_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNITUMI_8_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNITUMI_8_LC_13_9_3 .LUT_INIT=16'b1101111111001111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNITUMI_8_LC_13_9_3  (
            .in0(N__16424),
            .in1(N__15182),
            .in2(N__13968),
            .in3(N__15272),
            .lcout(\this_vga_signals.SUM_2_i_1_2_3 ),
            .ltout(\this_vga_signals.SUM_2_i_1_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_13_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_13_9_4 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_13_9_4  (
            .in0(N__16319),
            .in1(N__15245),
            .in2(N__14769),
            .in3(N__14765),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_N_2L1_LC_13_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_N_2L1_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_N_2L1_LC_13_9_7 .LUT_INIT=16'b0011111111111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_N_2L1_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__14782),
            .in2(N__15370),
            .in3(N__14805),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x0_LC_13_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x0_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x0_LC_13_10_0 .LUT_INIT=16'b1010001010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x0_LC_13_10_0  (
            .in0(N__16274),
            .in1(N__15141),
            .in2(N__14682),
            .in3(N__16412),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_ns_LC_13_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_ns_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_ns_LC_13_10_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_ns_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__14790),
            .in2(N__14754),
            .in3(N__14670),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_10_2 .LUT_INIT=16'b0001100011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_10_2  (
            .in0(N__15049),
            .in1(N__14661),
            .in2(N__14751),
            .in3(N__14732),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x1_LC_13_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x1_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x1_LC_13_10_3 .LUT_INIT=16'b1001001100010011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x1_LC_13_10_3  (
            .in0(N__16411),
            .in1(N__16273),
            .in2(N__15146),
            .in3(N__14678),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_13_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_13_10_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_13_10_4  (
            .in0(N__16486),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15216),
            .lcout(\this_vga_signals.vaddress_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.g2_0_a2_5_1_LC_13_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.g2_0_a2_5_1_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.g2_0_a2_5_1_LC_13_10_5 .LUT_INIT=16'b0100010010111011;
    LogicCell40 \this_vga_signals.g2_0_a2_5_1_LC_13_10_5  (
            .in0(N__14631),
            .in1(N__14620),
            .in2(_gnd_net_),
            .in3(N__14578),
            .lcout(),
            .ltout(\this_vga_signals.g2_0_a2_5Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIUR0A01_3_LC_13_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIUR0A01_3_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIUR0A01_3_LC_13_10_6 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIUR0A01_3_LC_13_10_6  (
            .in0(N__15985),
            .in1(N__16746),
            .in2(N__14541),
            .in3(N__14538),
            .lcout(\this_vga_signals.g2_0_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_LC_13_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_LC_13_11_0 .LUT_INIT=16'b0101001101001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_LC_13_11_0  (
            .in0(N__15105),
            .in1(N__16508),
            .in2(N__16619),
            .in3(N__16709),
            .lcout(\this_vga_signals.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_13_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_13_11_3 .LUT_INIT=16'b0111111010011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_3_LC_13_11_3  (
            .in0(N__16708),
            .in1(N__16511),
            .in2(N__16614),
            .in3(N__15104),
            .lcout(\this_vga_signals.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_13_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_13_11_5 .LUT_INIT=16'b1010010100001111;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_13_11_5  (
            .in0(N__15223),
            .in1(_gnd_net_),
            .in2(N__15186),
            .in3(N__16510),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m2_LC_13_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m2_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m2_LC_13_12_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_m2_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__15008),
            .in2(_gnd_net_),
            .in3(N__14959),
            .lcout(\this_vga_signals.if_m2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_13_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_13_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__17253),
            .in2(_gnd_net_),
            .in3(N__17067),
            .lcout(\this_vga_signals.N_1098_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_8_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15600),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34515),
            .ce(N__15504),
            .sr(N__15472));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_8_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15549),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34515),
            .ce(N__15504),
            .sr(N__15472));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_N_2L1_LC_14_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_N_2L1_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_N_2L1_LC_14_9_0 .LUT_INIT=16'b0001010101111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_N_2L1_LC_14_9_0  (
            .in0(N__14784),
            .in1(N__15366),
            .in2(N__14811),
            .in3(N__15263),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1_0_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15566),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34521),
            .ce(N__15513),
            .sr(N__15474));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_14_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_14_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15525),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34521),
            .ce(N__15513),
            .sr(N__15474));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIQE4H_LC_14_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIQE4H_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIQE4H_LC_14_9_4 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIQE4H_LC_14_9_4  (
            .in0(N__15177),
            .in1(N__15212),
            .in2(_gnd_net_),
            .in3(N__15365),
            .lcout(\this_vga_signals.vaddress_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_14_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_14_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15565),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34521),
            .ce(N__15513),
            .sr(N__15474));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_14_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_14_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15598),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34521),
            .ce(N__15513),
            .sr(N__15474));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_14_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_14_9_7 .LUT_INIT=16'b0110110110110111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_14_9_7  (
            .in0(N__16407),
            .in1(N__16266),
            .in2(N__15147),
            .in3(N__15178),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15599),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__15509),
            .sr(N__15476));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_14_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_14_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15578),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__15509),
            .sr(N__15476));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_10_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15547),
            .lcout(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__15509),
            .sr(N__15476));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_14_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_14_10_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_14_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_14_10_3  (
            .in0(N__15548),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__15509),
            .sr(N__15476));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_14_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_14_10_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_14_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15567),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__15509),
            .sr(N__15476));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_10_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_10_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_10_6  (
            .in0(N__15579),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__15509),
            .sr(N__15476));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_14_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_14_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__16320),
            .in2(_gnd_net_),
            .in3(N__16269),
            .lcout(),
            .ltout(\this_vga_signals.un6_vvisibilitylto8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_14_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_14_11_2 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_14_11_2  (
            .in0(N__16506),
            .in1(N__16603),
            .in2(N__15336),
            .in3(N__16710),
            .lcout(),
            .ltout(\this_vga_signals.un6_vvisibilitylt9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNINQIT3_5_LC_14_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNINQIT3_5_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNINQIT3_5_LC_14_11_3 .LUT_INIT=16'b0000101100000011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNINQIT3_5_LC_14_11_3  (
            .in0(N__16711),
            .in1(N__15282),
            .in2(N__15333),
            .in3(N__16507),
            .lcout(this_vga_signals_vvisibility_1),
            .ltout(this_vga_signals_vvisibility_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM8094_9_LC_14_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM8094_9_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM8094_9_LC_14_11_4 .LUT_INIT=16'b0011000000110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIM8094_9_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__16409),
            .in2(N__15330),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.vvisibility ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_14_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_14_11_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_14_11_6  (
            .in0(N__16268),
            .in1(N__16408),
            .in2(N__16337),
            .in3(N__16602),
            .lcout(\this_vga_signals.vaddress_ac0_9_0_a0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI01PG1_0_1_LC_14_12_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI01PG1_0_1_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI01PG1_0_1_LC_14_12_6 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_ppu.M_state_q_RNI01PG1_0_1_LC_14_12_6  (
            .in0(N__20977),
            .in1(N__18442),
            .in2(_gnd_net_),
            .in3(N__35075),
            .lcout(\this_ppu.N_1195_0_1 ),
            .ltout(\this_ppu.N_1195_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_0_LC_14_12_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_0_LC_14_12_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_0_LC_14_12_7 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \this_ppu.M_count_q_0_LC_14_12_7  (
            .in0(N__15645),
            .in1(N__20978),
            .in2(N__15276),
            .in3(N__21527),
            .lcout(\this_ppu.M_count_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34537),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_13_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__15644),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_13_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__15804),
            .in2(N__20081),
            .in3(N__15405),
            .lcout(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_13_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__20030),
            .in2(N__15825),
            .in3(N__15402),
            .lcout(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_13_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__20034),
            .in2(N__15722),
            .in3(N__15399),
            .lcout(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_13_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__15860),
            .in2(N__20083),
            .in3(N__15396),
            .lcout(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_13_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__15879),
            .in2(N__20082),
            .in3(N__15393),
            .lcout(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_13_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__15842),
            .in2(N__20084),
            .in3(N__15390),
            .lcout(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_7_LC_14_13_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_14_13_7 .LUT_INIT=16'b1111000000011110;
    LogicCell40 \this_ppu.M_count_q_RNO_0_7_LC_14_13_7  (
            .in0(N__21012),
            .in1(N__21533),
            .in2(N__15693),
            .in3(N__15387),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_14_14_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_14_14_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_14_14_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__34816),
            .in2(_gnd_net_),
            .in3(N__17475),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34553),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_14_16_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_14_16_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__34829),
            .in2(_gnd_net_),
            .in3(N__15384),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34567),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_14_18_3 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_14_18_3 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_14_18_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_14_18_3  (
            .in0(N__15450),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34581),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_14_18_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_14_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15420),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34581),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_14_18_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_14_18_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_14_18_6  (
            .in0(N__34837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15435),
            .lcout(\this_reset_cond.M_stage_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34581),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_14_18_7 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_14_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15426),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34581),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_15_8_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_15_8_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__17282),
            .in2(_gnd_net_),
            .in3(N__15480),
            .lcout(\this_vga_signals.N_852_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_15_9_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_15_9_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_15_9_0  (
            .in0(N__17284),
            .in1(N__16115),
            .in2(N__17117),
            .in3(N__17115),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__34516),
            .ce(),
            .sr(N__15473));
    defparam \this_vga_signals.M_vcounter_q_1_LC_15_9_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_15_9_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_15_9_1  (
            .in0(N__17286),
            .in1(N__16151),
            .in2(_gnd_net_),
            .in3(N__15414),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__34516),
            .ce(),
            .sr(N__15473));
    defparam \this_vga_signals.M_vcounter_q_2_LC_15_9_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_15_9_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_15_9_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_15_9_2  (
            .in0(N__17285),
            .in1(N__16047),
            .in2(_gnd_net_),
            .in3(N__15411),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__34516),
            .ce(),
            .sr(N__15473));
    defparam \this_vga_signals.M_vcounter_q_3_LC_15_9_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_15_9_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_15_9_3  (
            .in0(N__17287),
            .in1(N__15941),
            .in2(_gnd_net_),
            .in3(N__15408),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__34516),
            .ce(),
            .sr(N__15473));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_9_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__16715),
            .in2(_gnd_net_),
            .in3(N__15582),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_15_9_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_15_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__16509),
            .in2(_gnd_net_),
            .in3(N__15570),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_9_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__16610),
            .in2(_gnd_net_),
            .in3(N__15552),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_15_9_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_15_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__16336),
            .in2(_gnd_net_),
            .in3(N__15534),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_15_10_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_15_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__16272),
            .in2(_gnd_net_),
            .in3(N__15531),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_15_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_15_10_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_15_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__16410),
            .in2(_gnd_net_),
            .in3(N__15528),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34522),
            .ce(N__15505),
            .sr(N__15475));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_15_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_15_10_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_15_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15524),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34522),
            .ce(N__15505),
            .sr(N__15475));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_15_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_15_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_15_11_0  (
            .in0(N__16487),
            .in1(N__16335),
            .in2(N__16615),
            .in3(N__16267),
            .lcout(\this_vga_signals.M_vcounter_d7lto8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI4GQN4_0_LC_15_11_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI4GQN4_0_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI4GQN4_0_LC_15_11_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_ppu.M_state_q_RNI4GQN4_0_LC_15_11_3  (
            .in0(N__21575),
            .in1(N__21661),
            .in2(_gnd_net_),
            .in3(N__21616),
            .lcout(\this_ppu.N_132_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI4L615_0_LC_15_12_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI4L615_0_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI4L615_0_LC_15_12_0 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \this_ppu.M_state_q_RNI4L615_0_LC_15_12_0  (
            .in0(N__21628),
            .in1(N__21591),
            .in2(N__20995),
            .in3(N__21663),
            .lcout(\this_ppu.un16_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI4HJ86_0_LC_15_12_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI4HJ86_0_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI4HJ86_0_LC_15_12_2 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \this_ppu.M_state_q_RNI4HJ86_0_LC_15_12_2  (
            .in0(N__21627),
            .in1(N__21662),
            .in2(N__21602),
            .in3(N__15656),
            .lcout(\this_ppu.N_1195_0 ),
            .ltout(\this_ppu.N_1195_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_2_LC_15_12_3 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_2_LC_15_12_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_2_LC_15_12_3 .LUT_INIT=16'b1010000010010000;
    LogicCell40 \this_ppu.M_count_q_2_LC_15_12_3  (
            .in0(N__15824),
            .in1(N__15769),
            .in2(N__15666),
            .in3(N__15663),
            .lcout(\this_ppu.M_count_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34531),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_0_LC_15_12_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_0_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_0_LC_15_12_5 .LUT_INIT=16'b1011001111110011;
    LogicCell40 \this_ppu.M_state_q_0_LC_15_12_5  (
            .in0(N__21592),
            .in1(N__15657),
            .in2(N__21673),
            .in3(N__21629),
            .lcout(\this_ppu.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34531),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIL508_7_LC_15_13_0 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIL508_7_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIL508_7_LC_15_13_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_count_q_RNIL508_7_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__15686),
            .in2(_gnd_net_),
            .in3(N__15643),
            .lcout(\this_ppu.M_count_d_1_sqmuxa_1_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_1_LC_15_13_1 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_1_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_1_LC_15_13_1 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_1_LC_15_13_1  (
            .in0(N__15803),
            .in1(N__15770),
            .in2(N__15627),
            .in3(N__15737),
            .lcout(\this_ppu.M_count_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34538),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_5_LC_15_13_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_5_LC_15_13_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_5_LC_15_13_2 .LUT_INIT=16'b1010100000000010;
    LogicCell40 \this_ppu.M_count_q_5_LC_15_13_2  (
            .in0(N__15740),
            .in1(N__15618),
            .in2(N__15779),
            .in3(N__15878),
            .lcout(\this_ppu.M_count_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34538),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_4_LC_15_13_3 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_4_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_4_LC_15_13_3 .LUT_INIT=16'b1110000100000000;
    LogicCell40 \this_ppu.M_count_q_4_LC_15_13_3  (
            .in0(N__15612),
            .in1(N__15772),
            .in2(N__15864),
            .in3(N__15739),
            .lcout(\this_ppu.M_count_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34538),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_6_LC_15_13_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_6_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_6_LC_15_13_4 .LUT_INIT=16'b1010100000000010;
    LogicCell40 \this_ppu.M_count_q_6_LC_15_13_4  (
            .in0(N__15741),
            .in1(N__15606),
            .in2(N__15780),
            .in3(N__15841),
            .lcout(\this_ppu.M_count_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34538),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIDE0G_2_LC_15_13_5 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIDE0G_2_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIDE0G_2_LC_15_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_count_q_RNIDE0G_2_LC_15_13_5  (
            .in0(N__15877),
            .in1(N__15859),
            .in2(N__15843),
            .in3(N__15820),
            .lcout(),
            .ltout(\this_ppu.M_count_d_1_sqmuxa_1_i_a2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIKM001_1_LC_15_13_6 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIKM001_1_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIKM001_1_LC_15_13_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_ppu.M_count_q_RNIKM001_1_LC_15_13_6  (
            .in0(N__15715),
            .in1(N__15802),
            .in2(N__15789),
            .in3(N__15786),
            .lcout(\this_ppu.M_count_d_0_sqmuxa_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_3_LC_15_13_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_3_LC_15_13_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_3_LC_15_13_7 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_3_LC_15_13_7  (
            .in0(N__15723),
            .in1(N__15771),
            .in2(N__15750),
            .in3(N__15738),
            .lcout(\this_ppu.M_count_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34538),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_0_LC_15_14_0 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_15_14_0 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_15_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16821),
            .lcout(this_pixel_clk_M_counter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34546),
            .ce(),
            .sr(N__34994));
    defparam \this_ppu.M_count_q_7_LC_15_14_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_7_LC_15_14_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_7_LC_15_14_7 .LUT_INIT=16'b0101111101001100;
    LogicCell40 \this_ppu.M_count_q_7_LC_15_14_7  (
            .in0(N__18448),
            .in1(N__15699),
            .in2(N__21020),
            .in3(N__21534),
            .lcout(\this_ppu.M_count_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34546),
            .ce(),
            .sr(N__34994));
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_2_1_LC_15_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_2_1_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_2_1_LC_15_15_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_2_1_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__17859),
            .in2(_gnd_net_),
            .in3(N__35088),
            .lcout(\this_vga_signals.N_85 ),
            .ltout(\this_vga_signals.N_85_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_15_15_1.C_ON=1'b0;
    defparam M_this_state_q_5_LC_15_15_1.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_15_15_1.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_5_LC_15_15_1 (
            .in0(N__15672),
            .in1(N__21476),
            .in2(N__15675),
            .in3(N__22981),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34554),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_i_1_5_LC_15_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_i_1_5_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_i_1_5_LC_15_15_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_i_1_5_LC_15_15_4  (
            .in0(N__17837),
            .in1(N__17765),
            .in2(_gnd_net_),
            .in3(N__17682),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_444_i_i_o2_LC_15_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.N_444_i_i_o2_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_444_i_i_o2_LC_15_15_6 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \this_vga_signals.N_444_i_i_o2_LC_15_15_6  (
            .in0(N__20898),
            .in1(_gnd_net_),
            .in2(N__21765),
            .in3(N__23144),
            .lcout(\this_vga_signals.N_124_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_1_LC_15_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_1_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_1_LC_15_16_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_1_LC_15_16_0  (
            .in0(N__17761),
            .in1(N__16216),
            .in2(N__17838),
            .in3(N__17680),
            .lcout(this_vga_signals_M_this_state_q_srsts_0_1_i_a2_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_2_LC_15_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_2_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_2_LC_15_16_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_2_LC_15_16_4  (
            .in0(N__17836),
            .in1(N__16217),
            .in2(N__17766),
            .in3(N__17681),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_15_16_5.C_ON=1'b0;
    defparam M_this_state_q_2_LC_15_16_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_15_16_5.LUT_INIT=16'b1110101011000000;
    LogicCell40 M_this_state_q_2_LC_15_16_5 (
            .in0(N__21492),
            .in1(N__16898),
            .in2(N__16221),
            .in3(N__27607),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34561),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_LC_15_17_1.C_ON=1'b0;
    defparam M_this_substate_q_LC_15_17_1.SEQ_MODE=4'b1000;
    defparam M_this_substate_q_LC_15_17_1.LUT_INIT=16'b1110110010101010;
    LogicCell40 M_this_substate_q_LC_15_17_1 (
            .in0(N__16218),
            .in1(N__16928),
            .in2(N__17610),
            .in3(N__17858),
            .lcout(M_this_substate_qZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34568),
            .ce(),
            .sr(N__34990));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_i_1_6_LC_15_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_i_1_6_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_i_1_6_LC_15_17_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_i_1_6_LC_15_17_7  (
            .in0(N__17832),
            .in1(N__17755),
            .in2(_gnd_net_),
            .in3(N__17671),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_15_18_7 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_15_18_7 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_15_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16203),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34575),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_3_LC_15_25_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_3_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_3_LC_15_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_3_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(N__33730),
            .in2(_gnd_net_),
            .in3(N__17385),
            .lcout(M_this_map_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_2_LC_15_25_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_2_LC_15_25_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_2_LC_15_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_2_LC_15_25_6  (
            .in0(_gnd_net_),
            .in1(N__33845),
            .in2(_gnd_net_),
            .in3(N__17384),
            .lcout(M_this_map_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_16_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_16_9_4 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_16_9_4  (
            .in0(N__16141),
            .in1(N__16105),
            .in2(N__16048),
            .in3(N__15909),
            .lcout(\this_vga_signals.M_vcounter_d7lt8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_16_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_16_10_0 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_16_10_0  (
            .in0(N__16716),
            .in1(N__16791),
            .in2(N__16803),
            .in3(N__16418),
            .lcout(\this_vga_signals.M_vcounter_d8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_16_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_16_10_1 .LUT_INIT=16'b0000000100001111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_16_10_1  (
            .in0(N__16790),
            .in1(N__16717),
            .in2(N__16627),
            .in3(N__16516),
            .lcout(\this_vga_signals.un4_lvisibility_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_16_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_16_10_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_16_10_2  (
            .in0(N__16868),
            .in1(N__17146),
            .in2(_gnd_net_),
            .in3(N__16419),
            .lcout(\this_vga_signals.line_clk_1 ),
            .ltout(\this_vga_signals.line_clk_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICHRV3_7_LC_16_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICHRV3_7_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICHRV3_7_LC_16_10_3 .LUT_INIT=16'b1011000011010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICHRV3_7_LC_16_10_3  (
            .in0(N__16355),
            .in1(N__16341),
            .in2(N__16362),
            .in3(N__16270),
            .lcout(M_this_vga_signals_line_clk_0),
            .ltout(M_this_vga_signals_line_clk_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIGL6V4_0_LC_16_10_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIGL6V4_0_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIGL6V4_0_LC_16_10_4 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \this_ppu.M_state_q_RNIGL6V4_0_LC_16_10_4  (
            .in0(N__21576),
            .in1(N__21674),
            .in2(N__16359),
            .in3(N__35083),
            .lcout(\this_ppu.M_state_q_RNIGL6V4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_LC_16_10_5 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_LC_16_10_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.line_clk.M_last_q_LC_16_10_5 .LUT_INIT=16'b1011000011010000;
    LogicCell40 \this_ppu.line_clk.M_last_q_LC_16_10_5  (
            .in0(N__16356),
            .in1(N__16342),
            .in2(N__16287),
            .in3(N__16271),
            .lcout(\this_ppu.M_last_q ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34514),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_1_LC_16_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_1_LC_16_10_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_1_LC_16_10_6 .LUT_INIT=16'b0101011100001000;
    LogicCell40 \this_vga_signals.M_lcounter_q_1_LC_16_10_6  (
            .in0(N__17283),
            .in1(N__16839),
            .in2(N__17015),
            .in3(N__17147),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34514),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_1_LC_16_11_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_1_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_1_LC_16_11_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_1_LC_16_11_3  (
            .in0(N__29792),
            .in1(N__29951),
            .in2(_gnd_net_),
            .in3(N__20723),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34520),
            .ce(),
            .sr(N__19139));
    defparam \this_ppu.M_haddress_q_0_LC_16_11_7 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_0_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_0_LC_16_11_7 .LUT_INIT=16'b0000110111110010;
    LogicCell40 \this_ppu.M_haddress_q_0_LC_16_11_7  (
            .in0(N__21078),
            .in1(N__21114),
            .in2(N__31503),
            .in3(N__29950),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34520),
            .ce(),
            .sr(N__19139));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(N__16869),
            .in2(_gnd_net_),
            .in3(N__17118),
            .lcout(\this_vga_signals.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_10_LC_16_13_1.C_ON=1'b0;
    defparam M_this_state_q_10_LC_16_13_1.SEQ_MODE=4'b1000;
    defparam M_this_state_q_10_LC_16_13_1.LUT_INIT=16'b1101000000010000;
    LogicCell40 M_this_state_q_10_LC_16_13_1 (
            .in0(N__16971),
            .in1(N__23222),
            .in2(N__21444),
            .in3(N__27549),
            .lcout(M_this_state_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34530),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_16_13_4 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_16_13_4 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_16_13_4 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_16_13_4  (
            .in0(N__16830),
            .in1(N__16820),
            .in2(_gnd_net_),
            .in3(N__35071),
            .lcout(this_pixel_clk_M_counter_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34530),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.G_425_LC_16_13_6 .C_ON=1'b0;
    defparam \this_ppu.G_425_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.G_425_LC_16_13_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_ppu.G_425_LC_16_13_6  (
            .in0(N__16829),
            .in1(N__16819),
            .in2(_gnd_net_),
            .in3(N__35070),
            .lcout(G_425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_1_1_LC_16_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_1_1_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_1_1_LC_16_14_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_1_1_LC_16_14_3  (
            .in0(N__27550),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35079),
            .lcout(\this_vga_signals.N_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_o2_8_LC_16_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_o2_8_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_o2_8_LC_16_14_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_i_o2_8_LC_16_14_5  (
            .in0(N__23431),
            .in1(N__23148),
            .in2(_gnd_net_),
            .in3(N__21729),
            .lcout(),
            .ltout(\this_vga_signals.N_152_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_8_LC_16_14_6.C_ON=1'b0;
    defparam M_this_state_q_8_LC_16_14_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_8_LC_16_14_6.LUT_INIT=16'b0001000101010000;
    LogicCell40 M_this_state_q_8_LC_16_14_6 (
            .in0(N__35080),
            .in1(N__27551),
            .in2(N__16806),
            .in3(N__22928),
            .lcout(M_this_state_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34536),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_3_LC_16_15_0.C_ON=1'b0;
    defparam M_this_state_q_3_LC_16_15_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_16_15_0.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_3_LC_16_15_0 (
            .in0(N__16899),
            .in1(N__21469),
            .in2(N__17448),
            .in3(N__24422),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34544),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_2_0_LC_16_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_2_0_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_2_0_LC_16_15_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_0_a2_2_0_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__24421),
            .in2(_gnd_net_),
            .in3(N__28914),
            .lcout(\this_vga_signals.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_16_15_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_16_15_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_sprites_ram.mem_mem_4_0_wclke_3_LC_16_15_3  (
            .in0(N__30318),
            .in1(N__30239),
            .in2(N__30162),
            .in3(N__30048),
            .lcout(\this_sprites_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_16_15_5.C_ON=1'b0;
    defparam M_this_state_q_4_LC_16_15_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_16_15_5.LUT_INIT=16'b1110101011000000;
    LogicCell40 M_this_state_q_4_LC_16_15_5 (
            .in0(N__21470),
            .in1(N__16900),
            .in2(N__16878),
            .in3(N__25225),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34544),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_1_10_LC_16_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_1_10_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_1_10_LC_16_15_6 .LUT_INIT=16'b0001111100010101;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_i_1_10_LC_16_15_6  (
            .in0(N__20899),
            .in1(N__27537),
            .in2(N__22992),
            .in3(N__21728),
            .lcout(\this_vga_signals.M_this_state_q_srsts_i_i_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_15_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_15_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_15_7  (
            .in0(N__30317),
            .in1(N__30238),
            .in2(N__30161),
            .in3(N__30047),
            .lcout(\this_sprites_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_3_sn_m2_LC_16_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_3_sn_m2_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_3_sn_m2_LC_16_16_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_3_sn_m2_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__27584),
            .in2(_gnd_net_),
            .in3(N__22881),
            .lcout(N_383_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_16_16_2.C_ON=1'b0;
    defparam M_this_state_q_1_LC_16_16_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_16_16_2.LUT_INIT=16'b1110101011000000;
    LogicCell40 M_this_state_q_1_LC_16_16_2 (
            .in0(N__21483),
            .in1(N__16901),
            .in2(N__16932),
            .in3(N__22882),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34552),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_16_16_4.C_ON=1'b0;
    defparam M_this_state_q_6_LC_16_16_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_16_16_4.LUT_INIT=16'b1111100010001000;
    LogicCell40 M_this_state_q_6_LC_16_16_4 (
            .in0(N__21484),
            .in1(N__23315),
            .in2(N__16917),
            .in3(N__16902),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34552),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_i_1_4_LC_16_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_i_1_4_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_i_1_4_LC_16_16_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_i_1_4_LC_16_16_6  (
            .in0(N__17831),
            .in1(N__17757),
            .in2(_gnd_net_),
            .in3(N__17670),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_11_LC_16_16_7.C_ON=1'b0;
    defparam M_this_state_q_11_LC_16_16_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_11_LC_16_16_7.LUT_INIT=16'b1010000011100000;
    LogicCell40 M_this_state_q_11_LC_16_16_7 (
            .in0(N__23203),
            .in1(N__20901),
            .in2(N__17457),
            .in3(N__21730),
            .lcout(M_this_state_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34552),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_d_4_sqmuxa_0_a3_0_a2_0_LC_16_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_d_4_sqmuxa_0_a3_0_a2_0_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_d_4_sqmuxa_0_a3_0_a2_0_LC_16_17_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_data_count_d_4_sqmuxa_0_a3_0_a2_0_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__22991),
            .in2(_gnd_net_),
            .in3(N__27519),
            .lcout(N_164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_1_11_LC_16_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_1_11_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_1_11_LC_16_17_7 .LUT_INIT=16'b0000000001110010;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_1_11_LC_16_17_7  (
            .in0(N__23202),
            .in1(N__27520),
            .in2(N__23433),
            .in3(N__35089),
            .lcout(\this_vga_signals.M_this_state_q_srsts_i_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0_3_LC_16_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0_3_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0_3_LC_16_18_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0_3_LC_16_18_0  (
            .in0(N__17822),
            .in1(N__17756),
            .in2(_gnd_net_),
            .in3(N__17658),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_en_0_a3_0_LC_16_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_en_0_a3_0_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_en_0_a3_0_LC_16_19_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_en_0_a3_0_LC_16_19_0  (
            .in0(N__23210),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27536),
            .lcout(M_this_state_d_0_sqmuxa_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_7_LC_16_25_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_7_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_7_LC_16_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_7_LC_16_25_0  (
            .in0(_gnd_net_),
            .in1(N__35226),
            .in2(_gnd_net_),
            .in3(N__17375),
            .lcout(M_this_map_ram_write_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_32_3.C_ON=1'b0;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_32_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_32_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_32_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35076),
            .lcout(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_17_8_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_17_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_17_8_6  (
            .in0(N__17133),
            .in1(N__17272),
            .in2(_gnd_net_),
            .in3(N__17093),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_7_LC_17_9_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_7_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_7_LC_17_9_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_haddress_q_7_LC_17_9_1  (
            .in0(N__20454),
            .in1(N__20528),
            .in2(N__20401),
            .in3(N__18909),
            .lcout(M_this_ppu_map_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(N__19141));
    defparam \this_ppu.M_haddress_q_5_LC_17_10_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_5_LC_17_10_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_5_LC_17_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_haddress_q_5_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__20527),
            .in2(_gnd_net_),
            .in3(N__18907),
            .lcout(M_this_ppu_map_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34523),
            .ce(),
            .sr(N__19140));
    defparam \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_10_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_10_6  (
            .in0(N__17148),
            .in1(N__17132),
            .in2(_gnd_net_),
            .in3(N__17094),
            .lcout(\this_vga_signals.un1_M_hcounter_d7_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_2_LC_17_11_6.C_ON=1'b0;
    defparam M_this_data_count_q_2_LC_17_11_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_17_11_6.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_2_LC_17_11_6 (
            .in0(N__19293),
            .in1(N__19461),
            .in2(_gnd_net_),
            .in3(N__19315),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34526),
            .ce(N__19401),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_17_12_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_17_12_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_17_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_17_12_4  (
            .in0(N__34780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34532),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_5_LC_17_13_5.C_ON=1'b0;
    defparam M_this_data_count_q_5_LC_17_13_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_17_13_5.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_5_LC_17_13_5 (
            .in0(N__19456),
            .in1(N__19227),
            .in2(_gnd_net_),
            .in3(N__21301),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34539),
            .ce(N__19394),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_LC_17_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_LC_17_14_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_data_count_qlde_i_o2_LC_17_14_1  (
            .in0(N__21721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23430),
            .lcout(),
            .ltout(\this_vga_signals.N_153_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qlde_i_i_LC_17_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qlde_i_i_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qlde_i_i_LC_17_14_2 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \this_vga_signals.M_this_data_count_qlde_i_i_LC_17_14_2  (
            .in0(N__35084),
            .in1(N__35261),
            .in2(N__17463),
            .in3(N__17502),
            .lcout(M_this_data_count_qlde_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_9_8_LC_17_14_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_9_8_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_9_8_LC_17_14_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_9_8_LC_17_14_3  (
            .in0(N__19316),
            .in1(N__19342),
            .in2(N__19271),
            .in3(N__19360),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_17_14_4.C_ON=1'b0;
    defparam M_this_data_count_q_0_LC_17_14_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_17_14_4.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_0_LC_17_14_4 (
            .in0(N__19361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19446),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34547),
            .ce(N__19393),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_686_i_LC_17_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.N_686_i_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_686_i_LC_17_14_5 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \this_vga_signals.N_686_i_LC_17_14_5  (
            .in0(N__21722),
            .in1(N__23253),
            .in2(_gnd_net_),
            .in3(N__35085),
            .lcout(N_686_i),
            .ltout(N_686_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_1_LC_17_14_6.C_ON=1'b0;
    defparam M_this_data_count_q_1_LC_17_14_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_17_14_6.LUT_INIT=16'b0000101000000101;
    LogicCell40 M_this_data_count_q_1_LC_17_14_6 (
            .in0(N__19343),
            .in1(_gnd_net_),
            .in2(N__17460),
            .in3(N__19329),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34547),
            .ce(N__19393),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_10_LC_17_15_0.C_ON=1'b0;
    defparam M_this_data_count_q_10_LC_17_15_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_17_15_0.LUT_INIT=16'b0100010011100100;
    LogicCell40 M_this_data_count_q_10_LC_17_15_0 (
            .in0(N__19454),
            .in1(N__20160),
            .in2(N__17550),
            .in3(N__35096),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34555),
            .ce(N__19395),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_6_8_LC_17_15_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_6_8_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_6_8_LC_17_15_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_6_8_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__19183),
            .in2(_gnd_net_),
            .in3(N__19211),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_8_LC_17_15_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_8_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_8_LC_17_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_8_8_LC_17_15_3  (
            .in0(N__20113),
            .in1(N__20143),
            .in2(N__19514),
            .in3(N__20171),
            .lcout(),
            .ltout(\this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_LC_17_15_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_LC_17_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_8_LC_17_15_4  (
            .in0(N__17517),
            .in1(N__21240),
            .in2(N__17511),
            .in3(N__17508),
            .lcout(N_848),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_12_LC_17_15_5.C_ON=1'b0;
    defparam M_this_data_count_q_12_LC_17_15_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_17_15_5.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_12_LC_17_15_5 (
            .in0(N__20114),
            .in1(N__19524),
            .in2(_gnd_net_),
            .in3(N__19452),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34555),
            .ce(N__19395),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_6_LC_17_15_6.C_ON=1'b0;
    defparam M_this_data_count_q_6_LC_17_15_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_17_15_6.LUT_INIT=16'b0100010011100100;
    LogicCell40 M_this_data_count_q_6_LC_17_15_6 (
            .in0(N__19455),
            .in1(N__19200),
            .in2(N__26499),
            .in3(N__35097),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34555),
            .ce(N__19395),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_7_LC_17_15_7.C_ON=1'b0;
    defparam M_this_data_count_q_7_LC_17_15_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_17_15_7.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_7_LC_17_15_7 (
            .in0(N__19170),
            .in1(N__19453),
            .in2(_gnd_net_),
            .in3(N__19184),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34555),
            .ce(N__19395),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_0_LC_17_16_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_0_LC_17_16_0.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_0_LC_17_16_0.LUT_INIT=16'b0010001100100000;
    LogicCell40 M_this_sprites_address_q_0_LC_17_16_0 (
            .in0(N__23760),
            .in1(N__29111),
            .in2(N__28946),
            .in3(N__19485),
            .lcout(M_this_sprites_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34562),
            .ce(),
            .sr(N__28660));
    defparam \this_vga_signals.N_444_i_i_a2_LC_17_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.N_444_i_i_a2_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_444_i_i_a2_LC_17_16_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.N_444_i_i_a2_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__17501),
            .in2(_gnd_net_),
            .in3(N__21720),
            .lcout(\this_vga_signals.N_154 ),
            .ltout(\this_vga_signals.N_154_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_3_0_LC_17_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_3_0_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_3_0_LC_17_16_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_3_0_LC_17_16_5  (
            .in0(N__17606),
            .in1(N__18377),
            .in2(N__17478),
            .in3(N__34695),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_0_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_5_LC_17_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_5_LC_17_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_5_LC_17_17_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_ppu.M_state_q_5_LC_17_17_0  (
            .in0(N__35091),
            .in1(N__20367),
            .in2(_gnd_net_),
            .in3(N__20325),
            .lcout(\this_ppu.M_state_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34569),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0_0_LC_17_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0_0_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0_0_LC_17_17_1 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0_0_LC_17_17_1  (
            .in0(N__18384),
            .in1(N__27521),
            .in2(N__17879),
            .in3(N__35090),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_0_LC_17_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_0_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_0_LC_17_17_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_0_LC_17_17_2  (
            .in0(N__17906),
            .in1(N__23361),
            .in2(N__26540),
            .in3(N__18366),
            .lcout(),
            .ltout(\this_vga_signals.N_62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_17_17_3.C_ON=1'b0;
    defparam M_this_state_q_0_LC_17_17_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_0_LC_17_17_3.LUT_INIT=16'b0000101000001111;
    LogicCell40 M_this_state_q_0_LC_17_17_3 (
            .in0(N__18360),
            .in1(_gnd_net_),
            .in2(N__18354),
            .in3(N__18351),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34569),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI43UU_0_6_LC_17_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI43UU_0_6_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI43UU_0_6_LC_17_17_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \this_ppu.M_state_q_RNI43UU_0_6_LC_17_17_4  (
            .in0(N__18345),
            .in1(N__32010),
            .in2(N__31667),
            .in3(N__31452),
            .lcout(M_this_ppu_sprites_addr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI43UU_1_6_LC_17_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI43UU_1_6_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI43UU_1_6_LC_17_17_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \this_ppu.M_state_q_RNI43UU_1_6_LC_17_17_5  (
            .in0(N__31453),
            .in1(N__18117),
            .in2(N__31986),
            .in3(N__31642),
            .lcout(M_this_ppu_sprites_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_substate_d_0_sqmuxa_0_a3_0_a2_0_LC_17_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_substate_d_0_sqmuxa_0_a3_0_a2_0_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_substate_d_0_sqmuxa_0_a3_0_a2_0_LC_17_17_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.M_this_substate_d_0_sqmuxa_0_a3_0_a2_0_LC_17_17_6  (
            .in0(N__17907),
            .in1(N__17872),
            .in2(N__26541),
            .in3(N__23360),
            .lcout(N_84),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_m2_0_LC_17_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_m2_0_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_m2_0_LC_17_19_1 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_0_m2_0_LC_17_19_1  (
            .in0(N__17815),
            .in1(N__17737),
            .in2(_gnd_net_),
            .in3(N__17645),
            .lcout(N_36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI01PG1_1_LC_17_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI01PG1_1_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI01PG1_1_LC_17_19_4 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \this_ppu.M_state_q_RNI01PG1_1_LC_17_19_4  (
            .in0(N__21011),
            .in1(N__18456),
            .in2(_gnd_net_),
            .in3(N__35086),
            .lcout(\this_ppu.N_1156_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIE07J4_0_1_LC_17_19_6.C_ON=1'b0;
    defparam M_this_state_q_RNIE07J4_0_1_LC_17_19_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIE07J4_0_1_LC_17_19_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 M_this_state_q_RNIE07J4_0_1_LC_17_19_6 (
            .in0(N__21384),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(port_dmab_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_2_LC_17_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_2_LC_17_20_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_2_LC_17_20_0 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \this_ppu.M_oam_idx_q_2_LC_17_20_0  (
            .in0(N__18420),
            .in1(N__18995),
            .in2(N__19046),
            .in3(N__18410),
            .lcout(M_this_ppu_oam_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34589),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIGJUB2_3_LC_17_20_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIGJUB2_3_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIGJUB2_3_LC_17_20_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_state_q_RNIGJUB2_3_LC_17_20_1  (
            .in0(N__20361),
            .in1(N__18937),
            .in2(_gnd_net_),
            .in3(N__20319),
            .lcout(\this_ppu.un1_M_oam_idx_q_1_c1 ),
            .ltout(\this_ppu.un1_M_oam_idx_q_1_c1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_17_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_17_20_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__19038),
            .in2(N__18462),
            .in3(N__18993),
            .lcout(\this_ppu.un1_M_oam_idx_q_1_c3 ),
            .ltout(\this_ppu.un1_M_oam_idx_q_1_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_3_LC_17_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_3_LC_17_20_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_3_LC_17_20_3 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \this_ppu.M_oam_idx_q_3_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__20838),
            .in2(N__18459),
            .in3(N__18405),
            .lcout(M_this_ppu_oam_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34589),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_2_LC_17_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_2_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_2_LC_17_20_5 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \this_ppu.M_state_q_RNO_0_2_LC_17_20_5  (
            .in0(N__20362),
            .in1(N__21016),
            .in2(_gnd_net_),
            .in3(N__18455),
            .lcout(\this_ppu.N_148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_4_LC_17_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_4_LC_17_20_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_4_LC_17_20_6 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \this_ppu.M_oam_idx_q_4_LC_17_20_6  (
            .in0(N__18406),
            .in1(N__18968),
            .in2(N__20846),
            .in3(N__18426),
            .lcout(\this_ppu.M_oam_idx_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34589),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_1_LC_17_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_1_LC_17_20_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_1_LC_17_20_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_oam_idx_q_1_LC_17_20_7  (
            .in0(N__18994),
            .in1(N__18404),
            .in2(_gnd_net_),
            .in3(N__18419),
            .lcout(M_this_ppu_oam_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34589),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_0_LC_17_21_2 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_0_LC_17_21_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_0_LC_17_21_2 .LUT_INIT=16'b1010000000101000;
    LogicCell40 \this_ppu.M_oam_idx_q_0_LC_17_21_2  (
            .in0(N__18411),
            .in1(N__20366),
            .in2(N__18941),
            .in3(N__20324),
            .lcout(M_this_ppu_oam_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34595),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_RNI3VF_4_LC_17_21_3 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_RNI3VF_4_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_idx_q_RNI3VF_4_LC_17_21_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_ppu.M_oam_idx_q_RNI3VF_4_LC_17_21_3  (
            .in0(N__19045),
            .in1(N__18992),
            .in2(N__18969),
            .in3(N__18933),
            .lcout(\this_ppu.N_144_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_6_LC_18_9_7 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_6_LC_18_9_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_6_LC_18_9_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_6_LC_18_9_7  (
            .in0(N__20453),
            .in1(N__20529),
            .in2(_gnd_net_),
            .in3(N__18908),
            .lcout(M_this_ppu_map_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34524),
            .ce(),
            .sr(N__19155));
    defparam \this_ppu.M_haddress_q_RNIRHU1G_1_LC_18_10_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIRHU1G_1_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIRHU1G_1_LC_18_10_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNIRHU1G_1_LC_18_10_0  (
            .in0(N__29826),
            .in1(N__29961),
            .in2(_gnd_net_),
            .in3(N__20715),
            .lcout(\this_ppu.un1_M_haddress_q_3_c2 ),
            .ltout(\this_ppu.un1_M_haddress_q_3_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI81A2G_4_LC_18_10_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI81A2G_4_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI81A2G_4_LC_18_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNI81A2G_4_LC_18_10_1  (
            .in0(N__20597),
            .in1(N__20230),
            .in2(N__18912),
            .in3(N__29726),
            .lcout(\this_ppu.un1_M_haddress_q_3_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_10_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_10_5  (
            .in0(N__18891),
            .in1(N__18873),
            .in2(_gnd_net_),
            .in3(N__29630),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_6_LC_18_10_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_6_LC_18_10_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_6_LC_18_10_6 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \this_ppu.M_state_q_6_LC_18_10_6  (
            .in0(N__34721),
            .in1(N__20781),
            .in2(N__21087),
            .in3(N__21110),
            .lcout(\this_ppu.M_state_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34527),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_2_LC_18_11_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_2_LC_18_11_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_2_LC_18_11_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_haddress_q_2_LC_18_11_1  (
            .in0(N__29949),
            .in1(N__29804),
            .in2(N__29742),
            .in3(N__20722),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34533),
            .ce(),
            .sr(N__19154));
    defparam \this_ppu.M_haddress_q_RNI88B5_0_LC_18_11_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI88B5_0_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI88B5_0_LC_18_11_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_ppu.M_haddress_q_RNI88B5_0_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__29896),
            .in2(_gnd_net_),
            .in3(N__29947),
            .lcout(),
            .ltout(\this_ppu.un2_hscroll_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIVK7O_0_LC_18_11_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIVK7O_0_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIVK7O_0_LC_18_11_5 .LUT_INIT=16'b1010101010001011;
    LogicCell40 \this_ppu.M_haddress_q_RNIVK7O_0_LC_18_11_5  (
            .in0(N__29948),
            .in1(N__31552),
            .in2(N__18861),
            .in3(N__31480),
            .lcout(M_this_ppu_sprites_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_3_LC_18_11_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_3_LC_18_11_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_3_LC_18_11_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_3_LC_18_11_6  (
            .in0(N__20231),
            .in1(N__29727),
            .in2(_gnd_net_),
            .in3(N__19163),
            .lcout(M_this_ppu_map_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34533),
            .ce(),
            .sr(N__19154));
    defparam \this_ppu.M_haddress_q_4_LC_18_11_7 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_4_LC_18_11_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_4_LC_18_11_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_haddress_q_4_LC_18_11_7  (
            .in0(N__19164),
            .in1(N__20598),
            .in2(N__29743),
            .in3(N__20232),
            .lcout(M_this_ppu_map_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34533),
            .ce(),
            .sr(N__19154));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_12_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_12_0  (
            .in0(N__29628),
            .in1(N__19116),
            .in2(_gnd_net_),
            .in3(N__19101),
            .lcout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_18_12_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_18_12_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_wclke_3_LC_18_12_5  (
            .in0(N__30243),
            .in1(N__30294),
            .in2(N__30157),
            .in3(N__30054),
            .lcout(\this_sprites_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_3_LC_18_13_5.C_ON=1'b0;
    defparam M_this_data_count_q_3_LC_18_13_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_18_13_5.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_3_LC_18_13_5 (
            .in0(N__19248),
            .in1(N__19457),
            .in2(_gnd_net_),
            .in3(N__19270),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34548),
            .ce(N__19397),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_4_LC_18_14_1.C_ON=1'b0;
    defparam M_this_data_count_q_4_LC_18_14_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_18_14_1.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_4_LC_18_14_1 (
            .in0(N__19449),
            .in1(N__19236),
            .in2(_gnd_net_),
            .in3(N__21258),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34556),
            .ce(N__19396),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_9_LC_18_14_2.C_ON=1'b0;
    defparam M_this_data_count_q_9_LC_18_14_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_18_14_2.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_9_LC_18_14_2 (
            .in0(N__20184),
            .in1(N__19451),
            .in2(_gnd_net_),
            .in3(N__21280),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34556),
            .ce(N__19396),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_11_LC_18_14_4.C_ON=1'b0;
    defparam M_this_data_count_q_11_LC_18_14_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_18_14_4.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_11_LC_18_14_4 (
            .in0(N__20127),
            .in1(N__19447),
            .in2(_gnd_net_),
            .in3(N__20147),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34556),
            .ce(N__19396),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_18_14_5.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_18_14_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_18_14_5.LUT_INIT=16'b1110010001000100;
    LogicCell40 M_this_data_count_q_13_LC_18_14_5 (
            .in0(N__19448),
            .in1(N__19494),
            .in2(N__22839),
            .in3(N__25245),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34556),
            .ce(N__19396),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_8_LC_18_14_7.C_ON=1'b0;
    defparam M_this_data_count_q_8_LC_18_14_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_18_14_7.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_8_LC_18_14_7 (
            .in0(N__19450),
            .in1(N__20196),
            .in2(_gnd_net_),
            .in3(N__21332),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34556),
            .ce(N__19396),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_c_0_LC_18_15_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_c_0_LC_18_15_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_c_0_LC_18_15_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 M_this_data_count_q_cry_c_0_LC_18_15_0 (
            .in0(_gnd_net_),
            .in1(N__19362),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(M_this_data_count_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_18_15_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_18_15_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_18_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_0_THRU_LUT4_0_LC_18_15_1 (
            .in0(_gnd_net_),
            .in1(N__19841),
            .in2(N__19347),
            .in3(N__19323),
            .lcout(M_this_data_count_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_0),
            .carryout(M_this_data_count_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_18_15_2.C_ON=1'b1;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_18_15_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_18_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_1_THRU_LUT4_0_LC_18_15_2 (
            .in0(_gnd_net_),
            .in1(N__19320),
            .in2(N__19911),
            .in3(N__19281),
            .lcout(M_this_data_count_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_1),
            .carryout(M_this_data_count_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_18_15_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_18_15_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_18_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_2_THRU_LUT4_0_LC_18_15_3 (
            .in0(_gnd_net_),
            .in1(N__19845),
            .in2(N__19278),
            .in3(N__19239),
            .lcout(M_this_data_count_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_2),
            .carryout(M_this_data_count_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_18_15_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_18_15_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_18_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_3_THRU_LUT4_0_LC_18_15_4 (
            .in0(_gnd_net_),
            .in1(N__21257),
            .in2(N__19912),
            .in3(N__19230),
            .lcout(M_this_data_count_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_3),
            .carryout(M_this_data_count_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_18_15_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_18_15_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_18_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_4_THRU_LUT4_0_LC_18_15_5 (
            .in0(_gnd_net_),
            .in1(N__19849),
            .in2(N__21312),
            .in3(N__19215),
            .lcout(M_this_data_count_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_4),
            .carryout(M_this_data_count_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_6_LC_18_15_6.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_6_LC_18_15_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_6_LC_18_15_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_6_LC_18_15_6 (
            .in0(_gnd_net_),
            .in1(N__19212),
            .in2(N__19910),
            .in3(N__19194),
            .lcout(M_this_data_count_q_s_6),
            .ltout(),
            .carryin(M_this_data_count_q_cry_5),
            .carryout(M_this_data_count_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_18_15_7.C_ON=1'b1;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_18_15_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_18_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_6_THRU_LUT4_0_LC_18_15_7 (
            .in0(_gnd_net_),
            .in1(N__19850),
            .in2(N__19191),
            .in3(N__20199),
            .lcout(M_this_data_count_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_6),
            .carryout(M_this_data_count_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_7_THRU_LUT4_0_LC_18_16_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_7_THRU_LUT4_0_LC_18_16_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_7_THRU_LUT4_0_LC_18_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_7_THRU_LUT4_0_LC_18_16_0 (
            .in0(_gnd_net_),
            .in1(N__21333),
            .in2(N__19837),
            .in3(N__20187),
            .lcout(M_this_data_count_q_cry_7_THRU_CO),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(M_this_data_count_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_18_16_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_18_16_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_18_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_8_THRU_LUT4_0_LC_18_16_1 (
            .in0(_gnd_net_),
            .in1(N__19765),
            .in2(N__21285),
            .in3(N__20175),
            .lcout(M_this_data_count_q_cry_8_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_8),
            .carryout(M_this_data_count_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_10_LC_18_16_2.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_10_LC_18_16_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_10_LC_18_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_10_LC_18_16_2 (
            .in0(_gnd_net_),
            .in1(N__20172),
            .in2(N__19835),
            .in3(N__20154),
            .lcout(M_this_data_count_q_s_10),
            .ltout(),
            .carryin(M_this_data_count_q_cry_9),
            .carryout(M_this_data_count_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_18_16_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_18_16_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_18_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_10_THRU_LUT4_0_LC_18_16_3 (
            .in0(_gnd_net_),
            .in1(N__19758),
            .in2(N__20151),
            .in3(N__20118),
            .lcout(M_this_data_count_q_cry_10_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_10),
            .carryout(M_this_data_count_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_18_16_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_18_16_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_18_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_11_THRU_LUT4_0_LC_18_16_4 (
            .in0(_gnd_net_),
            .in1(N__20115),
            .in2(N__19836),
            .in3(N__19518),
            .lcout(M_this_data_count_q_cry_11_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_11),
            .carryout(M_this_data_count_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_13_LC_18_16_5.C_ON=1'b0;
    defparam M_this_data_count_q_RNO_0_13_LC_18_16_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_13_LC_18_16_5.LUT_INIT=16'b1100110000110011;
    LogicCell40 M_this_data_count_q_RNO_0_13_LC_18_16_5 (
            .in0(_gnd_net_),
            .in1(N__19515),
            .in2(_gnd_net_),
            .in3(N__19497),
            .lcout(M_this_data_count_q_s_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_0_LC_18_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_0_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_0_LC_18_16_7 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_0_LC_18_16_7  (
            .in0(N__23801),
            .in1(N__34173),
            .in2(N__27667),
            .in3(N__27554),
            .lcout(N_49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNILG0GD_0_LC_18_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNILG0GD_0_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNILG0GD_0_LC_18_17_3 .LUT_INIT=16'b1011111110101010;
    LogicCell40 \this_ppu.M_state_q_RNILG0GD_0_LC_18_17_3  (
            .in0(N__35081),
            .in1(N__21371),
            .in2(N__19479),
            .in3(N__21549),
            .lcout(\this_ppu.M_state_q_RNILG0GDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIPG425_1_LC_18_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIPG425_1_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIPG425_1_LC_18_17_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIPG425_1_LC_18_17_6  (
            .in0(N__21550),
            .in1(N__30683),
            .in2(_gnd_net_),
            .in3(N__30821),
            .lcout(\this_ppu.un1_M_vaddress_q_2_c2 ),
            .ltout(\this_ppu.un1_M_vaddress_q_2_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_18_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_18_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_18_17_7  (
            .in0(N__21892),
            .in1(N__21933),
            .in2(N__20286),
            .in3(N__30631),
            .lcout(\this_ppu.un1_M_vaddress_q_2_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_5_LC_18_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_5_LC_18_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_5_LC_18_18_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_ppu.M_vaddress_q_5_LC_18_18_4  (
            .in0(N__20282),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21843),
            .lcout(M_this_ppu_map_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34582),
            .ce(),
            .sr(N__21981));
    defparam \this_ppu.M_vaddress_q_7_LC_18_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_7_LC_18_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_7_LC_18_18_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \this_ppu.M_vaddress_q_7_LC_18_18_5  (
            .in0(N__21845),
            .in1(N__20281),
            .in2(N__21809),
            .in3(N__22124),
            .lcout(M_this_ppu_map_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34582),
            .ce(),
            .sr(N__21981));
    defparam \this_ppu.M_vaddress_q_6_LC_18_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_6_LC_18_18_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_6_LC_18_18_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_vaddress_q_6_LC_18_18_6  (
            .in0(N__20283),
            .in1(N__21802),
            .in2(_gnd_net_),
            .in3(N__21844),
            .lcout(M_this_ppu_map_addr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34582),
            .ce(),
            .sr(N__21981));
    defparam \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_18_19_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_18_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__22080),
            .in2(N__29901),
            .in3(N__29965),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_0 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_18_19_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_18_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__22068),
            .in2(N__31794),
            .in3(N__29820),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_0 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_18_19_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_18_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__31835),
            .in2(N__22056),
            .in3(N__29734),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_1 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_18_19_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_18_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__22037),
            .in2(N__24924),
            .in3(N__20248),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_0 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_2 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_18_19_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_18_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__22022),
            .in2(N__20343),
            .in3(N__20614),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_3 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_18_19_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_18_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__22007),
            .in2(N__20298),
            .in3(N__20545),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_4 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_18_19_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_18_19_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_18_19_6  (
            .in0(N__20467),
            .in1(N__22281),
            .in2(N__30897),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_3 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_5 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_18_19_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_18_19_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_18_19_7  (
            .in0(N__20411),
            .in1(N__24885),
            .in2(N__22269),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_4 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_6 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_18_20_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_18_20_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_18_20_0  (
            .in0(N__22101),
            .in1(N__22251),
            .in2(_gnd_net_),
            .in3(N__20370),
            .lcout(\this_ppu.vscroll8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_3_LC_18_20_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_3_LC_18_20_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_3_LC_18_20_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_3_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__20868),
            .in2(_gnd_net_),
            .in3(N__35094),
            .lcout(\this_ppu.M_state_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34596),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc1_LC_18_20_3 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc1_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc1_LC_18_20_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc1_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__31021),
            .in2(_gnd_net_),
            .in3(N__30944),
            .lcout(\this_ppu.un1_M_haddress_q_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_2_LC_18_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_2_LC_18_20_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_2_LC_18_20_5 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \this_ppu.M_state_q_2_LC_18_20_5  (
            .in0(N__20331),
            .in1(N__20323),
            .in2(N__21024),
            .in3(N__35093),
            .lcout(\this_ppu.M_state_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34596),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc2_LC_18_20_6 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc2_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc2_LC_18_20_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc2_LC_18_20_6  (
            .in0(N__30945),
            .in1(_gnd_net_),
            .in2(N__31026),
            .in3(N__31068),
            .lcout(\this_ppu.un1_M_haddress_q_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_4_LC_18_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_4_LC_18_20_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_4_LC_18_20_7 .LUT_INIT=16'b0000000010110000;
    LogicCell40 \this_ppu.M_state_q_4_LC_18_20_7  (
            .in0(N__20842),
            .in1(N__20811),
            .in2(N__20799),
            .in3(N__35095),
            .lcout(\this_ppu.M_state_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34596),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_6_LC_18_21_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_6_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_6_LC_18_21_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_ppu.M_state_q_RNO_0_6_LC_18_21_1  (
            .in0(N__20837),
            .in1(N__20810),
            .in2(N__20798),
            .in3(N__35077),
            .lcout(\this_ppu.N_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_7_LC_18_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_7_LC_18_21_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_7_LC_18_21_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_ppu.M_state_q_7_LC_18_21_4  (
            .in0(N__35078),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31671),
            .lcout(\this_ppu.M_state_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34602),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_19_11_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_19_11_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_19_11_0 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_19_11_0  (
            .in0(N__20769),
            .in1(N__24033),
            .in2(N__23700),
            .in3(N__21228),
            .lcout(M_this_ppu_vram_data_0),
            .ltout(M_this_ppu_vram_data_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vram_en_i_a2_0_LC_19_11_1 .C_ON=1'b0;
    defparam \this_ppu.vram_en_i_a2_0_LC_19_11_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vram_en_i_a2_0_LC_19_11_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.vram_en_i_a2_0_LC_19_11_1  (
            .in0(N__21125),
            .in1(N__22571),
            .in2(N__20742),
            .in3(N__22703),
            .lcout(\this_ppu.N_156 ),
            .ltout(\this_ppu.N_156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI22N1G_5_LC_19_11_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI22N1G_5_LC_19_11_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI22N1G_5_LC_19_11_2 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \this_ppu.M_state_q_RNI22N1G_5_LC_19_11_2  (
            .in0(_gnd_net_),
            .in1(N__31478),
            .in2(N__20739),
            .in3(N__21077),
            .lcout(M_this_ppu_vram_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_11_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_11_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_11_3  (
            .in0(N__29629),
            .in1(N__20697),
            .in2(_gnd_net_),
            .in3(N__20679),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_19_11_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_19_11_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_19_11_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_19_11_4  (
            .in0(N__29633),
            .in1(N__20667),
            .in2(_gnd_net_),
            .in3(N__20652),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_19_11_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_19_11_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_19_11_5 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_19_11_5  (
            .in0(N__22624),
            .in1(N__23691),
            .in2(N__21231),
            .in3(N__26850),
            .lcout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_13_LC_19_11_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_13_LC_19_11_6 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_13_LC_19_11_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \this_sprites_ram.mem_radreg_13_LC_19_11_6  (
            .in0(N__31582),
            .in1(N__31479),
            .in2(N__21222),
            .in3(N__32211),
            .lcout(\this_sprites_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34540),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_12_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_12_1  (
            .in0(N__21198),
            .in1(N__21177),
            .in2(_gnd_net_),
            .in3(N__29632),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_1_LC_19_12_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_19_12_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_19_12_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.M_state_q_RNO_0_1_LC_19_12_2  (
            .in0(N__31481),
            .in1(N__21079),
            .in2(_gnd_net_),
            .in3(N__21548),
            .lcout(\this_ppu.N_150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_12_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_12_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_12_3 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_12_3  (
            .in0(N__23697),
            .in1(N__21159),
            .in2(N__22632),
            .in3(N__21153),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_12_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_12_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_12_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_12_4  (
            .in0(N__23699),
            .in1(N__21147),
            .in2(N__21141),
            .in3(N__20907),
            .lcout(M_this_ppu_vram_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_1_LC_19_12_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_1_LC_19_12_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_1_LC_19_12_5 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \this_ppu.M_state_q_1_LC_19_12_5  (
            .in0(N__21109),
            .in1(N__21093),
            .in2(N__21086),
            .in3(N__34701),
            .lcout(\this_ppu.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34549),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_19_12_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_19_12_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_19_12_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_19_12_7  (
            .in0(N__20940),
            .in1(N__20925),
            .in2(_gnd_net_),
            .in3(N__29631),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIH92S_10_LC_19_13_0.C_ON=1'b0;
    defparam M_this_state_q_RNIH92S_10_LC_19_13_0.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIH92S_10_LC_19_13_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_state_q_RNIH92S_10_LC_19_13_0 (
            .in0(N__24476),
            .in1(N__21756),
            .in2(N__23620),
            .in3(N__20900),
            .lcout(),
            .ltout(M_this_state_q_RNIH92SZ0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI373A1_8_LC_19_13_1.C_ON=1'b0;
    defparam M_this_state_q_RNI373A1_8_LC_19_13_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI373A1_8_LC_19_13_1.LUT_INIT=16'b0000000000110000;
    LogicCell40 M_this_state_q_RNI373A1_8_LC_19_13_1 (
            .in0(_gnd_net_),
            .in1(N__23221),
            .in2(N__21495),
            .in3(N__22938),
            .lcout(M_this_state_q_RNI373A1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_13_LC_19_14_0.C_ON=1'b0;
    defparam M_this_state_q_13_LC_19_14_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_13_LC_19_14_0.LUT_INIT=16'b1111000010000000;
    LogicCell40 M_this_state_q_13_LC_19_14_0 (
            .in0(N__21687),
            .in1(N__23429),
            .in2(N__21491),
            .in3(N__23618),
            .lcout(M_this_state_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34563),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_12_LC_19_14_2.C_ON=1'b0;
    defparam M_this_state_q_12_LC_19_14_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_12_LC_19_14_2.LUT_INIT=16'b1100110011001000;
    LogicCell40 M_this_state_q_12_LC_19_14_2 (
            .in0(N__21686),
            .in1(N__21426),
            .in2(N__23345),
            .in3(N__23619),
            .lcout(M_this_state_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34563),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_7_i_a2_LC_19_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_7_i_a2_LC_19_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_7_i_a2_LC_19_14_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_7_i_a2_LC_19_14_3  (
            .in0(N__22929),
            .in1(N__24433),
            .in2(_gnd_net_),
            .in3(N__25244),
            .lcout(\this_vga_signals.N_485 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_i_o2_7_LC_19_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_i_o2_7_LC_19_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_i_o2_7_LC_19_14_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_a2_0_i_o2_7_LC_19_14_6  (
            .in0(_gnd_net_),
            .in1(N__23428),
            .in2(_gnd_net_),
            .in3(N__35082),
            .lcout(\this_vga_signals.N_94_0 ),
            .ltout(\this_vga_signals.N_94_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_0_12_LC_19_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_0_12_LC_19_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_0_12_LC_19_14_7 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_i_0_12_LC_19_14_7  (
            .in0(N__23617),
            .in1(N__21758),
            .in2(N__21429),
            .in3(N__27514),
            .lcout(\this_vga_signals.M_this_state_q_srsts_i_i_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un21_i_a3_1_1_LC_19_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un21_i_a3_1_1_LC_19_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un21_i_a3_1_1_LC_19_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.un21_i_a3_1_1_LC_19_15_0  (
            .in0(N__24432),
            .in1(N__23139),
            .in2(N__23344),
            .in3(N__27636),
            .lcout(),
            .ltout(this_vga_signals_un21_i_a3_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIE07J4_1_LC_19_15_1.C_ON=1'b0;
    defparam M_this_state_q_RNIE07J4_1_LC_19_15_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIE07J4_1_LC_19_15_1.LUT_INIT=16'b1010101010101000;
    LogicCell40 M_this_state_q_RNIE07J4_1_LC_19_15_1 (
            .in0(N__21420),
            .in1(N__21774),
            .in2(N__21411),
            .in3(N__23106),
            .lcout(port_dmab_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_7_8_LC_19_15_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_7_8_LC_19_15_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_7_8_LC_19_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_7_8_LC_19_15_2  (
            .in0(N__21328),
            .in1(N__21308),
            .in2(N__21281),
            .in3(N__21256),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_a3_0_0_7_LC_19_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a3_0_0_7_LC_19_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a3_0_0_7_LC_19_15_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_a3_0_0_7_LC_19_15_3  (
            .in0(N__23140),
            .in1(N__23432),
            .in2(_gnd_net_),
            .in3(N__24484),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_srsts_i_a3_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_0_7_LC_19_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_0_7_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_0_7_LC_19_15_4 .LUT_INIT=16'b0100010100000101;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_0_7_LC_19_15_4  (
            .in0(N__35092),
            .in1(N__27518),
            .in2(N__21780),
            .in3(N__25233),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_srsts_i_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_19_15_5.C_ON=1'b0;
    defparam M_this_state_q_7_LC_19_15_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_19_15_5.LUT_INIT=16'b1110000011110000;
    LogicCell40 M_this_state_q_7_LC_19_15_5 (
            .in0(N__25234),
            .in1(N__24485),
            .in2(N__21777),
            .in3(N__21732),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34570),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI6Q0S_5_LC_19_15_6.C_ON=1'b0;
    defparam M_this_state_q_RNI6Q0S_5_LC_19_15_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI6Q0S_5_LC_19_15_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_state_q_RNI6Q0S_5_LC_19_15_6 (
            .in0(N__22994),
            .in1(N__23138),
            .in2(N__23343),
            .in3(N__25232),
            .lcout(M_this_state_q_RNI6Q0SZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_o2_12_LC_19_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_o2_12_LC_19_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_o2_12_LC_19_15_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_i_o2_12_LC_19_15_7  (
            .in0(_gnd_net_),
            .in1(N__21757),
            .in2(_gnd_net_),
            .in3(N__21731),
            .lcout(\this_vga_signals.N_93_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_1_LC_19_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_1_LC_19_16_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_1_LC_19_16_2 .LUT_INIT=16'b0111100001111000;
    LogicCell40 \this_ppu.M_vaddress_q_1_LC_19_16_2  (
            .in0(N__30823),
            .in1(N__21551),
            .in2(N__30695),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_vaddress_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34576),
            .ce(),
            .sr(N__21974));
    defparam \this_ppu.M_vaddress_q_0_LC_19_16_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_0_LC_19_16_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_0_LC_19_16_3 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \this_ppu.M_vaddress_q_0_LC_19_16_3  (
            .in0(N__21678),
            .in1(N__21636),
            .in2(N__21603),
            .in3(N__30822),
            .lcout(M_this_ppu_vram_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34576),
            .ce(),
            .sr(N__21974));
    defparam \this_ppu.M_vaddress_q_2_LC_19_16_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_2_LC_19_16_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_2_LC_19_16_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_vaddress_q_2_LC_19_16_4  (
            .in0(N__30824),
            .in1(N__30633),
            .in2(N__30694),
            .in3(N__21552),
            .lcout(\this_ppu.M_vaddress_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34576),
            .ce(),
            .sr(N__21974));
    defparam \this_ppu.M_vaddress_q_3_LC_19_16_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_3_LC_19_16_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_3_LC_19_16_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_vaddress_q_3_LC_19_16_6  (
            .in0(N__21992),
            .in1(N__21934),
            .in2(_gnd_net_),
            .in3(N__30634),
            .lcout(M_this_ppu_map_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34576),
            .ce(),
            .sr(N__21974));
    defparam \this_ppu.M_vaddress_q_4_LC_19_16_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_4_LC_19_16_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_4_LC_19_16_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \this_ppu.M_vaddress_q_4_LC_19_16_7  (
            .in0(N__30632),
            .in1(N__21993),
            .in2(N__21941),
            .in3(N__21893),
            .lcout(M_this_ppu_map_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34576),
            .ce(),
            .sr(N__21974));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_19_17_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_19_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_19_17_0  (
            .in0(_gnd_net_),
            .in1(N__23567),
            .in2(N__30780),
            .in3(N__30812),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_7 ),
            .ltout(),
            .carryin(bfn_19_17_0_),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_19_17_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_19_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_19_17_1  (
            .in0(_gnd_net_),
            .in1(N__23552),
            .in2(N__31899),
            .in3(N__30676),
            .lcout(\this_ppu.M_vaddress_q_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_0 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_19_17_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_19_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_19_17_2  (
            .in0(_gnd_net_),
            .in1(N__23537),
            .in2(N__30597),
            .in3(N__30624),
            .lcout(\this_ppu.M_vaddress_q_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_1 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_19_17_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_19_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_19_17_3  (
            .in0(_gnd_net_),
            .in1(N__23519),
            .in2(N__24936),
            .in3(N__21932),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_5 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_2 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_19_17_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_19_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_19_17_4  (
            .in0(_gnd_net_),
            .in1(N__23501),
            .in2(N__22245),
            .in3(N__21891),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_6 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_3 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_19_17_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_19_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_19_17_5  (
            .in0(_gnd_net_),
            .in1(N__23483),
            .in2(N__33123),
            .in3(N__21842),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_7 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_4 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_19_17_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_19_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_19_17_6  (
            .in0(_gnd_net_),
            .in1(N__23465),
            .in2(N__32910),
            .in3(N__21801),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_8 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_5 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_19_17_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_19_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_19_17_7  (
            .in0(_gnd_net_),
            .in1(N__32094),
            .in2(N__23451),
            .in3(N__22123),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_9 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_6 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_19_18_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_19_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_19_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_19_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22104),
            .lcout(\this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_4_LC_19_18_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_4_LC_19_18_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_4_LC_19_18_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_4_LC_19_18_6  (
            .in0(N__34830),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22092),
            .lcout(\this_reset_cond.M_stage_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34590),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_19_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_19_0  (
            .in0(_gnd_net_),
            .in1(N__22079),
            .in2(N__29897),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_19_19_0_),
            .carryout(\this_ppu.un1_M_haddress_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_19_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_19_1  (
            .in0(_gnd_net_),
            .in1(N__22067),
            .in2(N__31790),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_0 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_19_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_19_2  (
            .in0(_gnd_net_),
            .in1(N__22049),
            .in2(N__31836),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_1 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_19_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_19_3  (
            .in0(_gnd_net_),
            .in1(N__30943),
            .in2(N__22038),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_2 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_19_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_19_4  (
            .in0(_gnd_net_),
            .in1(N__31025),
            .in2(N__22023),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_3 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_19_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_19_5  (
            .in0(_gnd_net_),
            .in1(N__31067),
            .in2(N__22008),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_4 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_19_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_19_6  (
            .in0(_gnd_net_),
            .in1(N__22280),
            .in2(N__30978),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_5 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_19_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_19_7  (
            .in0(_gnd_net_),
            .in1(N__22265),
            .in2(N__24912),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_6 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_19_20_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_19_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_19_20_0 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_19_20_0  (
            .in0(N__32157),
            .in1(N__31914),
            .in2(N__23733),
            .in3(N__22254),
            .lcout(\this_ppu.vscroll8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_4_LC_19_21_6.C_ON=1'b0;
    defparam M_this_oam_address_q_4_LC_19_21_6.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_4_LC_19_21_6.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_4_LC_19_21_6 (
            .in0(N__24853),
            .in1(N__26483),
            .in2(_gnd_net_),
            .in3(N__24833),
            .lcout(M_this_oam_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34605),
            .ce(),
            .sr(N__28657));
    defparam \this_ppu.un1_oam_data_axbxc1_LC_19_25_7 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc1_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc1_LC_19_25_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.un1_oam_data_axbxc1_LC_19_25_7  (
            .in0(_gnd_net_),
            .in1(N__33041),
            .in2(_gnd_net_),
            .in3(N__32966),
            .lcout(\this_ppu.un1_M_vaddress_q_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_20_9_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_20_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_20_9_4  (
            .in0(N__29648),
            .in1(N__22227),
            .in2(_gnd_net_),
            .in3(N__22212),
            .lcout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_9_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_9_7  (
            .in0(N__22194),
            .in1(N__22176),
            .in2(_gnd_net_),
            .in3(N__29649),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_12_LC_20_10_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_12_LC_20_10_2 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_12_LC_20_10_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \this_sprites_ram.mem_radreg_12_LC_20_10_2  (
            .in0(N__31501),
            .in1(N__31578),
            .in2(N__22164),
            .in3(N__32259),
            .lcout(\this_sprites_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34541),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_20_10_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_20_10_3 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_20_10_3  (
            .in0(N__23695),
            .in1(N__24099),
            .in2(N__22628),
            .in3(N__22146),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_10_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_10_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_10_4  (
            .in0(N__23696),
            .in1(N__22722),
            .in2(N__22716),
            .in3(N__29559),
            .lcout(M_this_ppu_vram_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_20_11_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_20_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_20_11_0  (
            .in0(N__22692),
            .in1(N__22674),
            .in2(_gnd_net_),
            .in3(N__29627),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_20_11_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_20_11_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_20_11_1  (
            .in0(N__22659),
            .in1(_gnd_net_),
            .in2(N__29650),
            .in3(N__22647),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_20_11_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_20_11_2 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_20_11_2  (
            .in0(N__23681),
            .in1(N__22620),
            .in2(N__22593),
            .in3(N__22287),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_20_11_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_20_11_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_20_11_3  (
            .in0(N__23698),
            .in1(N__22590),
            .in2(N__22584),
            .in3(N__24069),
            .lcout(M_this_ppu_vram_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI43UU_2_6_LC_20_11_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI43UU_2_6_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI43UU_2_6_LC_20_11_4 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \this_ppu.M_state_q_RNI43UU_2_6_LC_20_11_4  (
            .in0(N__22560),
            .in1(N__31492),
            .in2(N__31663),
            .in3(N__31941),
            .lcout(M_this_ppu_sprites_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_20_11_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_20_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_20_11_7  (
            .in0(N__29623),
            .in1(N__22314),
            .in2(_gnd_net_),
            .in3(N__22299),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_10_LC_20_12_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_10_LC_20_12_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_10_LC_20_12_4.LUT_INIT=16'b0000100000001010;
    LogicCell40 M_this_sprites_address_q_10_LC_20_12_4 (
            .in0(N__24024),
            .in1(N__24153),
            .in2(N__22848),
            .in3(N__29007),
            .lcout(M_this_sprites_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34557),
            .ce(),
            .sr(N__28665));
    defparam M_this_sprites_address_q_11_LC_20_12_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_11_LC_20_12_6.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_11_LC_20_12_6.LUT_INIT=16'b0000100000001010;
    LogicCell40 M_this_sprites_address_q_11_LC_20_12_6 (
            .in0(N__22854),
            .in1(N__24141),
            .in2(N__22863),
            .in3(N__29008),
            .lcout(M_this_sprites_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34557),
            .ce(),
            .sr(N__28665));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_11_LC_20_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_11_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_11_LC_20_13_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_11_LC_20_13_1  (
            .in0(N__27552),
            .in1(N__33608),
            .in2(N__29021),
            .in3(N__27681),
            .lcout(N_792),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_11_LC_20_13_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_11_LC_20_13_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_11_LC_20_13_2.LUT_INIT=16'b0000000011011101;
    LogicCell40 M_this_sprites_address_q_RNO_0_11_LC_20_13_2 (
            .in0(N__26298),
            .in1(N__30279),
            .in2(_gnd_net_),
            .in3(N__29091),
            .lcout(M_this_sprites_address_qc_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_10_LC_20_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_10_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_10_LC_20_13_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_10_LC_20_13_4  (
            .in0(N__27680),
            .in1(N__29003),
            .in2(N__33753),
            .in3(N__27553),
            .lcout(N_795),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_13_LC_20_14_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_13_LC_20_14_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_13_LC_20_14_2.LUT_INIT=16'b0000001100000001;
    LogicCell40 M_this_sprites_address_q_RNO_0_13_LC_20_14_2 (
            .in0(N__26310),
            .in1(N__29114),
            .in2(N__23157),
            .in3(N__30084),
            .lcout(M_this_sprites_address_qc_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_LC_20_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_LC_20_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_LC_20_14_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_LC_20_14_5  (
            .in0(_gnd_net_),
            .in1(N__27504),
            .in2(_gnd_net_),
            .in3(N__35087),
            .lcout(N_773_0),
            .ltout(N_773_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_9_LC_20_14_6.C_ON=1'b0;
    defparam M_this_state_q_9_LC_20_14_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_9_LC_20_14_6.LUT_INIT=16'b1111000000000000;
    LogicCell40 M_this_state_q_9_LC_20_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22827),
            .in3(N__22930),
            .lcout(M_this_state_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34571),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_443_i_LC_20_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.N_443_i_LC_20_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_443_i_LC_20_14_7 .LUT_INIT=16'b1111011111110011;
    LogicCell40 \this_vga_signals.N_443_i_LC_20_14_7  (
            .in0(N__22824),
            .in1(N__28947),
            .in2(N__24489),
            .in3(N__27503),
            .lcout(N_443_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_0_LC_20_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_0_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_0_LC_20_15_0 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_0_LC_20_15_0  (
            .in0(N__27297),
            .in1(N__34193),
            .in2(N__33609),
            .in3(N__27328),
            .lcout(N_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_13_LC_20_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_13_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_13_LC_20_15_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_13_LC_20_15_3  (
            .in0(N__28993),
            .in1(N__27668),
            .in2(N__35425),
            .in3(N__27505),
            .lcout(N_126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_en_0_i_0_0_LC_20_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_en_0_i_0_0_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_en_0_i_0_0_LC_20_15_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_en_0_i_0_0_LC_20_15_4  (
            .in0(N__27296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24483),
            .lcout(N_23_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIUK1S_3_LC_20_15_5.C_ON=1'b0;
    defparam M_this_state_q_RNIUK1S_3_LC_20_15_5.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIUK1S_3_LC_20_15_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_state_q_RNIUK1S_3_LC_20_15_5 (
            .in0(N__23217),
            .in1(N__22993),
            .in2(N__24437),
            .in3(N__23608),
            .lcout(),
            .ltout(port_dmab_ac0_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI392H1_1_LC_20_15_6.C_ON=1'b0;
    defparam M_this_state_q_RNI392H1_1_LC_20_15_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI392H1_1_LC_20_15_6.LUT_INIT=16'b0000000000010000;
    LogicCell40 M_this_state_q_RNI392H1_1_LC_20_15_6 (
            .in0(N__24490),
            .in1(N__23137),
            .in2(N__23109),
            .in3(N__22893),
            .lcout(port_dmab_ac0_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_2_LC_20_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_2_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_2_LC_20_15_7 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_2_LC_20_15_7  (
            .in0(N__27329),
            .in1(N__35410),
            .in2(N__33908),
            .in3(N__27298),
            .lcout(N_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_2_13_LC_20_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_2_13_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_2_13_LC_20_16_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_a2_2_13_LC_20_16_0  (
            .in0(N__27418),
            .in1(N__25247),
            .in2(_gnd_net_),
            .in3(N__28941),
            .lcout(N_809),
            .ltout(N_809_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_8_LC_20_16_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_8_LC_20_16_1.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_8_LC_20_16_1.LUT_INIT=16'b0000101000001111;
    LogicCell40 M_this_sprites_address_q_RNO_0_8_LC_20_16_1 (
            .in0(N__24525),
            .in1(_gnd_net_),
            .in2(N__22998),
            .in3(N__26285),
            .lcout(M_this_sprites_address_qc_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_394_0_i_i_o2_LC_20_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.N_394_0_i_i_o2_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_394_0_i_i_o2_LC_20_16_3 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \this_vga_signals.N_394_0_i_i_o2_LC_20_16_3  (
            .in0(N__22995),
            .in1(N__25246),
            .in2(N__23346),
            .in3(N__27417),
            .lcout(N_749_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2_0_a3_0_a2_0_a2_LC_20_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2_0_a3_0_a2_0_a2_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2_0_a3_0_a2_0_a2_LC_20_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2_0_a3_0_a2_0_a2_LC_20_16_5  (
            .in0(_gnd_net_),
            .in1(N__22937),
            .in2(_gnd_net_),
            .in3(N__27416),
            .lcout(\this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_4_13_LC_20_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_4_13_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_4_13_LC_20_16_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_a2_4_13_LC_20_16_7  (
            .in0(N__27625),
            .in1(N__22892),
            .in2(_gnd_net_),
            .in3(N__27419),
            .lcout(N_813),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.M_this_start_address_delay_out_i_0_i2_i_o2_0_LC_20_17_1 .C_ON=1'b0;
    defparam \this_start_address_delay.M_this_start_address_delay_out_i_0_i2_i_o2_0_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \this_start_address_delay.M_this_start_address_delay_out_i_0_i2_i_o2_0_LC_20_17_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_start_address_delay.M_this_start_address_delay_out_i_0_i2_i_o2_0_LC_20_17_1  (
            .in0(N__23283),
            .in1(N__23245),
            .in2(_gnd_net_),
            .in3(N__23581),
            .lcout(N_775_0),
            .ltout(N_775_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_1_0_LC_20_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_1_0_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_1_0_LC_20_17_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_1_0_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23382),
            .in3(N__23379),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_o2_LC_20_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_o2_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_o2_LC_20_17_3 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_o2_LC_20_17_3  (
            .in0(N__23643),
            .in1(N__23246),
            .in2(N__23289),
            .in3(N__23582),
            .lcout(N_122_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_o2_LC_20_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_o2_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_o2_LC_20_17_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_o2_LC_20_17_5  (
            .in0(N__23285),
            .in1(N__23244),
            .in2(_gnd_net_),
            .in3(N__23580),
            .lcout(N_87_0),
            .ltout(N_87_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a3_0_a2_0_LC_20_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a3_0_a2_0_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a3_0_a2_0_LC_20_17_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a3_0_a2_0_LC_20_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23349),
            .in3(N__23342),
            .lcout(N_163),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_20_17_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_20_17_7 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_20_17_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_20_17_7  (
            .in0(N__23284),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23583),
            .lcout(this_start_data_delay_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34591),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_5_LC_20_18_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_5_LC_20_18_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_5_LC_20_18_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_5_LC_20_18_1  (
            .in0(_gnd_net_),
            .in1(N__34831),
            .in2(_gnd_net_),
            .in3(N__23229),
            .lcout(\this_reset_cond.M_stage_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34597),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_9_0_i_LC_20_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_9_0_i_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_9_0_i_LC_20_18_2 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_9_0_i_LC_20_18_2  (
            .in0(N__23223),
            .in1(N__24495),
            .in2(N__23638),
            .in3(N__27457),
            .lcout(un1_M_this_state_q_9_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_20_18_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_20_18_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_20_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_20_18_5  (
            .in0(N__23166),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34597),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_19_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_19_0  (
            .in0(_gnd_net_),
            .in1(N__23568),
            .in2(N__30779),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_19_0_),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_19_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_19_1  (
            .in0(_gnd_net_),
            .in1(N__23553),
            .in2(N__31895),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_0 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_19_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_19_2  (
            .in0(_gnd_net_),
            .in1(N__23538),
            .in2(N__30590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_1 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_19_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_19_3  (
            .in0(_gnd_net_),
            .in1(N__32965),
            .in2(N__23523),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_2 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_19_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_19_4  (
            .in0(_gnd_net_),
            .in1(N__33042),
            .in2(N__23505),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_3 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_19_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_19_5  (
            .in0(_gnd_net_),
            .in1(N__33075),
            .in2(N__23487),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_4 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_19_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_19_6  (
            .in0(_gnd_net_),
            .in1(N__32997),
            .in2(N__23469),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_5 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_19_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_19_7  (
            .in0(_gnd_net_),
            .in1(N__23450),
            .in2(N__32124),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_6 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_20_20_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_20_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_20_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23736),
            .lcout(\this_ppu.un1_M_vaddress_q_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_11_LC_20_20_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_11_LC_20_20_2 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_11_LC_20_20_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \this_sprites_ram.mem_radreg_11_LC_20_20_2  (
            .in0(N__31672),
            .in1(N__31477),
            .in2(N__23724),
            .in3(N__32232),
            .lcout(\this_sprites_ram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34606),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIMU531_13_LC_20_20_4.C_ON=1'b0;
    defparam M_this_state_q_RNIMU531_13_LC_20_20_4.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIMU531_13_LC_20_20_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_state_q_RNIMU531_13_LC_20_20_4 (
            .in0(N__32769),
            .in1(N__23639),
            .in2(N__32691),
            .in3(N__27527),
            .lcout(un1_M_this_oam_address_q_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_1_LC_20_20_5.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_1_LC_20_20_5.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_1_LC_20_20_5.LUT_INIT=16'b1111111100100000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_1_LC_20_20_5 (
            .in0(N__32665),
            .in1(N__32774),
            .in2(N__32384),
            .in3(N__35074),
            .lcout(N_1174_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_20_20_6.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_20_20_6.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_20_20_6.LUT_INIT=16'b1010101010101110;
    LogicCell40 M_this_oam_address_q_RNI24IA1_1_1_LC_20_20_6 (
            .in0(N__35072),
            .in1(N__32336),
            .in2(N__32844),
            .in3(N__32664),
            .lcout(N_1190_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_20_20_7.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_20_20_7.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_20_20_7.LUT_INIT=16'b1111111100001000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_0_1_LC_20_20_7 (
            .in0(N__32335),
            .in1(N__32773),
            .in2(N__32692),
            .in3(N__35073),
            .lcout(N_1182_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNILNG41_3_LC_20_21_0.C_ON=1'b0;
    defparam M_this_oam_address_q_RNILNG41_3_LC_20_21_0.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNILNG41_3_LC_20_21_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 M_this_oam_address_q_RNILNG41_3_LC_20_21_0 (
            .in0(N__24772),
            .in1(N__26411),
            .in2(_gnd_net_),
            .in3(N__26437),
            .lcout(un1_M_this_oam_address_q_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_23_LC_20_25_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_23_LC_20_25_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_23_LC_20_25_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_23_LC_20_25_1 (
            .in0(N__35222),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34623),
            .ce(N__28325),
            .sr(N__34995));
    defparam M_this_data_tmp_q_esr_18_LC_20_25_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_18_LC_20_25_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_18_LC_20_25_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_18_LC_20_25_6 (
            .in0(N__33844),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34623),
            .ce(N__28325),
            .sr(N__34995));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_10_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_10_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_10_6  (
            .in0(N__29651),
            .in1(N__24126),
            .in2(_gnd_net_),
            .in3(N__24111),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_21_11_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_21_11_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_21_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_21_11_2  (
            .in0(N__24093),
            .in1(N__24081),
            .in2(_gnd_net_),
            .in3(N__29656),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_11_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_11_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_11_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_11_5  (
            .in0(N__29657),
            .in1(_gnd_net_),
            .in2(N__24063),
            .in3(N__24048),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_10_LC_21_12_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_10_LC_21_12_1.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_10_LC_21_12_1.LUT_INIT=16'b0000000010111011;
    LogicCell40 M_this_sprites_address_q_RNO_0_10_LC_21_12_1 (
            .in0(N__24181),
            .in1(N__26308),
            .in2(_gnd_net_),
            .in3(N__29112),
            .lcout(M_this_sprites_address_qc_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_21_12_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_21_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_wclke_3_LC_21_12_2  (
            .in0(N__30219),
            .in1(N__30280),
            .in2(N__30123),
            .in3(N__30053),
            .lcout(\this_sprites_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_0_LC_21_13_0.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_0_0_LC_21_13_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_0_LC_21_13_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_0_0_LC_21_13_0 (
            .in0(_gnd_net_),
            .in1(N__23824),
            .in2(N__23775),
            .in3(N__23774),
            .lcout(M_this_sprites_address_q_RNO_0Z0Z_0),
            .ltout(),
            .carryin(bfn_21_13_0_),
            .carryout(un1_M_this_sprites_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_21_13_1.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_21_13_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_21_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_21_13_1 (
            .in0(_gnd_net_),
            .in1(N__27740),
            .in2(_gnd_net_),
            .in3(N__23745),
            .lcout(un1_M_this_sprites_address_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_0),
            .carryout(un1_M_this_sprites_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_2_LC_21_13_2.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_0_2_LC_21_13_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_2_LC_21_13_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_0_2_LC_21_13_2 (
            .in0(_gnd_net_),
            .in1(N__25410),
            .in2(_gnd_net_),
            .in3(N__23742),
            .lcout(M_this_sprites_address_q_RNO_0Z0Z_2),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_1),
            .carryout(un1_M_this_sprites_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_3_LC_21_13_3.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_0_3_LC_21_13_3.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_3_LC_21_13_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_0_3_LC_21_13_3 (
            .in0(_gnd_net_),
            .in1(N__25828),
            .in2(_gnd_net_),
            .in3(N__23739),
            .lcout(M_this_sprites_address_q_RNO_0Z0Z_3),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_2),
            .carryout(un1_M_this_sprites_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_4_LC_21_13_4.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_0_4_LC_21_13_4.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_4_LC_21_13_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_0_4_LC_21_13_4 (
            .in0(_gnd_net_),
            .in1(N__26654),
            .in2(_gnd_net_),
            .in3(N__24384),
            .lcout(M_this_sprites_address_q_RNO_0Z0Z_4),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_3),
            .carryout(un1_M_this_sprites_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_5_LC_21_13_5.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_0_5_LC_21_13_5.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_5_LC_21_13_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_0_5_LC_21_13_5 (
            .in0(_gnd_net_),
            .in1(N__28764),
            .in2(_gnd_net_),
            .in3(N__24381),
            .lcout(M_this_sprites_address_q_RNO_0Z0Z_5),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_4),
            .carryout(un1_M_this_sprites_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_6_LC_21_13_6.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_0_6_LC_21_13_6.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_6_LC_21_13_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_0_6_LC_21_13_6 (
            .in0(_gnd_net_),
            .in1(N__27928),
            .in2(_gnd_net_),
            .in3(N__24378),
            .lcout(M_this_sprites_address_q_RNO_0Z0Z_6),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_5),
            .carryout(un1_M_this_sprites_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_7_LC_21_13_7.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_7_LC_21_13_7.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_7_LC_21_13_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_7_LC_21_13_7 (
            .in0(_gnd_net_),
            .in1(N__25018),
            .in2(_gnd_net_),
            .in3(N__24375),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_7),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_6),
            .carryout(un1_M_this_sprites_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_8_LC_21_14_0.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_8_LC_21_14_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_8_LC_21_14_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_8_LC_21_14_0 (
            .in0(_gnd_net_),
            .in1(N__24524),
            .in2(_gnd_net_),
            .in3(N__24372),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_8),
            .ltout(),
            .carryin(bfn_21_14_0_),
            .carryout(un1_M_this_sprites_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_9_LC_21_14_1.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_9_LC_21_14_1.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_9_LC_21_14_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_9_LC_21_14_1 (
            .in0(_gnd_net_),
            .in1(N__26050),
            .in2(_gnd_net_),
            .in3(N__24369),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_9),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_8),
            .carryout(un1_M_this_sprites_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_10_LC_21_14_2.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_10_LC_21_14_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_10_LC_21_14_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_10_LC_21_14_2 (
            .in0(_gnd_net_),
            .in1(N__24194),
            .in2(_gnd_net_),
            .in3(N__24144),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_10),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_9),
            .carryout(un1_M_this_sprites_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_11_LC_21_14_3.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_11_LC_21_14_3.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_11_LC_21_14_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_11_LC_21_14_3 (
            .in0(_gnd_net_),
            .in1(N__30293),
            .in2(_gnd_net_),
            .in3(N__24132),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_11),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_10),
            .carryout(un1_M_this_sprites_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_12_LC_21_14_4.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_0_12_LC_21_14_4.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_12_LC_21_14_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_0_12_LC_21_14_4 (
            .in0(_gnd_net_),
            .in1(N__30198),
            .in2(_gnd_net_),
            .in3(N__24129),
            .lcout(M_this_sprites_address_q_RNO_0Z0Z_12),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_11),
            .carryout(un1_M_this_sprites_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_13_LC_21_14_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_13_LC_21_14_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_13_LC_21_14_5.LUT_INIT=16'b0100110010001100;
    LogicCell40 M_this_sprites_address_q_13_LC_21_14_5 (
            .in0(N__30102),
            .in1(N__24753),
            .in2(N__29022),
            .in3(N__24747),
            .lcout(M_this_sprites_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34577),
            .ce(),
            .sr(N__28664));
    defparam M_this_sprites_address_q_12_LC_21_15_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_12_LC_21_15_0.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_12_LC_21_15_0.LUT_INIT=16'b0100010101000000;
    LogicCell40 M_this_sprites_address_q_12_LC_21_15_0 (
            .in0(N__29087),
            .in1(N__24744),
            .in2(N__29020),
            .in3(N__24501),
            .lcout(M_this_sprites_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34583),
            .ce(),
            .sr(N__28663));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_7_LC_21_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_7_LC_21_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_7_LC_21_15_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_7_LC_21_15_4  (
            .in0(N__27678),
            .in1(N__28994),
            .in2(N__34197),
            .in3(N__27544),
            .lcout(),
            .ltout(N_807_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_7_LC_21_15_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_7_LC_21_15_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_7_LC_21_15_5.LUT_INIT=16'b0000101000000010;
    LogicCell40 M_this_sprites_address_q_7_LC_21_15_5 (
            .in0(N__24942),
            .in1(N__28999),
            .in2(N__24738),
            .in3(N__24735),
            .lcout(M_this_sprites_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34583),
            .ce(),
            .sr(N__28663));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_8_LC_21_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_8_LC_21_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_8_LC_21_15_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_8_LC_21_15_6  (
            .in0(N__27679),
            .in1(N__34016),
            .in2(N__29019),
            .in3(N__27545),
            .lcout(),
            .ltout(N_803_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_8_LC_21_15_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_8_LC_21_15_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_8_LC_21_15_7.LUT_INIT=16'b0000110100000000;
    LogicCell40 M_this_sprites_address_q_8_LC_21_15_7 (
            .in0(N__28995),
            .in1(N__24726),
            .in2(N__24720),
            .in3(N__24717),
            .lcout(M_this_sprites_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34583),
            .ce(),
            .sr(N__28663));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_9_LC_21_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_9_LC_21_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_9_LC_21_16_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_9_LC_21_16_0  (
            .in0(N__27459),
            .in1(N__33904),
            .in2(N__27666),
            .in3(N__28942),
            .lcout(N_799),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_3_0_12_LC_21_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_3_0_12_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_3_0_12_LC_21_16_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_3_0_12_LC_21_16_3  (
            .in0(N__27632),
            .in1(N__30197),
            .in2(N__33457),
            .in3(N__27460),
            .lcout(N_602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_3_0_i_0_o2_LC_21_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_3_0_i_0_o2_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_3_0_i_0_o2_LC_21_16_5 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_3_0_i_0_o2_LC_21_16_5  (
            .in0(N__24494),
            .in1(N__24438),
            .in2(_gnd_net_),
            .in3(N__27458),
            .lcout(\this_vga_signals.un1_M_this_state_q_3_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_7_LC_21_16_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_7_LC_21_16_6.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_7_LC_21_16_6.LUT_INIT=16'b0000000010111011;
    LogicCell40 M_this_sprites_address_q_RNO_0_7_LC_21_16_6 (
            .in0(N__25001),
            .in1(N__26286),
            .in2(_gnd_net_),
            .in3(N__29071),
            .lcout(M_this_sprites_address_qc_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_17_2 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32967),
            .lcout(M_this_oam_ram_read_data_i_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_19_2 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_19_2 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30942),
            .lcout(M_this_oam_ram_read_data_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc4_LC_21_19_6 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc4_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc4_LC_21_19_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc4_LC_21_19_6  (
            .in0(N__30974),
            .in1(N__31063),
            .in2(N__24908),
            .in3(N__26505),
            .lcout(\this_ppu.un1_M_haddress_q_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_2_LC_21_20_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_2_LC_21_20_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_2_LC_21_20_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_2_LC_21_20_1 (
            .in0(N__33892),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34609),
            .ce(N__26374),
            .sr(N__34987));
    defparam M_this_data_tmp_q_esr_1_LC_21_20_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_1_LC_21_20_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_1_LC_21_20_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_1_LC_21_20_6 (
            .in0(N__34042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34609),
            .ce(N__26374),
            .sr(N__34987));
    defparam M_this_oam_address_q_0_LC_21_21_1.C_ON=1'b0;
    defparam M_this_oam_address_q_0_LC_21_21_1.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_0_LC_21_21_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_0_LC_21_21_1 (
            .in0(N__32383),
            .in1(N__26496),
            .in2(_gnd_net_),
            .in3(N__32842),
            .lcout(M_this_oam_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34612),
            .ce(),
            .sr(N__28658));
    defparam M_this_oam_address_q_5_LC_21_21_3.C_ON=1'b0;
    defparam M_this_oam_address_q_5_LC_21_21_3.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_5_LC_21_21_3.LUT_INIT=16'b0000000001111000;
    LogicCell40 M_this_oam_address_q_5_LC_21_21_3 (
            .in0(N__24860),
            .in1(N__24834),
            .in2(N__24809),
            .in3(N__26498),
            .lcout(M_this_oam_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34612),
            .ce(),
            .sr(N__28658));
    defparam M_this_oam_address_q_3_LC_21_21_4.C_ON=1'b0;
    defparam M_this_oam_address_q_3_LC_21_21_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_3_LC_21_21_4.LUT_INIT=16'b0001010001010000;
    LogicCell40 M_this_oam_address_q_3_LC_21_21_4 (
            .in0(N__26497),
            .in1(N__26407),
            .in2(N__24779),
            .in3(N__26441),
            .lcout(M_this_oam_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34612),
            .ce(),
            .sr(N__28658));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_21_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_21_22_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_21_22_2  (
            .in0(N__32376),
            .in1(N__32778),
            .in2(N__25290),
            .in3(N__32571),
            .lcout(N_746_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_5_LC_21_23_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_5_LC_21_23_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_5_LC_21_23_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 M_this_data_tmp_q_esr_5_LC_21_23_0 (
            .in0(_gnd_net_),
            .in1(N__33463),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34617),
            .ce(N__26381),
            .sr(N__34991));
    defparam M_this_data_tmp_q_esr_0_LC_21_23_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_0_LC_21_23_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_0_LC_21_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_0_LC_21_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34123),
            .lcout(M_this_data_tmp_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34617),
            .ce(N__26381),
            .sr(N__34991));
    defparam M_this_data_tmp_q_esr_4_LC_21_23_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_4_LC_21_23_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_4_LC_21_23_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_4_LC_21_23_3 (
            .in0(N__33604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34617),
            .ce(N__26381),
            .sr(N__34991));
    defparam M_this_data_tmp_q_esr_7_LC_21_23_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_7_LC_21_23_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_7_LC_21_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_7_LC_21_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35200),
            .lcout(M_this_data_tmp_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34617),
            .ce(N__26381),
            .sr(N__34991));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a2_28_LC_21_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a2_28_LC_21_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a2_28_LC_21_24_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a2_28_LC_21_24_6  (
            .in0(N__32377),
            .in1(N__32689),
            .in2(N__33606),
            .in3(N__32845),
            .lcout(M_this_oam_ram_write_data_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_21_LC_21_25_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_21_LC_21_25_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_21_LC_21_25_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_21_LC_21_25_4 (
            .in0(N__33458),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34624),
            .ce(N__28327),
            .sr(N__34993));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_4_LC_22_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_4_LC_22_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_4_LC_22_13_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_4_LC_22_13_5  (
            .in0(N__26647),
            .in1(N__27682),
            .in2(N__33607),
            .in3(N__27546),
            .lcout(N_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_3_bm_1_LC_22_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_3_bm_1_LC_22_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_3_bm_1_LC_22_13_7 .LUT_INIT=16'b0000011101110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_3_bm_1_LC_22_13_7  (
            .in0(N__25251),
            .in1(N__27547),
            .in2(N__27770),
            .in3(N__25182),
            .lcout(\this_vga_signals.M_this_sprites_address_q_3_bmZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_2_LC_22_14_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_2_LC_22_14_0.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_2_LC_22_14_0.LUT_INIT=16'b0100010001010000;
    LogicCell40 M_this_sprites_address_q_2_LC_22_14_0 (
            .in0(N__29115),
            .in1(N__26316),
            .in2(N__25380),
            .in3(N__29010),
            .lcout(M_this_sprites_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__28666));
    defparam M_this_sprites_address_q_RNO_0_9_LC_22_14_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_9_LC_22_14_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_9_LC_22_14_2.LUT_INIT=16'b0000000010111011;
    LogicCell40 M_this_sprites_address_q_RNO_0_9_LC_22_14_2 (
            .in0(N__26051),
            .in1(N__26309),
            .in2(_gnd_net_),
            .in3(N__29113),
            .lcout(),
            .ltout(M_this_sprites_address_qc_11_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_9_LC_22_14_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_9_LC_22_14_3.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_9_LC_22_14_3.LUT_INIT=16'b0011000000010000;
    LogicCell40 M_this_sprites_address_q_9_LC_22_14_3 (
            .in0(N__29009),
            .in1(N__26259),
            .in2(N__26247),
            .in3(N__26244),
            .lcout(M_this_sprites_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__28666));
    defparam M_this_sprites_address_q_3_LC_22_14_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_3_LC_22_14_6.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_3_LC_22_14_6.LUT_INIT=16'b0100010001010000;
    LogicCell40 M_this_sprites_address_q_3_LC_22_14_6 (
            .in0(N__29116),
            .in1(N__26028),
            .in2(N__25794),
            .in3(N__29011),
            .lcout(M_this_sprites_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__28666));
    defparam \this_vga_signals.M_this_sprites_address_q_3_0_i_m2_3_LC_22_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_3_0_i_m2_3_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_3_0_i_m2_3_LC_22_15_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_3_0_i_m2_3_LC_22_15_2  (
            .in0(N__25874),
            .in1(N__27677),
            .in2(N__33749),
            .in3(N__27543),
            .lcout(N_50),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIS5A21_0_LC_22_15_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIS5A21_0_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIS5A21_0_LC_22_15_3 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \this_ppu.M_vaddress_q_RNIS5A21_0_LC_22_15_3  (
            .in0(N__27186),
            .in1(N__31457),
            .in2(N__31653),
            .in3(N__30842),
            .lcout(M_this_ppu_sprites_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_2_LC_22_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_2_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_2_LC_22_15_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_2_LC_22_15_6  (
            .in0(N__25411),
            .in1(N__27676),
            .in2(N__33909),
            .in3(N__27542),
            .lcout(N_103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_1_LC_22_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_1_LC_22_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_1_LC_22_16_0 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_1_LC_22_16_0  (
            .in0(N__33416),
            .in1(N__27327),
            .in2(N__34050),
            .in3(N__27305),
            .lcout(M_this_sprites_ram_write_data_iv_i_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_15_LC_22_19_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_15_LC_22_19_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_15_LC_22_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_15_LC_22_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35168),
            .lcout(M_this_data_tmp_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34610),
            .ce(N__28217),
            .sr(N__34984));
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_5_0_LC_22_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_5_0_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_5_0_LC_22_20_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_5_0_LC_22_20_4  (
            .in0(N__26616),
            .in1(N__26598),
            .in2(N__26586),
            .in3(N__26556),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_0_a2_1_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_8_LC_22_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_8_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_8_LC_22_20_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_8_LC_22_20_5  (
            .in0(N__32375),
            .in1(N__32572),
            .in2(N__28227),
            .in3(N__32779),
            .lcout(N_54_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_ac0_1_LC_22_20_6 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_ac0_1_LC_22_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_ac0_1_LC_22_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_ac0_1_LC_22_20_6  (
            .in0(_gnd_net_),
            .in1(N__31012),
            .in2(_gnd_net_),
            .in3(N__30930),
            .lcout(\this_ppu.un1_oam_data_1_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_1_LC_22_21_0.C_ON=1'b0;
    defparam M_this_oam_address_q_1_LC_22_21_0.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_1_LC_22_21_0.LUT_INIT=16'b0001010001010000;
    LogicCell40 M_this_oam_address_q_1_LC_22_21_0 (
            .in0(N__26492),
            .in1(N__32426),
            .in2(N__32690),
            .in3(N__32843),
            .lcout(M_this_oam_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34615),
            .ce(),
            .sr(N__28661));
    defparam M_this_oam_address_q_2_LC_22_21_5.C_ON=1'b0;
    defparam M_this_oam_address_q_2_LC_22_21_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_2_LC_22_21_5.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_2_LC_22_21_5 (
            .in0(N__26406),
            .in1(N__26491),
            .in2(_gnd_net_),
            .in3(N__26445),
            .lcout(M_this_oam_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34615),
            .ce(),
            .sr(N__28661));
    defparam M_this_data_tmp_q_esr_6_LC_22_22_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_6_LC_22_22_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_6_LC_22_22_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_6_LC_22_22_0 (
            .in0(N__35427),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34618),
            .ce(N__26382),
            .sr(N__34988));
    defparam M_this_data_tmp_q_esr_3_LC_22_22_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_3_LC_22_22_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_3_LC_22_22_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_3_LC_22_22_4 (
            .in0(N__33718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34618),
            .ce(N__26382),
            .sr(N__34988));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_22_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_22_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_22_23_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_22_23_0  (
            .in0(N__32437),
            .in1(N__32853),
            .in2(N__26352),
            .in3(N__32587),
            .lcout(N_742_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_22_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_22_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_22_23_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_22_23_2  (
            .in0(N__32435),
            .in1(N__32850),
            .in2(N__33896),
            .in3(N__32582),
            .lcout(N_34_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_22_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_22_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_22_23_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_22_23_4  (
            .in0(N__32436),
            .in1(N__32851),
            .in2(N__26961),
            .in3(N__32586),
            .lcout(N_744_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_23_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_23_7  (
            .in0(N__32852),
            .in1(N__26940),
            .in2(N__32657),
            .in3(N__32438),
            .lcout(N_56_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_16_LC_22_24_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_16_LC_22_24_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_16_LC_22_24_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_16_LC_22_24_1 (
            .in0(N__34159),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34625),
            .ce(N__28328),
            .sr(N__34992));
    defparam M_this_data_tmp_q_esr_22_LC_22_24_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_22_LC_22_24_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_22_LC_22_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_22_LC_22_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35437),
            .lcout(M_this_data_tmp_qZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34625),
            .ce(N__28328),
            .sr(N__34992));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_16_LC_22_25_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_16_LC_22_25_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_16_LC_22_25_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_16_LC_22_25_0  (
            .in0(N__32453),
            .in1(N__32652),
            .in2(N__26919),
            .in3(N__32880),
            .lcout(N_738_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_22_LC_22_25_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_22_LC_22_25_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_22_LC_22_25_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_22_LC_22_25_2  (
            .in0(N__32454),
            .in1(N__32653),
            .in2(N__26898),
            .in3(N__32881),
            .lcout(N_40_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_11_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_11_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_11_7  (
            .in0(N__29652),
            .in1(N__26877),
            .in2(_gnd_net_),
            .in3(N__26862),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_4_LC_23_13_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_4_LC_23_13_0.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_4_LC_23_13_0.LUT_INIT=16'b0011001000010000;
    LogicCell40 M_this_sprites_address_q_4_LC_23_13_0 (
            .in0(N__29016),
            .in1(N__29125),
            .in2(N__26841),
            .in3(N__26832),
            .lcout(M_this_sprites_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__28667));
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_6_LC_23_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_6_LC_23_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_6_LC_23_13_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_6_LC_23_13_3  (
            .in0(N__27921),
            .in1(N__27684),
            .in2(N__35406),
            .in3(N__27548),
            .lcout(),
            .ltout(N_101_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_6_LC_23_13_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_6_LC_23_13_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_6_LC_23_13_4.LUT_INIT=16'b0011001000010000;
    LogicCell40 M_this_sprites_address_q_6_LC_23_13_4 (
            .in0(N__29017),
            .in1(N__29126),
            .in2(N__28113),
            .in3(N__28110),
            .lcout(M_this_sprites_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__28667));
    defparam M_this_sprites_address_q_1_LC_23_13_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_1_LC_23_13_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_1_LC_23_13_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 M_this_sprites_address_q_1_LC_23_13_7 (
            .in0(N__27345),
            .in1(N__29018),
            .in2(_gnd_net_),
            .in3(N__27897),
            .lcout(M_this_sprites_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__28667));
    defparam \this_vga_signals.M_this_sprites_address_q_3_0_5_LC_23_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_3_0_5_LC_23_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_3_0_5_LC_23_14_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_3_0_5_LC_23_14_3  (
            .in0(N__28701),
            .in1(N__27683),
            .in2(N__33468),
            .in3(N__27555),
            .lcout(N_595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_3_am_1_LC_23_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_3_am_1_LC_23_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_3_am_1_LC_23_15_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_3_am_1_LC_23_15_5  (
            .in0(N__27766),
            .in1(N__27669),
            .in2(N__34036),
            .in3(N__27538),
            .lcout(\this_vga_signals.M_this_sprites_address_q_3_amZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_3_LC_23_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_3_LC_23_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_3_LC_23_15_7 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_3_LC_23_15_7  (
            .in0(N__33742),
            .in1(N__27336),
            .in2(N__35211),
            .in3(N__27309),
            .lcout(M_this_sprites_ram_write_data_iv_i_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_16_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_16_0  (
            .in0(_gnd_net_),
            .in1(N__30778),
            .in2(_gnd_net_),
            .in3(N__30841),
            .lcout(\this_ppu.un2_vscroll_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_19_LC_23_18_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_19_LC_23_18_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_19_LC_23_18_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_19_LC_23_18_3 (
            .in0(N__33732),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34611),
            .ce(N__28326),
            .sr(N__34983));
    defparam \this_ppu.M_haddress_q_RNI4S061_1_LC_23_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI4S061_1_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI4S061_1_LC_23_19_2 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_haddress_q_RNI4S061_1_LC_23_19_2  (
            .in0(N__31500),
            .in1(N__29766),
            .in2(N__31683),
            .in3(N__29838),
            .lcout(M_this_ppu_sprites_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_10_LC_23_20_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_10_LC_23_20_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_10_LC_23_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_10_LC_23_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33897),
            .lcout(M_this_data_tmp_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34616),
            .ce(N__28213),
            .sr(N__34985));
    defparam M_this_data_tmp_q_esr_12_LC_23_20_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_12_LC_23_20_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_12_LC_23_20_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_12_LC_23_20_2 (
            .in0(N__33605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34616),
            .ce(N__28213),
            .sr(N__34985));
    defparam M_this_data_tmp_q_esr_13_LC_23_20_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_13_LC_23_20_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_13_LC_23_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_13_LC_23_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33447),
            .lcout(M_this_data_tmp_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34616),
            .ce(N__28213),
            .sr(N__34985));
    defparam M_this_data_tmp_q_esr_14_LC_23_20_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_14_LC_23_20_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_14_LC_23_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_14_LC_23_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35426),
            .lcout(M_this_data_tmp_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34616),
            .ce(N__28213),
            .sr(N__34985));
    defparam M_this_data_tmp_q_esr_8_LC_23_20_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_8_LC_23_20_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_8_LC_23_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_8_LC_23_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34166),
            .lcout(M_this_data_tmp_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34616),
            .ce(N__28213),
            .sr(N__34985));
    defparam M_this_data_tmp_q_esr_9_LC_23_21_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_9_LC_23_21_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_9_LC_23_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_9_LC_23_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34037),
            .lcout(M_this_data_tmp_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34619),
            .ce(N__28218),
            .sr(N__34986));
    defparam M_this_data_tmp_q_esr_11_LC_23_21_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_11_LC_23_21_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_11_LC_23_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_11_LC_23_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33731),
            .lcout(M_this_data_tmp_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34619),
            .ce(N__28218),
            .sr(N__34986));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_22_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_22_5  (
            .in0(N__32459),
            .in1(N__32574),
            .in2(N__28182),
            .in3(N__32893),
            .lcout(N_745_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_14_LC_23_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_14_LC_23_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_14_LC_23_22_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_14_LC_23_22_7  (
            .in0(N__32458),
            .in1(N__32573),
            .in2(N__28161),
            .in3(N__32892),
            .lcout(N_739_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_23_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_23_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_23_23_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_23_23_1  (
            .in0(N__32859),
            .in1(N__32441),
            .in2(N__28137),
            .in3(N__32679),
            .lcout(N_743_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_27_LC_23_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_27_LC_23_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_27_LC_23_23_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_27_LC_23_23_2  (
            .in0(N__32439),
            .in1(N__32667),
            .in2(N__33701),
            .in3(N__32860),
            .lcout(N_32_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_11_LC_23_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_11_LC_23_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_11_LC_23_23_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_11_LC_23_23_6  (
            .in0(N__32442),
            .in1(N__32668),
            .in2(N__28395),
            .in3(N__32861),
            .lcout(M_this_oam_ram_write_data_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_23_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_23_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_23_23_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_23_23_7  (
            .in0(N__32858),
            .in1(N__32440),
            .in2(N__28374),
            .in3(N__32678),
            .lcout(N_748_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_23_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_23_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_23_24_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_23_24_2  (
            .in0(N__32666),
            .in1(N__32443),
            .in2(N__28338),
            .in3(N__32862),
            .lcout(N_44_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_17_LC_23_24_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_17_LC_23_24_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_17_LC_23_24_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_17_LC_23_24_3 (
            .in0(N__34020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34628),
            .ce(N__28329),
            .sr(N__34989));
    defparam M_this_data_tmp_q_esr_20_LC_23_24_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_20_LC_23_24_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_20_LC_23_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_20_LC_23_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33585),
            .lcout(M_this_data_tmp_qZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34628),
            .ce(N__28329),
            .sr(N__34989));
    defparam \this_vga_signals.M_this_oam_ram_write_data_23_LC_23_25_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_23_LC_23_25_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_23_LC_23_25_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_23_LC_23_25_2  (
            .in0(N__32863),
            .in1(N__28269),
            .in2(N__32693),
            .in3(N__32456),
            .lcout(M_this_oam_ram_write_data_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_23_25_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_23_25_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_23_25_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_23_25_3  (
            .in0(N__32455),
            .in1(N__32669),
            .in2(N__28248),
            .in3(N__32864),
            .lcout(N_42_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a2_30_LC_23_25_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a2_30_LC_23_25_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a2_30_LC_23_25_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a2_30_LC_23_25_6  (
            .in0(N__32865),
            .in1(N__35438),
            .in2(N__32694),
            .in3(N__32457),
            .lcout(M_this_oam_ram_write_data_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_24_10_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_24_10_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_24_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_24_10_0  (
            .in0(N__29676),
            .in1(N__29670),
            .in2(_gnd_net_),
            .in3(N__29658),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI70261_2_LC_24_11_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI70261_2_LC_24_11_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI70261_2_LC_24_11_3 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_haddress_q_RNI70261_2_LC_24_11_3  (
            .in0(N__31502),
            .in1(N__31803),
            .in2(N__31678),
            .in3(N__29741),
            .lcout(M_this_ppu_sprites_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_12_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_12_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_12_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_12_3  (
            .in0(N__30241),
            .in1(N__30295),
            .in2(N__30158),
            .in3(N__30051),
            .lcout(\this_sprites_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_13_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_13_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_13_3  (
            .in0(N__30319),
            .in1(N__30240),
            .in2(N__30144),
            .in3(N__30050),
            .lcout(\this_sprites_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_24_13_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_24_13_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_24_13_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_24_13_6  (
            .in0(N__31464),
            .in1(N__30552),
            .in2(N__31652),
            .in3(N__30642),
            .lcout(M_this_ppu_sprites_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_5_LC_24_14_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_5_LC_24_14_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_5_LC_24_14_5.LUT_INIT=16'b0100010001010000;
    LogicCell40 M_this_sprites_address_q_5_LC_24_14_5 (
            .in0(N__29127),
            .in1(N__29043),
            .in2(N__29031),
            .in3(N__29012),
            .lcout(M_this_sprites_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34598),
            .ce(),
            .sr(N__28668));
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_15_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_15_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_15_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_15_3  (
            .in0(N__30320),
            .in1(N__30220),
            .in2(N__30159),
            .in3(N__30049),
            .lcout(\this_sprites_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_24_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_24_15_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_24_15_6  (
            .in0(N__31499),
            .in1(N__30651),
            .in2(N__31677),
            .in3(N__30699),
            .lcout(M_this_ppu_sprites_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_vscroll_cry_0_c_inv_LC_24_16_0 .C_ON=1'b1;
    defparam \this_ppu.un2_vscroll_cry_0_c_inv_LC_24_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_vscroll_cry_0_c_inv_LC_24_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un2_vscroll_cry_0_c_inv_LC_24_16_0  (
            .in0(_gnd_net_),
            .in1(N__30840),
            .in2(N__30708),
            .in3(N__30765),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_16 ),
            .ltout(),
            .carryin(bfn_24_16_0_),
            .carryout(\this_ppu.un2_vscroll_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_24_16_1 .C_ON=1'b1;
    defparam \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_24_16_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_24_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_24_16_1  (
            .in0(_gnd_net_),
            .in1(N__30690),
            .in2(N__31848),
            .in3(N__30645),
            .lcout(\this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0 ),
            .ltout(),
            .carryin(\this_ppu.un2_vscroll_cry_0 ),
            .carryout(\this_ppu.un2_vscroll_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_24_16_2 .C_ON=1'b0;
    defparam \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_24_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_24_16_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_24_16_2  (
            .in0(N__30635),
            .in1(N__30589),
            .in2(_gnd_net_),
            .in3(N__30555),
            .lcout(\this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI53UU_6_LC_24_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI53UU_6_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI53UU_6_LC_24_17_1 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \this_ppu.M_state_q_RNI53UU_6_LC_24_17_1  (
            .in0(N__30543),
            .in1(N__31482),
            .in2(N__31673),
            .in3(N__32178),
            .lcout(M_this_ppu_sprites_addr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_17_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_17_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_17_3  (
            .in0(N__30324),
            .in1(N__30242),
            .in2(N__30160),
            .in3(N__30052),
            .lcout(\this_sprites_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_19_0 .C_ON=1'b1;
    defparam \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_19_0  (
            .in0(_gnd_net_),
            .in1(N__29973),
            .in2(N__29847),
            .in3(N__29895),
            .lcout(\this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ),
            .ltout(),
            .carryin(bfn_24_19_0_),
            .carryout(\this_ppu.un2_hscroll_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_19_1 .C_ON=1'b1;
    defparam \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_19_1  (
            .in0(_gnd_net_),
            .in1(N__29837),
            .in2(N__31755),
            .in3(N__29760),
            .lcout(\this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0 ),
            .ltout(),
            .carryin(\this_ppu.un2_hscroll_cry_0 ),
            .carryout(\this_ppu.un2_hscroll_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_19_2 .C_ON=1'b0;
    defparam \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_19_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_19_2  (
            .in0(N__29753),
            .in1(N__31825),
            .in2(_gnd_net_),
            .in3(N__31806),
            .lcout(\this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_19_3 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31789),
            .lcout(M_this_oam_ram_read_data_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_24_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_24_20_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_24_20_2  (
            .in0(N__32373),
            .in1(N__32687),
            .in2(N__31746),
            .in3(N__32854),
            .lcout(N_747_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_10_LC_24_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_10_LC_24_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_10_LC_24_20_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_10_LC_24_20_6  (
            .in0(N__32374),
            .in1(N__32688),
            .in2(N__31722),
            .in3(N__32855),
            .lcout(M_this_oam_ram_write_data_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI43UU_6_LC_24_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI43UU_6_LC_24_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI43UU_6_LC_24_21_4 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \this_ppu.M_state_q_RNI43UU_6_LC_24_21_4  (
            .in0(N__31959),
            .in1(N__31704),
            .in2(N__31682),
            .in3(N__31437),
            .lcout(M_this_ppu_sprites_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_24_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_24_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_24_22_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_24_22_0  (
            .in0(N__32857),
            .in1(N__32432),
            .in2(N__31089),
            .in3(N__32677),
            .lcout(N_740_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc3_LC_24_22_2 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc3_LC_24_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc3_LC_24_22_2 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc3_LC_24_22_2  (
            .in0(N__31050),
            .in1(N__31002),
            .in2(N__30970),
            .in3(N__30918),
            .lcout(\this_ppu.un1_M_haddress_q_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_19_LC_24_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_19_LC_24_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_19_LC_24_22_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_19_LC_24_22_4  (
            .in0(N__32856),
            .in1(N__32431),
            .in2(N__30882),
            .in3(N__32676),
            .lcout(M_this_oam_ram_write_data_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un9lto7_4_LC_24_22_6 .C_ON=1'b0;
    defparam \this_ppu.un9lto7_4_LC_24_22_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un9lto7_4_LC_24_22_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un9lto7_4_LC_24_22_6  (
            .in0(N__32255),
            .in1(N__32225),
            .in2(N__32201),
            .in3(N__32174),
            .lcout(\this_ppu.un9lto7Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_24_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_24_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_24_23_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_24_23_0  (
            .in0(N__32429),
            .in1(N__32656),
            .in2(N__32142),
            .in3(N__32849),
            .lcout(N_741_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_ac0_1_LC_24_23_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_ac0_1_LC_24_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_ac0_1_LC_24_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.un1_oam_data_ac0_1_LC_24_23_1  (
            .in0(_gnd_net_),
            .in1(N__33030),
            .in2(_gnd_net_),
            .in3(N__32943),
            .lcout(),
            .ltout(\this_ppu.un1_oam_data_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc4_LC_24_23_2 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc4_LC_24_23_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc4_LC_24_23_2 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.un1_oam_data_axbxc4_LC_24_23_2  (
            .in0(N__33071),
            .in1(N__32111),
            .in2(N__32097),
            .in3(N__32996),
            .lcout(\this_ppu.un1_M_vaddress_q_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_13_LC_24_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_13_LC_24_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_13_LC_24_23_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_13_LC_24_23_3  (
            .in0(N__32847),
            .in1(N__32430),
            .in2(N__32079),
            .in3(N__32686),
            .lcout(M_this_oam_ram_write_data_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_15_LC_24_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_15_LC_24_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_15_LC_24_23_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_15_LC_24_23_4  (
            .in0(N__32428),
            .in1(N__32655),
            .in2(N__32061),
            .in3(N__32848),
            .lcout(M_this_oam_ram_write_data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o2_LC_24_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o2_LC_24_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o2_LC_24_23_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o2_LC_24_23_6  (
            .in0(N__32427),
            .in1(N__32654),
            .in2(_gnd_net_),
            .in3(N__32846),
            .lcout(N_123_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un9lto7_5_LC_24_23_7 .C_ON=1'b0;
    defparam \this_ppu.un9lto7_5_LC_24_23_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un9lto7_5_LC_24_23_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un9lto7_5_LC_24_23_7  (
            .in0(N__32009),
            .in1(N__31973),
            .in2(N__31958),
            .in3(N__31925),
            .lcout(\this_ppu.un9lto7Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_24_0 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_24_0 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_24_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_24_0  (
            .in0(N__31873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_oam_ram_read_data_i_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_18_LC_24_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_18_LC_24_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_18_LC_24_24_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_18_LC_24_24_3  (
            .in0(N__32433),
            .in1(N__32680),
            .in2(N__33147),
            .in3(N__32876),
            .lcout(M_this_oam_ram_write_data_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc2_LC_24_24_4 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc2_LC_24_24_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc2_LC_24_24_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.un1_oam_data_axbxc2_LC_24_24_4  (
            .in0(N__33067),
            .in1(N__33034),
            .in2(_gnd_net_),
            .in3(N__32949),
            .lcout(\this_ppu.un1_M_vaddress_q_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_24_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_24_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_24_24_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_24_24_5  (
            .in0(N__32434),
            .in1(N__32681),
            .in2(N__34191),
            .in3(N__32877),
            .lcout(N_38_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a2_31_LC_24_25_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a2_31_LC_24_25_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a2_31_LC_24_25_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a2_31_LC_24_25_0  (
            .in0(N__32460),
            .in1(N__32682),
            .in2(N__35221),
            .in3(N__32878),
            .lcout(M_this_oam_ram_write_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_24_25_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_24_25_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_24_25_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_24_25_1  (
            .in0(N__32895),
            .in1(N__32685),
            .in2(N__33467),
            .in3(N__32463),
            .lcout(N_736_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_24_25_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_24_25_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_24_25_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_24_25_2  (
            .in0(N__32461),
            .in1(N__32683),
            .in2(N__34041),
            .in3(N__32879),
            .lcout(N_737_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc3_LC_24_25_4 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc3_LC_24_25_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc3_LC_24_25_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.un1_oam_data_axbxc3_LC_24_25_4  (
            .in0(N__33066),
            .in1(N__33029),
            .in2(N__32995),
            .in3(N__32942),
            .lcout(\this_ppu.un1_M_vaddress_q_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_21_LC_24_25_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_21_LC_24_25_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_21_LC_24_25_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_21_LC_24_25_7  (
            .in0(N__32894),
            .in1(N__32684),
            .in2(N__32475),
            .in3(N__32462),
            .lcout(M_this_oam_ram_write_data_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_8_LC_26_18_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_8_LC_26_18_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_8_LC_26_18_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_8_LC_26_18_2  (
            .in0(_gnd_net_),
            .in1(N__34850),
            .in2(_gnd_net_),
            .in3(N__33312),
            .lcout(\this_reset_cond.M_stage_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34622),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_6_LC_26_18_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_6_LC_26_18_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_6_LC_26_18_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_6_LC_26_18_3  (
            .in0(N__34848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33327),
            .lcout(\this_reset_cond.M_stage_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34622),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_7_LC_26_18_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_7_LC_26_18_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_7_LC_26_18_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_7_LC_26_18_7  (
            .in0(N__34849),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33318),
            .lcout(\this_reset_cond.M_stage_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34622),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_0_LC_28_21_0.C_ON=1'b1;
    defparam M_this_external_address_q_0_LC_28_21_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_0_LC_28_21_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_0_LC_28_21_0 (
            .in0(N__35302),
            .in1(N__33269),
            .in2(N__33306),
            .in3(N__33305),
            .lcout(M_this_external_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_28_21_0_),
            .carryout(un1_M_this_external_address_q_cry_0),
            .clk(N__34631),
            .ce(),
            .sr(N__34981));
    defparam M_this_external_address_q_1_LC_28_21_1.C_ON=1'b1;
    defparam M_this_external_address_q_1_LC_28_21_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_1_LC_28_21_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_1_LC_28_21_1 (
            .in0(N__35311),
            .in1(N__33245),
            .in2(_gnd_net_),
            .in3(N__33234),
            .lcout(M_this_external_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_0),
            .carryout(un1_M_this_external_address_q_cry_1),
            .clk(N__34631),
            .ce(),
            .sr(N__34981));
    defparam M_this_external_address_q_2_LC_28_21_2.C_ON=1'b1;
    defparam M_this_external_address_q_2_LC_28_21_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_2_LC_28_21_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_2_LC_28_21_2 (
            .in0(N__35303),
            .in1(N__33224),
            .in2(_gnd_net_),
            .in3(N__33213),
            .lcout(M_this_external_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_1),
            .carryout(un1_M_this_external_address_q_cry_2),
            .clk(N__34631),
            .ce(),
            .sr(N__34981));
    defparam M_this_external_address_q_3_LC_28_21_3.C_ON=1'b1;
    defparam M_this_external_address_q_3_LC_28_21_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_3_LC_28_21_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_3_LC_28_21_3 (
            .in0(N__35312),
            .in1(N__33200),
            .in2(_gnd_net_),
            .in3(N__33189),
            .lcout(M_this_external_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_2),
            .carryout(un1_M_this_external_address_q_cry_3),
            .clk(N__34631),
            .ce(),
            .sr(N__34981));
    defparam M_this_external_address_q_4_LC_28_21_4.C_ON=1'b1;
    defparam M_this_external_address_q_4_LC_28_21_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_4_LC_28_21_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_4_LC_28_21_4 (
            .in0(N__35304),
            .in1(N__33179),
            .in2(_gnd_net_),
            .in3(N__33168),
            .lcout(M_this_external_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_3),
            .carryout(un1_M_this_external_address_q_cry_4),
            .clk(N__34631),
            .ce(),
            .sr(N__34981));
    defparam M_this_external_address_q_5_LC_28_21_5.C_ON=1'b1;
    defparam M_this_external_address_q_5_LC_28_21_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_5_LC_28_21_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_5_LC_28_21_5 (
            .in0(N__35313),
            .in1(N__33161),
            .in2(_gnd_net_),
            .in3(N__33150),
            .lcout(M_this_external_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_4),
            .carryout(un1_M_this_external_address_q_cry_5),
            .clk(N__34631),
            .ce(),
            .sr(N__34981));
    defparam M_this_external_address_q_6_LC_28_21_6.C_ON=1'b1;
    defparam M_this_external_address_q_6_LC_28_21_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_6_LC_28_21_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_6_LC_28_21_6 (
            .in0(N__35305),
            .in1(N__34241),
            .in2(_gnd_net_),
            .in3(N__34230),
            .lcout(M_this_external_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_5),
            .carryout(un1_M_this_external_address_q_cry_6),
            .clk(N__34631),
            .ce(),
            .sr(N__34981));
    defparam M_this_external_address_q_7_LC_28_21_7.C_ON=1'b1;
    defparam M_this_external_address_q_7_LC_28_21_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_7_LC_28_21_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_7_LC_28_21_7 (
            .in0(N__35310),
            .in1(N__34211),
            .in2(_gnd_net_),
            .in3(N__34200),
            .lcout(M_this_external_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_6),
            .carryout(un1_M_this_external_address_q_cry_7),
            .clk(N__34631),
            .ce(),
            .sr(N__34981));
    defparam M_this_external_address_q_8_LC_28_22_0.C_ON=1'b1;
    defparam M_this_external_address_q_8_LC_28_22_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_8_LC_28_22_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_external_address_q_8_LC_28_22_0 (
            .in0(N__34192),
            .in1(N__35298),
            .in2(N__34070),
            .in3(N__34053),
            .lcout(M_this_external_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_28_22_0_),
            .carryout(un1_M_this_external_address_q_cry_8),
            .clk(N__34637),
            .ce(),
            .sr(N__34982));
    defparam M_this_external_address_q_9_LC_28_22_1.C_ON=1'b1;
    defparam M_this_external_address_q_9_LC_28_22_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_9_LC_28_22_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_external_address_q_9_LC_28_22_1 (
            .in0(N__34046),
            .in1(N__35306),
            .in2(N__33929),
            .in3(N__33912),
            .lcout(M_this_external_address_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_8),
            .carryout(un1_M_this_external_address_q_cry_9),
            .clk(N__34637),
            .ce(),
            .sr(N__34982));
    defparam M_this_external_address_q_10_LC_28_22_2.C_ON=1'b1;
    defparam M_this_external_address_q_10_LC_28_22_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_10_LC_28_22_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_external_address_q_10_LC_28_22_2 (
            .in0(N__33879),
            .in1(N__35299),
            .in2(N__33773),
            .in3(N__33756),
            .lcout(M_this_external_address_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_9),
            .carryout(un1_M_this_external_address_q_cry_10),
            .clk(N__34637),
            .ce(),
            .sr(N__34982));
    defparam M_this_external_address_q_11_LC_28_22_3.C_ON=1'b1;
    defparam M_this_external_address_q_11_LC_28_22_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_11_LC_28_22_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_external_address_q_11_LC_28_22_3 (
            .in0(N__33697),
            .in1(N__35307),
            .in2(N__33629),
            .in3(N__33612),
            .lcout(M_this_external_address_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_10),
            .carryout(un1_M_this_external_address_q_cry_11),
            .clk(N__34637),
            .ce(),
            .sr(N__34982));
    defparam M_this_external_address_q_12_LC_28_22_4.C_ON=1'b1;
    defparam M_this_external_address_q_12_LC_28_22_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_12_LC_28_22_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_external_address_q_12_LC_28_22_4 (
            .in0(N__33584),
            .in1(N__35300),
            .in2(N__33488),
            .in3(N__33471),
            .lcout(M_this_external_address_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_11),
            .carryout(un1_M_this_external_address_q_cry_12),
            .clk(N__34637),
            .ce(),
            .sr(N__34982));
    defparam M_this_external_address_q_13_LC_28_22_5.C_ON=1'b1;
    defparam M_this_external_address_q_13_LC_28_22_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_13_LC_28_22_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_external_address_q_13_LC_28_22_5 (
            .in0(N__33405),
            .in1(N__35308),
            .in2(N__33344),
            .in3(N__35442),
            .lcout(M_this_external_address_qZ0Z_13),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_12),
            .carryout(un1_M_this_external_address_q_cry_13),
            .clk(N__34637),
            .ce(),
            .sr(N__34982));
    defparam M_this_external_address_q_14_LC_28_22_6.C_ON=1'b1;
    defparam M_this_external_address_q_14_LC_28_22_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_14_LC_28_22_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_external_address_q_14_LC_28_22_6 (
            .in0(N__35383),
            .in1(N__35301),
            .in2(N__35333),
            .in3(N__35316),
            .lcout(M_this_external_address_qZ0Z_14),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_13),
            .carryout(un1_M_this_external_address_q_cry_14),
            .clk(N__34637),
            .ce(),
            .sr(N__34982));
    defparam M_this_external_address_q_15_LC_28_22_7.C_ON=1'b0;
    defparam M_this_external_address_q_15_LC_28_22_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_15_LC_28_22_7.LUT_INIT=16'b1101000111100010;
    LogicCell40 M_this_external_address_q_15_LC_28_22_7 (
            .in0(N__35108),
            .in1(N__35309),
            .in2(N__35201),
            .in3(N__35127),
            .lcout(M_this_external_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34637),
            .ce(),
            .sr(N__34982));
    defparam \this_reset_cond.M_stage_q_9_LC_32_18_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_9_LC_32_18_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_9_LC_32_18_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_9_LC_32_18_4  (
            .in0(N__34854),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34746),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34638),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
